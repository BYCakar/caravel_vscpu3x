magic
tech sky130A
magscale 1 2
timestamp 1655420456
<< metal1 >>
rect 235166 700272 235172 700324
rect 235224 700312 235230 700324
rect 304258 700312 304264 700324
rect 235224 700284 304264 700312
rect 235224 700272 235230 700284
rect 304258 700272 304264 700284
rect 304316 700272 304322 700324
rect 137738 683136 137744 683188
rect 137796 683176 137802 683188
rect 580166 683176 580172 683188
rect 137796 683148 580172 683176
rect 137796 683136 137802 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 59078 649272 59084 649324
rect 59136 649312 59142 649324
rect 542354 649312 542360 649324
rect 59136 649284 542360 649312
rect 59136 649272 59142 649284
rect 542354 649272 542360 649284
rect 542412 649272 542418 649324
rect 104894 647844 104900 647896
rect 104952 647884 104958 647896
rect 429378 647884 429384 647896
rect 104952 647856 429384 647884
rect 104952 647844 104958 647856
rect 429378 647844 429384 647856
rect 429436 647844 429442 647896
rect 299474 646484 299480 646536
rect 299532 646524 299538 646536
rect 401134 646524 401140 646536
rect 299532 646496 401140 646524
rect 299532 646484 299538 646496
rect 401134 646484 401140 646496
rect 401192 646484 401198 646536
rect 169754 645124 169760 645176
rect 169812 645164 169818 645176
rect 430574 645164 430580 645176
rect 169812 645136 430580 645164
rect 169812 645124 169818 645136
rect 430574 645124 430580 645136
rect 430632 645124 430638 645176
rect 364334 643696 364340 643748
rect 364392 643736 364398 643748
rect 423674 643736 423680 643748
rect 364392 643708 423680 643736
rect 364392 643696 364398 643708
rect 423674 643696 423680 643708
rect 423732 643696 423738 643748
rect 317046 643152 317052 643204
rect 317104 643192 317110 643204
rect 430758 643192 430764 643204
rect 317104 643164 430764 643192
rect 317104 643152 317110 643164
rect 430758 643152 430764 643164
rect 430816 643152 430822 643204
rect 284938 643084 284944 643136
rect 284996 643124 285002 643136
rect 430666 643124 430672 643136
rect 284996 643096 430672 643124
rect 284996 643084 285002 643096
rect 430666 643084 430672 643096
rect 430724 643084 430730 643136
rect 318794 642336 318800 642388
rect 318852 642376 318858 642388
rect 494054 642376 494060 642388
rect 318852 642348 494060 642376
rect 318852 642336 318858 642348
rect 494054 642336 494060 642348
rect 494112 642336 494118 642388
rect 289814 641724 289820 641776
rect 289872 641764 289878 641776
rect 435358 641764 435364 641776
rect 289872 641736 435364 641764
rect 289872 641724 289878 641736
rect 435358 641724 435364 641736
rect 435416 641724 435422 641776
rect 287698 641180 287704 641232
rect 287756 641220 287762 641232
rect 378594 641220 378600 641232
rect 287756 641192 378600 641220
rect 287756 641180 287762 641192
rect 378594 641180 378600 641192
rect 378652 641180 378658 641232
rect 311250 641112 311256 641164
rect 311308 641152 311314 641164
rect 332870 641152 332876 641164
rect 311308 641124 332876 641152
rect 311308 641112 311314 641124
rect 332870 641112 332876 641124
rect 332928 641112 332934 641164
rect 312630 641044 312636 641096
rect 312688 641084 312694 641096
rect 337378 641084 337384 641096
rect 312688 641056 337384 641084
rect 312688 641044 312694 641056
rect 337378 641044 337384 641056
rect 337436 641044 337442 641096
rect 319622 640976 319628 641028
rect 319680 641016 319686 641028
rect 355410 641016 355416 641028
rect 319680 640988 355416 641016
rect 319680 640976 319686 640988
rect 355410 640976 355416 640988
rect 355468 640976 355474 641028
rect 315298 640908 315304 640960
rect 315356 640948 315362 640960
rect 359918 640948 359924 640960
rect 315356 640920 359924 640948
rect 315356 640908 315362 640920
rect 359918 640908 359924 640920
rect 359976 640908 359982 640960
rect 316678 640840 316684 640892
rect 316736 640880 316742 640892
rect 364426 640880 364432 640892
rect 316736 640852 364432 640880
rect 316736 640840 316742 640852
rect 364426 640840 364432 640852
rect 364484 640840 364490 640892
rect 302878 640772 302884 640824
rect 302936 640812 302942 640824
rect 350902 640812 350908 640824
rect 302936 640784 350908 640812
rect 302936 640772 302942 640784
rect 350902 640772 350908 640784
rect 350960 640772 350966 640824
rect 319806 640704 319812 640756
rect 319864 640744 319870 640756
rect 373442 640744 373448 640756
rect 319864 640716 373448 640744
rect 319864 640704 319870 640716
rect 373442 640704 373448 640716
rect 373500 640704 373506 640756
rect 314010 640636 314016 640688
rect 314068 640676 314074 640688
rect 368934 640676 368940 640688
rect 314068 640648 368940 640676
rect 314068 640636 314074 640648
rect 368934 640636 368940 640648
rect 368992 640636 368998 640688
rect 316862 640568 316868 640620
rect 316920 640608 316926 640620
rect 387610 640608 387616 640620
rect 316920 640580 387616 640608
rect 316920 640568 316926 640580
rect 387610 640568 387616 640580
rect 387668 640568 387674 640620
rect 309778 640500 309784 640552
rect 309836 640540 309842 640552
rect 383102 640540 383108 640552
rect 309836 640512 383108 640540
rect 309836 640500 309842 640512
rect 383102 640500 383108 640512
rect 383160 640500 383166 640552
rect 316954 640432 316960 640484
rect 317012 640472 317018 640484
rect 396626 640472 396632 640484
rect 317012 640444 396632 640472
rect 317012 640432 317018 640444
rect 396626 640432 396632 640444
rect 396684 640432 396690 640484
rect 318150 640364 318156 640416
rect 318208 640404 318214 640416
rect 428182 640404 428188 640416
rect 318208 640376 428188 640404
rect 318208 640364 318214 640376
rect 428182 640364 428188 640376
rect 428240 640364 428246 640416
rect 319530 640296 319536 640348
rect 319588 640336 319594 640348
rect 323854 640336 323860 640348
rect 319588 640308 323860 640336
rect 319588 640296 319594 640308
rect 323854 640296 323860 640308
rect 323912 640296 323918 640348
rect 414658 640296 414664 640348
rect 414716 640336 414722 640348
rect 457438 640336 457444 640348
rect 414716 640308 457444 640336
rect 414716 640296 414722 640308
rect 457438 640296 457444 640308
rect 457496 640296 457502 640348
rect 280706 639616 280712 639668
rect 280764 639656 280770 639668
rect 341886 639656 341892 639668
rect 280764 639628 341892 639656
rect 280764 639616 280770 639628
rect 341886 639616 341892 639628
rect 341944 639616 341950 639668
rect 298094 639548 298100 639600
rect 298152 639588 298158 639600
rect 428458 639588 428464 639600
rect 298152 639560 428464 639588
rect 298152 639548 298158 639560
rect 428458 639548 428464 639560
rect 428516 639548 428522 639600
rect 296714 639480 296720 639532
rect 296772 639520 296778 639532
rect 432598 639520 432604 639532
rect 296772 639492 432604 639520
rect 296772 639480 296778 639492
rect 432598 639480 432604 639492
rect 432656 639480 432662 639532
rect 291194 639412 291200 639464
rect 291252 639452 291258 639464
rect 429838 639452 429844 639464
rect 291252 639424 429844 639452
rect 291252 639412 291258 639424
rect 429838 639412 429844 639424
rect 429896 639412 429902 639464
rect 318334 639344 318340 639396
rect 318392 639384 318398 639396
rect 457530 639384 457536 639396
rect 318392 639356 457536 639384
rect 318392 639344 318398 639356
rect 457530 639344 457536 639356
rect 457588 639344 457594 639396
rect 319438 639276 319444 639328
rect 319496 639316 319502 639328
rect 470594 639316 470600 639328
rect 319496 639288 470600 639316
rect 319496 639276 319502 639288
rect 470594 639276 470600 639288
rect 470652 639276 470658 639328
rect 293954 639208 293960 639260
rect 294012 639248 294018 639260
rect 511994 639248 512000 639260
rect 294012 639220 512000 639248
rect 294012 639208 294018 639220
rect 511994 639208 512000 639220
rect 512052 639208 512058 639260
rect 287054 639140 287060 639192
rect 287112 639180 287118 639192
rect 510614 639180 510620 639192
rect 287112 639152 510620 639180
rect 287112 639140 287118 639152
rect 510614 639140 510620 639152
rect 510672 639140 510678 639192
rect 219158 639072 219164 639124
rect 219216 639112 219222 639124
rect 580258 639112 580264 639124
rect 219216 639084 580264 639112
rect 219216 639072 219222 639084
rect 580258 639072 580264 639084
rect 580316 639072 580322 639124
rect 18598 639004 18604 639056
rect 18656 639044 18662 639056
rect 409874 639044 409880 639056
rect 18656 639016 409880 639044
rect 18656 639004 18662 639016
rect 409874 639004 409880 639016
rect 409932 639004 409938 639056
rect 218698 638936 218704 638988
rect 218756 638976 218762 638988
rect 414566 638976 414572 638988
rect 218756 638948 414572 638976
rect 218756 638936 218762 638948
rect 414566 638936 414572 638948
rect 414624 638936 414630 638988
rect 311158 637644 311164 637696
rect 311216 637684 311222 637696
rect 317966 637684 317972 637696
rect 311216 637656 317972 637684
rect 311216 637644 311222 637656
rect 317966 637644 317972 637656
rect 318024 637644 318030 637696
rect 288434 637576 288440 637628
rect 288492 637616 288498 637628
rect 512086 637616 512092 637628
rect 288492 637588 512092 637616
rect 288492 637576 288498 637588
rect 512086 637576 512092 637588
rect 512144 637576 512150 637628
rect 3418 636828 3424 636880
rect 3476 636868 3482 636880
rect 316770 636868 316776 636880
rect 3476 636840 316776 636868
rect 3476 636828 3482 636840
rect 316770 636828 316776 636840
rect 316828 636828 316834 636880
rect 114186 634040 114192 634092
rect 114244 634080 114250 634092
rect 121638 634080 121644 634092
rect 114244 634052 121644 634080
rect 114244 634040 114250 634052
rect 121638 634040 121644 634052
rect 121696 634040 121702 634092
rect 131114 634040 131120 634092
rect 131172 634080 131178 634092
rect 151262 634080 151268 634092
rect 131172 634052 151268 634080
rect 131172 634040 131178 634052
rect 151262 634040 151268 634052
rect 151320 634040 151326 634092
rect 210418 634040 210424 634092
rect 210476 634080 210482 634092
rect 219710 634080 219716 634092
rect 210476 634052 219716 634080
rect 210476 634040 210482 634052
rect 219710 634040 219716 634052
rect 219768 634040 219774 634092
rect 115658 633972 115664 634024
rect 115716 634012 115722 634024
rect 124582 634012 124588 634024
rect 115716 633984 124588 634012
rect 115716 633972 115722 633984
rect 124582 633972 124588 633984
rect 124640 633972 124646 634024
rect 135254 633972 135260 634024
rect 135312 634012 135318 634024
rect 183554 634012 183560 634024
rect 135312 633984 183560 634012
rect 135312 633972 135318 633984
rect 183554 633972 183560 633984
rect 183612 633972 183618 634024
rect 213914 633972 213920 634024
rect 213972 634012 213978 634024
rect 225414 634012 225420 634024
rect 213972 633984 225420 634012
rect 213972 633972 213978 633984
rect 225414 633972 225420 633984
rect 225472 633972 225478 634024
rect 112530 633904 112536 633956
rect 112588 633944 112594 633956
rect 123018 633944 123024 633956
rect 112588 633916 123024 633944
rect 112588 633904 112594 633916
rect 123018 633904 123024 633916
rect 123076 633904 123082 633956
rect 135162 633904 135168 633956
rect 135220 633944 135226 633956
rect 160278 633944 160284 633956
rect 135220 633916 160284 633944
rect 135220 633904 135226 633916
rect 160278 633904 160284 633916
rect 160336 633904 160342 633956
rect 212534 633904 212540 633956
rect 212592 633944 212598 633956
rect 271874 633944 271880 633956
rect 212592 633916 271880 633944
rect 212592 633904 212598 633916
rect 271874 633904 271880 633916
rect 271932 633904 271938 633956
rect 69290 633836 69296 633888
rect 69348 633876 69354 633888
rect 127066 633876 127072 633888
rect 69348 633848 127072 633876
rect 69348 633836 69354 633848
rect 127066 633836 127072 633848
rect 127124 633836 127130 633888
rect 136542 633836 136548 633888
rect 136600 633876 136606 633888
rect 162854 633876 162860 633888
rect 136600 633848 162860 633876
rect 136600 633836 136606 633848
rect 162854 633836 162860 633848
rect 162912 633836 162918 633888
rect 217870 633836 217876 633888
rect 217928 633876 217934 633888
rect 242894 633876 242900 633888
rect 217928 633848 242900 633876
rect 217928 633836 217934 633848
rect 242894 633836 242900 633848
rect 242952 633836 242958 633888
rect 106642 633768 106648 633820
rect 106700 633808 106706 633820
rect 121454 633808 121460 633820
rect 106700 633780 121460 633808
rect 106700 633768 106706 633780
rect 121454 633768 121460 633780
rect 121512 633768 121518 633820
rect 139118 633768 139124 633820
rect 139176 633808 139182 633820
rect 166166 633808 166172 633820
rect 139176 633780 166172 633808
rect 139176 633768 139182 633780
rect 166166 633768 166172 633780
rect 166224 633768 166230 633820
rect 218882 633768 218888 633820
rect 218940 633808 218946 633820
rect 251910 633808 251916 633820
rect 218940 633780 251916 633808
rect 218940 633768 218946 633780
rect 251910 633768 251916 633780
rect 251968 633768 251974 633820
rect 122834 633740 122840 633752
rect 114296 633712 122840 633740
rect 56502 633632 56508 633684
rect 56560 633672 56566 633684
rect 77294 633672 77300 633684
rect 56560 633644 77300 633672
rect 56560 633632 56566 633644
rect 77294 633632 77300 633644
rect 77352 633632 77358 633684
rect 104066 633632 104072 633684
rect 104124 633672 104130 633684
rect 114186 633672 114192 633684
rect 104124 633644 114192 633672
rect 104124 633632 104130 633644
rect 114186 633632 114192 633644
rect 114244 633632 114250 633684
rect 54846 633564 54852 633616
rect 54904 633604 54910 633616
rect 88702 633604 88708 633616
rect 54904 633576 88708 633604
rect 54904 633564 54910 633576
rect 88702 633564 88708 633576
rect 88760 633564 88766 633616
rect 100662 633564 100668 633616
rect 100720 633604 100726 633616
rect 114296 633604 114324 633712
rect 122834 633700 122840 633712
rect 122892 633700 122898 633752
rect 139210 633700 139216 633752
rect 139268 633740 139274 633752
rect 174446 633740 174452 633752
rect 139268 633712 174452 633740
rect 139268 633700 139274 633712
rect 174446 633700 174452 633712
rect 174504 633700 174510 633752
rect 218790 633700 218796 633752
rect 218848 633740 218854 633752
rect 263594 633740 263600 633752
rect 218848 633712 263600 633740
rect 218848 633700 218854 633712
rect 263594 633700 263600 633712
rect 263652 633700 263658 633752
rect 118234 633632 118240 633684
rect 118292 633672 118298 633684
rect 124306 633672 124312 633684
rect 118292 633644 124312 633672
rect 118292 633632 118298 633644
rect 124306 633632 124312 633644
rect 124364 633632 124370 633684
rect 134886 633632 134892 633684
rect 134944 633672 134950 633684
rect 180334 633672 180340 633684
rect 134944 633644 180340 633672
rect 134944 633632 134950 633644
rect 180334 633632 180340 633644
rect 180392 633632 180398 633684
rect 189994 633632 190000 633684
rect 190052 633672 190058 633684
rect 204438 633672 204444 633684
rect 190052 633644 204444 633672
rect 190052 633632 190058 633644
rect 204438 633632 204444 633644
rect 204496 633632 204502 633684
rect 209774 633632 209780 633684
rect 209832 633672 209838 633684
rect 260190 633672 260196 633684
rect 209832 633644 260196 633672
rect 209832 633632 209838 633644
rect 260190 633632 260196 633644
rect 260248 633632 260254 633684
rect 100720 633576 114324 633604
rect 100720 633564 100726 633576
rect 124214 633564 124220 633616
rect 124272 633604 124278 633616
rect 171870 633604 171876 633616
rect 124272 633576 171876 633604
rect 124272 633564 124278 633576
rect 171870 633564 171876 633576
rect 171928 633564 171934 633616
rect 214006 633564 214012 633616
rect 214064 633604 214070 633616
rect 269206 633604 269212 633616
rect 214064 633576 269212 633604
rect 214064 633564 214070 633576
rect 269206 633564 269212 633576
rect 269264 633564 269270 633616
rect 55122 633496 55128 633548
rect 55180 633536 55186 633548
rect 91830 633536 91836 633548
rect 55180 633508 91836 633536
rect 55180 633496 55186 633508
rect 91830 633496 91836 633508
rect 91888 633496 91894 633548
rect 95050 633496 95056 633548
rect 95108 633536 95114 633548
rect 120902 633536 120908 633548
rect 95108 633508 120908 633536
rect 95108 633496 95114 633508
rect 120902 633496 120908 633508
rect 120960 633496 120966 633548
rect 137646 633496 137652 633548
rect 137704 633536 137710 633548
rect 137704 633508 139808 633536
rect 137704 633496 137710 633508
rect 109954 633428 109960 633480
rect 110012 633468 110018 633480
rect 120994 633468 121000 633480
rect 110012 633440 121000 633468
rect 110012 633428 110018 633440
rect 120994 633428 121000 633440
rect 121052 633428 121058 633480
rect 133874 633428 133880 633480
rect 133932 633468 133938 633480
rect 139670 633468 139676 633480
rect 133932 633440 139676 633468
rect 133932 633428 133938 633440
rect 139670 633428 139676 633440
rect 139728 633428 139734 633480
rect 139780 633400 139808 633508
rect 140130 633496 140136 633548
rect 140188 633536 140194 633548
rect 157518 633536 157524 633548
rect 140188 633508 157524 633536
rect 140188 633496 140194 633508
rect 157518 633496 157524 633508
rect 157576 633496 157582 633548
rect 192570 633496 192576 633548
rect 192628 633536 192634 633548
rect 201678 633536 201684 633548
rect 192628 633508 201684 633536
rect 192628 633496 192634 633508
rect 201678 633496 201684 633508
rect 201736 633496 201742 633548
rect 219342 633496 219348 633548
rect 219400 633536 219406 633548
rect 275094 633536 275100 633548
rect 219400 633508 275100 633536
rect 219400 633496 219406 633508
rect 275094 633496 275100 633508
rect 275152 633496 275158 633548
rect 186498 633468 186504 633480
rect 140056 633440 186504 633468
rect 140056 633400 140084 633440
rect 186498 633428 186504 633440
rect 186556 633428 186562 633480
rect 195698 633428 195704 633480
rect 195756 633468 195762 633480
rect 200850 633468 200856 633480
rect 195756 633440 200856 633468
rect 195756 633428 195762 633440
rect 200850 633428 200856 633440
rect 200908 633428 200914 633480
rect 217318 633428 217324 633480
rect 217376 633468 217382 633480
rect 231302 633468 231308 633480
rect 217376 633440 231308 633468
rect 217376 633428 217382 633440
rect 231302 633428 231308 633440
rect 231360 633428 231366 633480
rect 270402 633428 270408 633480
rect 270460 633468 270466 633480
rect 277670 633468 277676 633480
rect 270460 633440 277676 633468
rect 270460 633428 270466 633440
rect 277670 633428 277676 633440
rect 277728 633428 277734 633480
rect 139780 633372 140084 633400
rect 204254 632680 204260 632732
rect 204312 632720 204318 632732
rect 270402 632720 270408 632732
rect 204312 632692 270408 632720
rect 204312 632680 204318 632692
rect 270402 632680 270408 632692
rect 270460 632680 270466 632732
rect 215294 632272 215300 632324
rect 215352 632312 215358 632324
rect 234614 632312 234620 632324
rect 215352 632284 234620 632312
rect 215352 632272 215358 632284
rect 234614 632272 234620 632284
rect 234672 632272 234678 632324
rect 208394 632204 208400 632256
rect 208452 632244 208458 632256
rect 240318 632244 240324 632256
rect 208452 632216 240324 632244
rect 208452 632204 208458 632216
rect 240318 632204 240324 632216
rect 240376 632204 240382 632256
rect 206278 632136 206284 632188
rect 206336 632176 206342 632188
rect 254486 632176 254492 632188
rect 206336 632148 254492 632176
rect 206336 632136 206342 632148
rect 254486 632136 254492 632148
rect 254544 632136 254550 632188
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 313918 632108 313924 632120
rect 3476 632080 313924 632108
rect 3476 632068 3482 632080
rect 313918 632068 313924 632080
rect 313976 632068 313982 632120
rect 59354 631320 59360 631372
rect 59412 631360 59418 631372
rect 97718 631360 97724 631372
rect 59412 631332 97724 631360
rect 59412 631320 59418 631332
rect 97718 631320 97724 631332
rect 97776 631320 97782 631372
rect 134978 631048 134984 631100
rect 135036 631088 135042 631100
rect 142982 631088 142988 631100
rect 135036 631060 142988 631088
rect 135036 631048 135042 631060
rect 142982 631048 142988 631060
rect 143040 631048 143046 631100
rect 217962 631048 217968 631100
rect 218020 631088 218026 631100
rect 228726 631088 228732 631100
rect 218020 631060 228732 631088
rect 218020 631048 218026 631060
rect 228726 631048 228732 631060
rect 228784 631048 228790 631100
rect 124858 630980 124864 631032
rect 124916 631020 124922 631032
rect 178126 631020 178132 631032
rect 124916 630992 178132 631020
rect 124916 630980 124922 630992
rect 178126 630980 178132 630992
rect 178184 630980 178190 631032
rect 204346 630980 204352 631032
rect 204404 631020 204410 631032
rect 222838 631020 222844 631032
rect 204404 630992 222844 631020
rect 204404 630980 204410 630992
rect 222838 630980 222844 630992
rect 222896 630980 222902 631032
rect 57790 630912 57796 630964
rect 57848 630952 57854 630964
rect 80238 630952 80244 630964
rect 57848 630924 80244 630952
rect 57848 630912 57854 630924
rect 80238 630912 80244 630924
rect 80296 630912 80302 630964
rect 136450 630912 136456 630964
rect 136508 630952 136514 630964
rect 149146 630952 149152 630964
rect 136508 630924 149152 630952
rect 136508 630912 136514 630924
rect 149146 630912 149152 630924
rect 149204 630912 149210 630964
rect 204898 630912 204904 630964
rect 204956 630952 204962 630964
rect 237282 630952 237288 630964
rect 204956 630924 237288 630952
rect 204956 630912 204962 630924
rect 237282 630912 237288 630924
rect 237340 630912 237346 630964
rect 59262 630844 59268 630896
rect 59320 630884 59326 630896
rect 65518 630884 65524 630896
rect 59320 630856 65524 630884
rect 59320 630844 59326 630856
rect 65518 630844 65524 630856
rect 65576 630844 65582 630896
rect 135070 630844 135076 630896
rect 135128 630884 135134 630896
rect 154574 630884 154580 630896
rect 135128 630856 154580 630884
rect 135128 630844 135134 630856
rect 154574 630844 154580 630856
rect 154632 630844 154638 630896
rect 206370 630844 206376 630896
rect 206428 630884 206434 630896
rect 248690 630884 248696 630896
rect 206428 630856 248696 630884
rect 206428 630844 206434 630856
rect 248690 630844 248696 630856
rect 248748 630844 248754 630896
rect 56410 630776 56416 630828
rect 56468 630816 56474 630828
rect 71222 630816 71228 630828
rect 56468 630788 71228 630816
rect 56468 630776 56474 630788
rect 71222 630776 71228 630788
rect 71280 630776 71286 630828
rect 136634 630776 136640 630828
rect 136692 630816 136698 630828
rect 168742 630816 168748 630828
rect 136692 630788 168748 630816
rect 136692 630776 136698 630788
rect 168742 630776 168748 630788
rect 168800 630776 168806 630828
rect 213178 630776 213184 630828
rect 213236 630816 213242 630828
rect 257614 630816 257620 630828
rect 213236 630788 257620 630816
rect 213236 630776 213242 630788
rect 257614 630776 257620 630788
rect 257672 630776 257678 630828
rect 54938 630708 54944 630760
rect 54996 630748 55002 630760
rect 74626 630748 74632 630760
rect 54996 630720 74632 630748
rect 54996 630708 55002 630720
rect 74626 630708 74632 630720
rect 74684 630708 74690 630760
rect 86770 630708 86776 630760
rect 86828 630748 86834 630760
rect 124490 630748 124496 630760
rect 86828 630720 124496 630748
rect 86828 630708 86834 630720
rect 124490 630708 124496 630720
rect 124548 630708 124554 630760
rect 137830 630708 137836 630760
rect 137888 630748 137894 630760
rect 145558 630748 145564 630760
rect 137888 630720 145564 630748
rect 137888 630708 137894 630720
rect 145558 630708 145564 630720
rect 145616 630708 145622 630760
rect 211798 630708 211804 630760
rect 211856 630748 211862 630760
rect 266262 630748 266268 630760
rect 211856 630720 266268 630748
rect 211856 630708 211862 630720
rect 266262 630708 266268 630720
rect 266320 630708 266326 630760
rect 55030 630640 55036 630692
rect 55088 630680 55094 630692
rect 62942 630680 62948 630692
rect 55088 630652 62948 630680
rect 55088 630640 55094 630652
rect 62942 630640 62948 630652
rect 63000 630640 63006 630692
rect 83458 630640 83464 630692
rect 83516 630680 83522 630692
rect 124398 630680 124404 630692
rect 83516 630652 124404 630680
rect 83516 630640 83522 630652
rect 124398 630640 124404 630652
rect 124456 630640 124462 630692
rect 137922 630640 137928 630692
rect 137980 630680 137986 630692
rect 218698 630680 218704 630692
rect 137980 630652 218704 630680
rect 137980 630640 137986 630652
rect 218698 630640 218704 630652
rect 218756 630640 218762 630692
rect 219434 630640 219440 630692
rect 219492 630680 219498 630692
rect 246022 630680 246028 630692
rect 219492 630652 246028 630680
rect 219492 630640 219498 630652
rect 246022 630640 246028 630652
rect 246080 630640 246086 630692
rect 280706 630504 280712 630556
rect 280764 630504 280770 630556
rect 139854 630368 139860 630420
rect 139912 630408 139918 630420
rect 140130 630408 140136 630420
rect 139912 630380 140136 630408
rect 139912 630368 139918 630380
rect 140130 630368 140136 630380
rect 140188 630368 140194 630420
rect 198274 630368 198280 630420
rect 198332 630408 198338 630420
rect 201586 630408 201592 630420
rect 198332 630380 201592 630408
rect 198332 630368 198338 630380
rect 201586 630368 201592 630380
rect 201644 630368 201650 630420
rect 280724 630352 280752 630504
rect 280706 630300 280712 630352
rect 280764 630300 280770 630352
rect 435358 630028 435364 630080
rect 435416 630068 435422 630080
rect 483198 630068 483204 630080
rect 435416 630040 483204 630068
rect 435416 630028 435422 630040
rect 483198 630028 483204 630040
rect 483256 630028 483262 630080
rect 432598 629960 432604 630012
rect 432656 630000 432662 630012
rect 494790 630000 494796 630012
rect 432656 629972 494796 630000
rect 432656 629960 432662 629972
rect 494790 629960 494796 629972
rect 494848 629960 494854 630012
rect 428458 629892 428464 629944
rect 428516 629932 428522 629944
rect 501230 629932 501236 629944
rect 428516 629904 501236 629932
rect 428516 629892 428522 629904
rect 501230 629892 501236 629904
rect 501288 629892 501294 629944
rect 294598 627920 294604 627972
rect 294656 627960 294662 627972
rect 317690 627960 317696 627972
rect 294656 627932 317696 627960
rect 294656 627920 294662 627932
rect 317690 627920 317696 627932
rect 317748 627920 317754 627972
rect 465442 627920 465448 627972
rect 465500 627960 465506 627972
rect 580258 627960 580264 627972
rect 465500 627932 580264 627960
rect 465500 627920 465506 627932
rect 580258 627920 580264 627932
rect 580316 627920 580322 627972
rect 429838 627852 429844 627904
rect 429896 627892 429902 627904
rect 456794 627892 456800 627904
rect 429896 627864 456800 627892
rect 429896 627852 429902 627864
rect 456794 627852 456800 627864
rect 456852 627852 456858 627904
rect 208486 625132 208492 625184
rect 208544 625172 208550 625184
rect 216674 625172 216680 625184
rect 208544 625144 216680 625172
rect 208544 625132 208550 625144
rect 216674 625132 216680 625144
rect 216732 625132 216738 625184
rect 312538 623772 312544 623824
rect 312596 623812 312602 623824
rect 317414 623812 317420 623824
rect 312596 623784 317420 623812
rect 312596 623772 312602 623784
rect 317414 623772 317420 623784
rect 317472 623772 317478 623824
rect 206462 619624 206468 619676
rect 206520 619664 206526 619676
rect 216674 619664 216680 619676
rect 206520 619636 216680 619664
rect 206520 619624 206526 619636
rect 216674 619624 216680 619636
rect 216732 619624 216738 619676
rect 307018 618264 307024 618316
rect 307076 618304 307082 618316
rect 317598 618304 317604 618316
rect 307076 618276 317604 618304
rect 307076 618264 307082 618276
rect 317598 618264 317604 618276
rect 317656 618264 317662 618316
rect 132494 615884 132500 615936
rect 132552 615924 132558 615936
rect 136726 615924 136732 615936
rect 132552 615896 136732 615924
rect 132552 615884 132558 615896
rect 136726 615884 136732 615896
rect 136784 615884 136790 615936
rect 204990 615476 204996 615528
rect 205048 615516 205054 615528
rect 216674 615516 216680 615528
rect 205048 615488 216680 615516
rect 205048 615476 205054 615488
rect 216674 615476 216680 615488
rect 216732 615476 216738 615528
rect 287790 614116 287796 614168
rect 287848 614156 287854 614168
rect 317966 614156 317972 614168
rect 287848 614128 317972 614156
rect 287848 614116 287854 614128
rect 317966 614116 317972 614128
rect 318024 614116 318030 614168
rect 295978 608608 295984 608660
rect 296036 608648 296042 608660
rect 317966 608648 317972 608660
rect 296036 608620 317972 608648
rect 296036 608608 296042 608620
rect 317966 608608 317972 608620
rect 318024 608608 318030 608660
rect 286318 604460 286324 604512
rect 286376 604500 286382 604512
rect 317966 604500 317972 604512
rect 286376 604472 317972 604500
rect 286376 604460 286382 604472
rect 317966 604460 317972 604472
rect 318024 604460 318030 604512
rect 126238 597524 126244 597576
rect 126296 597564 126302 597576
rect 136726 597564 136732 597576
rect 126296 597536 136732 597564
rect 126296 597524 126302 597536
rect 136726 597524 136732 597536
rect 136784 597524 136790 597576
rect 213270 597524 213276 597576
rect 213328 597564 213334 597576
rect 216674 597564 216680 597576
rect 213328 597536 216680 597564
rect 213328 597524 213334 597536
rect 216674 597524 216680 597536
rect 216732 597524 216738 597576
rect 302234 596776 302240 596828
rect 302292 596816 302298 596828
rect 318334 596816 318340 596828
rect 302292 596788 318340 596816
rect 302292 596776 302298 596788
rect 318334 596776 318340 596788
rect 318392 596776 318398 596828
rect 203242 596640 203248 596692
rect 203300 596680 203306 596692
rect 204530 596680 204536 596692
rect 203300 596652 204536 596680
rect 203300 596640 203306 596652
rect 204530 596640 204536 596652
rect 204588 596640 204594 596692
rect 124122 596164 124128 596216
rect 124180 596204 124186 596216
rect 134518 596204 134524 596216
rect 124180 596176 134524 596204
rect 124180 596164 124186 596176
rect 134518 596164 134524 596176
rect 134576 596164 134582 596216
rect 283650 596164 283656 596216
rect 283708 596204 283714 596216
rect 302234 596204 302240 596216
rect 283708 596176 302240 596204
rect 283708 596164 283714 596176
rect 302234 596164 302240 596176
rect 302292 596164 302298 596216
rect 211154 594804 211160 594856
rect 211212 594844 211218 594856
rect 216674 594844 216680 594856
rect 211212 594816 216680 594844
rect 211212 594804 211218 594816
rect 216674 594804 216680 594816
rect 216732 594804 216738 594856
rect 285030 594804 285036 594856
rect 285088 594844 285094 594856
rect 317966 594844 317972 594856
rect 285088 594816 317972 594844
rect 285088 594804 285094 594816
rect 317966 594804 317972 594816
rect 318024 594804 318030 594856
rect 210510 590656 210516 590708
rect 210568 590696 210574 590708
rect 216674 590696 216680 590708
rect 210568 590668 216680 590696
rect 210568 590656 210574 590668
rect 216674 590656 216680 590668
rect 216732 590656 216738 590708
rect 286410 589296 286416 589348
rect 286468 589336 286474 589348
rect 317966 589336 317972 589348
rect 286468 589308 317972 589336
rect 286468 589296 286474 589308
rect 317966 589296 317972 589308
rect 318024 589296 318030 589348
rect 125594 585148 125600 585200
rect 125652 585188 125658 585200
rect 136726 585188 136732 585200
rect 125652 585160 136732 585188
rect 125652 585148 125658 585160
rect 136726 585148 136732 585160
rect 136784 585148 136790 585200
rect 289078 585148 289084 585200
rect 289136 585188 289142 585200
rect 317966 585188 317972 585200
rect 289136 585160 317972 585188
rect 289136 585148 289142 585160
rect 317966 585148 317972 585160
rect 318024 585148 318030 585200
rect 128998 582360 129004 582412
rect 129056 582400 129062 582412
rect 136726 582400 136732 582412
rect 129056 582372 136732 582400
rect 129056 582360 129062 582372
rect 136726 582360 136732 582372
rect 136784 582360 136790 582412
rect 206554 582360 206560 582412
rect 206612 582400 206618 582412
rect 216674 582400 216680 582412
rect 206612 582372 216680 582400
rect 206612 582360 206618 582372
rect 216674 582360 216680 582372
rect 216732 582360 216738 582412
rect 209038 579640 209044 579692
rect 209096 579680 209102 579692
rect 216674 579680 216680 579692
rect 209096 579652 216680 579680
rect 209096 579640 209102 579652
rect 216674 579640 216680 579652
rect 216732 579640 216738 579692
rect 287882 579640 287888 579692
rect 287940 579680 287946 579692
rect 317966 579680 317972 579692
rect 287940 579652 317972 579680
rect 287940 579640 287946 579652
rect 317966 579640 317972 579652
rect 318024 579640 318030 579692
rect 513006 579640 513012 579692
rect 513064 579680 513070 579692
rect 560938 579680 560944 579692
rect 513064 579652 560944 579680
rect 513064 579640 513070 579652
rect 560938 579640 560944 579652
rect 560996 579640 561002 579692
rect 138566 572296 138572 572348
rect 138624 572336 138630 572348
rect 139118 572336 139124 572348
rect 138624 572308 139124 572336
rect 138624 572296 138630 572308
rect 139118 572296 139124 572308
rect 139176 572296 139182 572348
rect 207014 570596 207020 570648
rect 207072 570636 207078 570648
rect 217410 570636 217416 570648
rect 207072 570608 217416 570636
rect 207072 570596 207078 570608
rect 217410 570596 217416 570608
rect 217468 570596 217474 570648
rect 137370 569848 137376 569900
rect 137428 569888 137434 569900
rect 139762 569888 139768 569900
rect 137428 569860 139768 569888
rect 137428 569848 137434 569860
rect 139762 569848 139768 569860
rect 139820 569848 139826 569900
rect 200942 569848 200948 569900
rect 201000 569888 201006 569900
rect 202966 569888 202972 569900
rect 201000 569860 202972 569888
rect 201000 569848 201006 569860
rect 202966 569848 202972 569860
rect 203024 569848 203030 569900
rect 57882 569168 57888 569220
rect 57940 569208 57946 569220
rect 138014 569208 138020 569220
rect 57940 569180 138020 569208
rect 57940 569168 57946 569180
rect 138014 569168 138020 569180
rect 138072 569168 138078 569220
rect 57238 569100 57244 569152
rect 57296 569140 57302 569152
rect 59906 569140 59912 569152
rect 57296 569112 59912 569140
rect 57296 569100 57302 569112
rect 59906 569100 59912 569112
rect 59964 569100 59970 569152
rect 217686 568556 217692 568608
rect 217744 568596 217750 568608
rect 219894 568596 219900 568608
rect 217744 568568 219900 568596
rect 217744 568556 217750 568568
rect 219894 568556 219900 568568
rect 219952 568556 219958 568608
rect 3418 568488 3424 568540
rect 3476 568528 3482 568540
rect 286410 568528 286416 568540
rect 3476 568500 286416 568528
rect 3476 568488 3482 568500
rect 286410 568488 286416 568500
rect 286468 568488 286474 568540
rect 58710 568420 58716 568472
rect 58768 568460 58774 568472
rect 60734 568460 60740 568472
rect 58768 568432 60740 568460
rect 58768 568420 58774 568432
rect 60734 568420 60740 568432
rect 60792 568420 60798 568472
rect 134518 568420 134524 568472
rect 134576 568460 134582 568472
rect 204530 568460 204536 568472
rect 134576 568432 204536 568460
rect 134576 568420 134582 568432
rect 204530 568420 204536 568432
rect 204588 568460 204594 568472
rect 302234 568460 302240 568472
rect 204588 568432 302240 568460
rect 204588 568420 204594 568432
rect 302234 568420 302240 568432
rect 302292 568420 302298 568472
rect 57146 568352 57152 568404
rect 57204 568392 57210 568404
rect 61378 568392 61384 568404
rect 57204 568364 61384 568392
rect 57204 568352 57210 568364
rect 61378 568352 61384 568364
rect 61436 568352 61442 568404
rect 106274 568216 106280 568268
rect 106332 568256 106338 568268
rect 124582 568256 124588 568268
rect 106332 568228 124588 568256
rect 106332 568216 106338 568228
rect 124582 568216 124588 568228
rect 124640 568216 124646 568268
rect 164326 568216 164332 568268
rect 164384 568256 164390 568268
rect 200850 568256 200856 568268
rect 164384 568228 200856 568256
rect 164384 568216 164390 568228
rect 200850 568216 200856 568228
rect 200908 568216 200914 568268
rect 99558 568148 99564 568200
rect 99616 568188 99622 568200
rect 122190 568188 122196 568200
rect 99616 568160 122196 568188
rect 99616 568148 99622 568160
rect 122190 568148 122196 568160
rect 122248 568148 122254 568200
rect 137646 568148 137652 568200
rect 137704 568188 137710 568200
rect 145282 568188 145288 568200
rect 137704 568160 145288 568188
rect 137704 568148 137710 568160
rect 145282 568148 145288 568160
rect 145340 568148 145346 568200
rect 182358 568148 182364 568200
rect 182416 568188 182422 568200
rect 218882 568188 218888 568200
rect 182416 568160 218888 568188
rect 182416 568148 182422 568160
rect 218882 568148 218888 568160
rect 218940 568148 218946 568200
rect 96706 568080 96712 568132
rect 96764 568120 96770 568132
rect 123018 568120 123024 568132
rect 96764 568092 123024 568120
rect 96764 568080 96770 568092
rect 123018 568080 123024 568092
rect 123076 568080 123082 568132
rect 139026 568080 139032 568132
rect 139084 568120 139090 568132
rect 150618 568120 150624 568132
rect 139084 568092 150624 568120
rect 139084 568080 139090 568092
rect 150618 568080 150624 568092
rect 150676 568080 150682 568132
rect 154574 568080 154580 568132
rect 154632 568120 154638 568132
rect 201678 568120 201684 568132
rect 154632 568092 201684 568120
rect 154632 568080 154638 568092
rect 201678 568080 201684 568092
rect 201736 568080 201742 568132
rect 54846 568012 54852 568064
rect 54904 568052 54910 568064
rect 78766 568052 78772 568064
rect 54904 568024 78772 568052
rect 54904 568012 54910 568024
rect 78766 568012 78772 568024
rect 78824 568012 78830 568064
rect 93854 568012 93860 568064
rect 93912 568052 93918 568064
rect 122834 568052 122840 568064
rect 93912 568024 122840 568052
rect 93912 568012 93918 568024
rect 122834 568012 122840 568024
rect 122892 568012 122898 568064
rect 134886 568012 134892 568064
rect 134944 568052 134950 568064
rect 151814 568052 151820 568064
rect 134944 568024 151820 568052
rect 134944 568012 134950 568024
rect 151814 568012 151820 568024
rect 151872 568012 151878 568064
rect 156046 568012 156052 568064
rect 156104 568052 156110 568064
rect 204438 568052 204444 568064
rect 156104 568024 204444 568052
rect 156104 568012 156110 568024
rect 204438 568012 204444 568024
rect 204496 568012 204502 568064
rect 219342 568012 219348 568064
rect 219400 568052 219406 568064
rect 223574 568052 223580 568064
rect 219400 568024 223580 568052
rect 219400 568012 219406 568024
rect 223574 568012 223580 568024
rect 223632 568012 223638 568064
rect 242158 568012 242164 568064
rect 242216 568052 242222 568064
rect 281074 568052 281080 568064
rect 242216 568024 281080 568052
rect 242216 568012 242222 568024
rect 281074 568012 281080 568024
rect 281132 568012 281138 568064
rect 58802 567944 58808 567996
rect 58860 567984 58866 567996
rect 91094 567984 91100 567996
rect 58860 567956 91100 567984
rect 58860 567944 58866 567956
rect 91094 567944 91100 567956
rect 91152 567944 91158 567996
rect 98086 567944 98092 567996
rect 98144 567984 98150 567996
rect 120994 567984 121000 567996
rect 98144 567956 121000 567984
rect 98144 567944 98150 567956
rect 120994 567944 121000 567956
rect 121052 567944 121058 567996
rect 122190 567944 122196 567996
rect 122248 567984 122254 567996
rect 201770 567984 201776 567996
rect 122248 567956 201776 567984
rect 122248 567944 122254 567956
rect 201770 567944 201776 567956
rect 201828 567944 201834 567996
rect 217870 567944 217876 567996
rect 217928 567984 217934 567996
rect 222194 567984 222200 567996
rect 217928 567956 222200 567984
rect 217928 567944 217934 567956
rect 222194 567944 222200 567956
rect 222252 567944 222258 567996
rect 260834 567944 260840 567996
rect 260892 567984 260898 567996
rect 317046 567984 317052 567996
rect 260892 567956 317052 567984
rect 260892 567944 260898 567956
rect 317046 567944 317052 567956
rect 317104 567944 317110 567996
rect 58526 567876 58532 567928
rect 58584 567916 58590 567928
rect 67634 567916 67640 567928
rect 58584 567888 67640 567916
rect 58584 567876 58590 567888
rect 67634 567876 67640 567888
rect 67692 567876 67698 567928
rect 78674 567876 78680 567928
rect 78732 567916 78738 567928
rect 122282 567916 122288 567928
rect 78732 567888 122288 567916
rect 78732 567876 78738 567888
rect 122282 567876 122288 567888
rect 122340 567876 122346 567928
rect 139210 567876 139216 567928
rect 139268 567916 139274 567928
rect 158714 567916 158720 567928
rect 139268 567888 158720 567916
rect 139268 567876 139274 567888
rect 158714 567876 158720 567888
rect 158772 567876 158778 567928
rect 194594 567876 194600 567928
rect 194652 567916 194658 567928
rect 283558 567916 283564 567928
rect 194652 567888 283564 567916
rect 194652 567876 194658 567888
rect 283558 567876 283564 567888
rect 283616 567876 283622 567928
rect 64874 567808 64880 567860
rect 64932 567848 64938 567860
rect 123386 567848 123392 567860
rect 64932 567820 123392 567848
rect 64932 567808 64938 567820
rect 123386 567808 123392 567820
rect 123444 567808 123450 567860
rect 138566 567808 138572 567860
rect 138624 567848 138630 567860
rect 161658 567848 161664 567860
rect 138624 567820 161664 567848
rect 138624 567808 138630 567820
rect 161658 567808 161664 567820
rect 161716 567808 161722 567860
rect 179414 567808 179420 567860
rect 179472 567848 179478 567860
rect 282178 567848 282184 567860
rect 179472 567820 282184 567848
rect 179472 567808 179478 567820
rect 282178 567808 282184 567820
rect 282236 567808 282242 567860
rect 139118 567604 139124 567656
rect 139176 567644 139182 567656
rect 142154 567644 142160 567656
rect 139176 567616 142160 567644
rect 139176 567604 139182 567616
rect 142154 567604 142160 567616
rect 142212 567604 142218 567656
rect 87046 566788 87052 566840
rect 87104 566828 87110 566840
rect 121454 566828 121460 566840
rect 87104 566800 121460 566828
rect 87104 566788 87110 566800
rect 121454 566788 121460 566800
rect 121512 566788 121518 566840
rect 157978 566788 157984 566840
rect 158036 566828 158042 566840
rect 203150 566828 203156 566840
rect 158036 566800 203156 566828
rect 158036 566788 158042 566800
rect 203150 566788 203156 566800
rect 203208 566788 203214 566840
rect 111886 566720 111892 566772
rect 111944 566760 111950 566772
rect 121546 566760 121552 566772
rect 111944 566732 121552 566760
rect 111944 566720 111950 566732
rect 121546 566720 121552 566732
rect 121604 566720 121610 566772
rect 125686 566720 125692 566772
rect 125744 566760 125750 566772
rect 200758 566760 200764 566772
rect 125744 566732 200764 566760
rect 125744 566720 125750 566732
rect 200758 566720 200764 566732
rect 200816 566720 200822 566772
rect 58986 566652 58992 566704
rect 59044 566692 59050 566704
rect 77294 566692 77300 566704
rect 59044 566664 77300 566692
rect 59044 566652 59050 566664
rect 77294 566652 77300 566664
rect 77352 566652 77358 566704
rect 84194 566652 84200 566704
rect 84252 566692 84258 566704
rect 122098 566692 122104 566704
rect 84252 566664 122104 566692
rect 84252 566652 84258 566664
rect 122098 566652 122104 566664
rect 122156 566652 122162 566704
rect 200298 566652 200304 566704
rect 200356 566692 200362 566704
rect 283466 566692 283472 566704
rect 200356 566664 283472 566692
rect 200356 566652 200362 566664
rect 283466 566652 283472 566664
rect 283524 566652 283530 566704
rect 57514 566584 57520 566636
rect 57572 566624 57578 566636
rect 82906 566624 82912 566636
rect 57572 566596 82912 566624
rect 57572 566584 57578 566596
rect 82906 566584 82912 566596
rect 82964 566584 82970 566636
rect 86954 566584 86960 566636
rect 87012 566624 87018 566636
rect 124306 566624 124312 566636
rect 87012 566596 124312 566624
rect 87012 566584 87018 566596
rect 124306 566584 124312 566596
rect 124364 566584 124370 566636
rect 187786 566584 187792 566636
rect 187844 566624 187850 566636
rect 281718 566624 281724 566636
rect 187844 566596 281724 566624
rect 187844 566584 187850 566596
rect 281718 566584 281724 566596
rect 281776 566584 281782 566636
rect 69014 566516 69020 566568
rect 69072 566556 69078 566568
rect 123478 566556 123484 566568
rect 69072 566528 123484 566556
rect 69072 566516 69078 566528
rect 123478 566516 123484 566528
rect 123536 566516 123542 566568
rect 180886 566516 180892 566568
rect 180944 566556 180950 566568
rect 281902 566556 281908 566568
rect 180944 566528 281908 566556
rect 180944 566516 180950 566528
rect 281902 566516 281908 566528
rect 281960 566516 281966 566568
rect 67726 566448 67732 566500
rect 67784 566488 67790 566500
rect 121914 566488 121920 566500
rect 67784 566460 121920 566488
rect 67784 566448 67790 566460
rect 121914 566448 121920 566460
rect 121972 566448 121978 566500
rect 137186 566448 137192 566500
rect 137244 566488 137250 566500
rect 160094 566488 160100 566500
rect 137244 566460 160100 566488
rect 137244 566448 137250 566460
rect 160094 566448 160100 566460
rect 160152 566448 160158 566500
rect 180794 566448 180800 566500
rect 180852 566488 180858 566500
rect 281810 566488 281816 566500
rect 180852 566460 281816 566488
rect 180852 566448 180858 566460
rect 281810 566448 281816 566460
rect 281868 566448 281874 566500
rect 137554 566244 137560 566296
rect 137612 566284 137618 566296
rect 140774 566284 140780 566296
rect 137612 566256 140780 566284
rect 137612 566244 137618 566256
rect 140774 566244 140780 566256
rect 140832 566244 140838 566296
rect 139854 566040 139860 566092
rect 139912 566080 139918 566092
rect 140866 566080 140872 566092
rect 139912 566052 140872 566080
rect 139912 566040 139918 566052
rect 140866 566040 140872 566052
rect 140924 566040 140930 566092
rect 59078 565972 59084 566024
rect 59136 566012 59142 566024
rect 62114 566012 62120 566024
rect 59136 565984 62120 566012
rect 59136 565972 59142 565984
rect 62114 565972 62120 565984
rect 62172 565972 62178 566024
rect 267734 565836 267740 565888
rect 267792 565876 267798 565888
rect 317966 565876 317972 565888
rect 267792 565848 317972 565876
rect 267792 565836 267798 565848
rect 317966 565836 317972 565848
rect 318024 565836 318030 565888
rect 151354 565632 151360 565684
rect 151412 565672 151418 565684
rect 160738 565672 160744 565684
rect 151412 565644 160744 565672
rect 151412 565632 151418 565644
rect 160738 565632 160744 565644
rect 160796 565632 160802 565684
rect 148778 565564 148784 565616
rect 148836 565604 148842 565616
rect 159358 565604 159364 565616
rect 148836 565576 159364 565604
rect 148836 565564 148842 565576
rect 159358 565564 159364 565576
rect 159416 565564 159422 565616
rect 143534 565496 143540 565548
rect 143592 565536 143598 565548
rect 156414 565536 156420 565548
rect 143592 565508 156420 565536
rect 143592 565496 143598 565508
rect 156414 565496 156420 565508
rect 156472 565496 156478 565548
rect 159910 565496 159916 565548
rect 159968 565536 159974 565548
rect 164878 565536 164884 565548
rect 159968 565508 164884 565536
rect 159968 565496 159974 565508
rect 164878 565496 164884 565508
rect 164936 565496 164942 565548
rect 82722 565428 82728 565480
rect 82780 565468 82786 565480
rect 89806 565468 89812 565480
rect 82780 565440 89812 565468
rect 82780 565428 82786 565440
rect 89806 565428 89812 565440
rect 89864 565428 89870 565480
rect 147766 565428 147772 565480
rect 147824 565468 147830 565480
rect 162302 565468 162308 565480
rect 147824 565440 162308 565468
rect 147824 565428 147830 565440
rect 162302 565428 162308 565440
rect 162360 565428 162366 565480
rect 231854 565428 231860 565480
rect 231912 565468 231918 565480
rect 259638 565468 259644 565480
rect 231912 565440 259644 565468
rect 231912 565428 231918 565440
rect 259638 565428 259644 565440
rect 259696 565428 259702 565480
rect 74534 565360 74540 565412
rect 74592 565400 74598 565412
rect 96982 565400 96988 565412
rect 74592 565372 96988 565400
rect 74592 565360 74598 565372
rect 96982 565360 96988 565372
rect 97040 565360 97046 565412
rect 100202 565360 100208 565412
rect 100260 565400 100266 565412
rect 115198 565400 115204 565412
rect 100260 565372 115204 565400
rect 100260 565360 100266 565372
rect 115198 565360 115204 565372
rect 115256 565360 115262 565412
rect 154666 565360 154672 565412
rect 154724 565400 154730 565412
rect 171318 565400 171324 565412
rect 154724 565372 171324 565400
rect 154724 565360 154730 565372
rect 171318 565360 171324 565372
rect 171376 565360 171382 565412
rect 182818 565360 182824 565412
rect 182876 565400 182882 565412
rect 182876 565372 190454 565400
rect 182876 565360 182882 565372
rect 77018 565292 77024 565344
rect 77076 565332 77082 565344
rect 84838 565332 84844 565344
rect 77076 565304 84844 565332
rect 77076 565292 77082 565304
rect 84838 565292 84844 565304
rect 84896 565292 84902 565344
rect 86034 565292 86040 565344
rect 86092 565332 86098 565344
rect 108298 565332 108304 565344
rect 86092 565304 108304 565332
rect 86092 565292 86098 565304
rect 108298 565292 108304 565304
rect 108356 565292 108362 565344
rect 129734 565292 129740 565344
rect 129792 565332 129798 565344
rect 153838 565332 153844 565344
rect 129792 565304 153844 565332
rect 129792 565292 129798 565304
rect 153838 565292 153844 565304
rect 153896 565292 153902 565344
rect 158806 565292 158812 565344
rect 158864 565332 158870 565344
rect 182910 565332 182916 565344
rect 158864 565304 182916 565332
rect 158864 565292 158870 565304
rect 182910 565292 182916 565304
rect 182968 565292 182974 565344
rect 190426 565332 190454 565372
rect 222378 565360 222384 565412
rect 222436 565400 222442 565412
rect 253934 565400 253940 565412
rect 222436 565372 253940 565400
rect 222436 565360 222442 565372
rect 253934 565360 253940 565372
rect 253992 565360 253998 565412
rect 203334 565332 203340 565344
rect 190426 565304 203340 565332
rect 203334 565292 203340 565304
rect 203392 565292 203398 565344
rect 212626 565292 212632 565344
rect 212684 565332 212690 565344
rect 251266 565332 251272 565344
rect 212684 565304 251272 565332
rect 212684 565292 212690 565304
rect 251266 565292 251272 565304
rect 251324 565292 251330 565344
rect 252554 565292 252560 565344
rect 252612 565332 252618 565344
rect 316954 565332 316960 565344
rect 252612 565304 316960 565332
rect 252612 565292 252618 565304
rect 316954 565292 316960 565304
rect 317012 565292 317018 565344
rect 68738 565224 68744 565276
rect 68796 565264 68802 565276
rect 105538 565264 105544 565276
rect 68796 565236 105544 565264
rect 68796 565224 68802 565236
rect 105538 565224 105544 565236
rect 105596 565224 105602 565276
rect 118694 565224 118700 565276
rect 118752 565264 118758 565276
rect 145098 565264 145104 565276
rect 118752 565236 145104 565264
rect 118752 565224 118758 565236
rect 145098 565224 145104 565236
rect 145156 565224 145162 565276
rect 147674 565224 147680 565276
rect 147732 565264 147738 565276
rect 185486 565264 185492 565276
rect 147732 565236 185492 565264
rect 147732 565224 147738 565236
rect 185486 565224 185492 565236
rect 185544 565224 185550 565276
rect 190638 565224 190644 565276
rect 190696 565264 190702 565276
rect 257062 565264 257068 565276
rect 190696 565236 257068 565264
rect 190696 565224 190702 565236
rect 257062 565224 257068 565236
rect 257120 565224 257126 565276
rect 269114 565224 269120 565276
rect 269172 565264 269178 565276
rect 289078 565264 289084 565276
rect 269172 565236 289084 565264
rect 269172 565224 269178 565236
rect 289078 565224 289084 565236
rect 289136 565224 289142 565276
rect 71314 565156 71320 565208
rect 71372 565196 71378 565208
rect 108390 565196 108396 565208
rect 71372 565168 108396 565196
rect 71372 565156 71378 565168
rect 108390 565156 108396 565168
rect 108448 565156 108454 565208
rect 110414 565156 110420 565208
rect 110472 565196 110478 565208
rect 120718 565196 120724 565208
rect 110472 565168 120724 565196
rect 110472 565156 110478 565168
rect 120718 565156 120724 565168
rect 120776 565156 120782 565208
rect 133966 565156 133972 565208
rect 134024 565196 134030 565208
rect 197446 565196 197452 565208
rect 134024 565168 197452 565196
rect 134024 565156 134030 565168
rect 197446 565156 197452 565168
rect 197504 565156 197510 565208
rect 227714 565156 227720 565208
rect 227772 565196 227778 565208
rect 245654 565196 245660 565208
rect 227772 565168 245660 565196
rect 227772 565156 227778 565168
rect 245654 565156 245660 565168
rect 245712 565156 245718 565208
rect 247034 565156 247040 565208
rect 247092 565196 247098 565208
rect 319806 565196 319812 565208
rect 247092 565168 319812 565196
rect 247092 565156 247098 565168
rect 319806 565156 319812 565168
rect 319864 565156 319870 565208
rect 62850 565088 62856 565140
rect 62908 565128 62914 565140
rect 72418 565128 72424 565140
rect 62908 565100 72424 565128
rect 62908 565088 62914 565100
rect 72418 565088 72424 565100
rect 72476 565088 72482 565140
rect 75914 565088 75920 565140
rect 75972 565128 75978 565140
rect 117406 565128 117412 565140
rect 75972 565100 117412 565128
rect 75972 565088 75978 565100
rect 117406 565088 117412 565100
rect 117464 565088 117470 565140
rect 132586 565088 132592 565140
rect 132644 565128 132650 565140
rect 177022 565128 177028 565140
rect 132644 565100 177028 565128
rect 132644 565088 132650 565100
rect 177022 565088 177028 565100
rect 177080 565088 177086 565140
rect 191834 565088 191840 565140
rect 191892 565128 191898 565140
rect 276934 565128 276940 565140
rect 191892 565100 276940 565128
rect 191892 565088 191898 565100
rect 276934 565088 276940 565100
rect 276992 565088 276998 565140
rect 60274 565020 60280 565072
rect 60332 565060 60338 565072
rect 62574 565060 62580 565072
rect 60332 565032 62580 565060
rect 60332 565020 60338 565032
rect 62574 565020 62580 565032
rect 62632 565020 62638 565072
rect 94498 564884 94504 564936
rect 94556 564924 94562 564936
rect 102778 564924 102784 564936
rect 94556 564896 102784 564924
rect 94556 564884 94562 564896
rect 102778 564884 102784 564896
rect 102836 564884 102842 564936
rect 187694 564884 187700 564936
rect 187752 564924 187758 564936
rect 191190 564924 191196 564936
rect 187752 564896 191196 564924
rect 187752 564884 187758 564896
rect 191190 564884 191196 564896
rect 191248 564884 191254 564936
rect 113174 564476 113180 564528
rect 113232 564516 113238 564528
rect 121178 564516 121184 564528
rect 113232 564488 121184 564516
rect 113232 564476 113238 564488
rect 121178 564476 121184 564488
rect 121236 564476 121242 564528
rect 71774 564408 71780 564460
rect 71832 564448 71838 564460
rect 73798 564448 73804 564460
rect 71832 564420 73804 564448
rect 71832 564408 71838 564420
rect 73798 564408 73804 564420
rect 73856 564408 73862 564460
rect 100754 564408 100760 564460
rect 100812 564448 100818 564460
rect 102870 564448 102876 564460
rect 100812 564420 102876 564448
rect 100812 564408 100818 564420
rect 102870 564408 102876 564420
rect 102928 564408 102934 564460
rect 106918 564408 106924 564460
rect 106976 564448 106982 564460
rect 108574 564448 108580 564460
rect 106976 564420 108580 564448
rect 106976 564408 106982 564420
rect 108574 564408 108580 564420
rect 108632 564408 108638 564460
rect 116578 564408 116584 564460
rect 116636 564448 116642 564460
rect 120166 564448 120172 564460
rect 116636 564420 120172 564448
rect 116636 564408 116642 564420
rect 120166 564408 120172 564420
rect 120224 564408 120230 564460
rect 173158 564408 173164 564460
rect 173216 564448 173222 564460
rect 173986 564448 173992 564460
rect 173216 564420 173992 564448
rect 173216 564408 173222 564420
rect 173986 564408 173992 564420
rect 174044 564408 174050 564460
rect 197998 564408 198004 564460
rect 198056 564448 198062 564460
rect 200206 564448 200212 564460
rect 198056 564420 200212 564448
rect 198056 564408 198062 564420
rect 200206 564408 200212 564420
rect 200264 564408 200270 564460
rect 225138 564408 225144 564460
rect 225196 564448 225202 564460
rect 227990 564448 227996 564460
rect 225196 564420 227996 564448
rect 225196 564408 225202 564420
rect 227990 564408 227996 564420
rect 228048 564408 228054 564460
rect 260098 564408 260104 564460
rect 260156 564448 260162 564460
rect 262766 564448 262772 564460
rect 260156 564420 262772 564448
rect 260156 564408 260162 564420
rect 262766 564408 262772 564420
rect 262824 564408 262830 564460
rect 264238 564408 264244 564460
rect 264296 564448 264302 564460
rect 265342 564448 265348 564460
rect 264296 564420 265348 564448
rect 264296 564408 264302 564420
rect 265342 564408 265348 564420
rect 265400 564408 265406 564460
rect 266998 564408 267004 564460
rect 267056 564448 267062 564460
rect 268654 564448 268660 564460
rect 267056 564420 268660 564448
rect 267056 564408 267062 564420
rect 268654 564408 268660 564420
rect 268712 564408 268718 564460
rect 269758 564408 269764 564460
rect 269816 564448 269822 564460
rect 271230 564448 271236 564460
rect 269816 564420 271236 564448
rect 269816 564408 269822 564420
rect 271230 564408 271236 564420
rect 271288 564408 271294 564460
rect 278038 564408 278044 564460
rect 278096 564448 278102 564460
rect 280246 564448 280252 564460
rect 278096 564420 280252 564448
rect 278096 564408 278102 564420
rect 280246 564408 280252 564420
rect 280304 564408 280310 564460
rect 274818 563932 274824 563984
rect 274876 563972 274882 563984
rect 312630 563972 312636 563984
rect 274876 563944 312636 563972
rect 274876 563932 274882 563944
rect 312630 563932 312636 563944
rect 312688 563932 312694 563984
rect 57422 563864 57428 563916
rect 57480 563904 57486 563916
rect 87598 563904 87604 563916
rect 57480 563876 87604 563904
rect 57480 563864 57486 563876
rect 87598 563864 87604 563876
rect 87656 563864 87662 563916
rect 128354 563864 128360 563916
rect 128412 563904 128418 563916
rect 201954 563904 201960 563916
rect 128412 563876 201960 563904
rect 128412 563864 128418 563876
rect 201954 563864 201960 563876
rect 202012 563864 202018 563916
rect 226426 563864 226432 563916
rect 226484 563904 226490 563916
rect 280798 563904 280804 563916
rect 226484 563876 280804 563904
rect 226484 563864 226490 563876
rect 280798 563864 280804 563876
rect 280856 563864 280862 563916
rect 85666 563796 85672 563848
rect 85724 563836 85730 563848
rect 121822 563836 121828 563848
rect 85724 563808 121828 563836
rect 85724 563796 85730 563808
rect 121822 563796 121828 563808
rect 121880 563796 121886 563848
rect 122834 563796 122840 563848
rect 122892 563836 122898 563848
rect 201034 563836 201040 563848
rect 122892 563808 201040 563836
rect 122892 563796 122898 563808
rect 201034 563796 201040 563808
rect 201092 563796 201098 563848
rect 219250 563796 219256 563848
rect 219308 563836 219314 563848
rect 223666 563836 223672 563848
rect 219308 563808 223672 563836
rect 219308 563796 219314 563808
rect 223666 563796 223672 563808
rect 223724 563796 223730 563848
rect 255314 563796 255320 563848
rect 255372 563836 255378 563848
rect 318242 563836 318248 563848
rect 255372 563808 318248 563836
rect 255372 563796 255378 563808
rect 318242 563796 318248 563808
rect 318300 563796 318306 563848
rect 59446 563728 59452 563780
rect 59504 563768 59510 563780
rect 76006 563768 76012 563780
rect 59504 563740 76012 563768
rect 59504 563728 59510 563740
rect 76006 563728 76012 563740
rect 76064 563728 76070 563780
rect 80054 563728 80060 563780
rect 80112 563768 80118 563780
rect 123294 563768 123300 563780
rect 80112 563740 123300 563768
rect 80112 563728 80118 563740
rect 123294 563728 123300 563740
rect 123352 563728 123358 563780
rect 195974 563728 195980 563780
rect 196032 563768 196038 563780
rect 283282 563768 283288 563780
rect 196032 563740 283288 563768
rect 196032 563728 196038 563740
rect 283282 563728 283288 563740
rect 283340 563728 283346 563780
rect 63494 563660 63500 563712
rect 63552 563700 63558 563712
rect 123662 563700 123668 563712
rect 63552 563672 123668 563700
rect 63552 563660 63558 563672
rect 123662 563660 123668 563672
rect 123720 563660 123726 563712
rect 138842 563660 138848 563712
rect 138900 563700 138906 563712
rect 160186 563700 160192 563712
rect 138900 563672 160192 563700
rect 138900 563660 138906 563672
rect 160186 563660 160192 563672
rect 160244 563660 160250 563712
rect 179598 563660 179604 563712
rect 179656 563700 179662 563712
rect 281534 563700 281540 563712
rect 179656 563672 281540 563700
rect 179656 563660 179662 563672
rect 281534 563660 281540 563672
rect 281592 563660 281598 563712
rect 266354 562572 266360 562624
rect 266412 562612 266418 562624
rect 302878 562612 302884 562624
rect 266412 562584 302884 562612
rect 266412 562572 266418 562584
rect 302878 562572 302884 562584
rect 302936 562572 302942 562624
rect 120166 562504 120172 562556
rect 120224 562544 120230 562556
rect 187694 562544 187700 562556
rect 120224 562516 187700 562544
rect 120224 562504 120230 562516
rect 187694 562504 187700 562516
rect 187752 562504 187758 562556
rect 198734 562504 198740 562556
rect 198792 562544 198798 562556
rect 206462 562544 206468 562556
rect 198792 562516 206468 562544
rect 198792 562504 198798 562516
rect 206462 562504 206468 562516
rect 206520 562504 206526 562556
rect 215386 562504 215392 562556
rect 215444 562544 215450 562556
rect 282086 562544 282092 562556
rect 215444 562516 282092 562544
rect 215444 562504 215450 562516
rect 282086 562504 282092 562516
rect 282144 562504 282150 562556
rect 80146 562436 80152 562488
rect 80204 562476 80210 562488
rect 121086 562476 121092 562488
rect 80204 562448 121092 562476
rect 80204 562436 80210 562448
rect 121086 562436 121092 562448
rect 121144 562436 121150 562488
rect 126974 562436 126980 562488
rect 127032 562476 127038 562488
rect 201494 562476 201500 562488
rect 127032 562448 201500 562476
rect 127032 562436 127038 562448
rect 201494 562436 201500 562448
rect 201552 562436 201558 562488
rect 234614 562436 234620 562488
rect 234672 562476 234678 562488
rect 319714 562476 319720 562488
rect 234672 562448 319720 562476
rect 234672 562436 234678 562448
rect 319714 562436 319720 562448
rect 319772 562436 319778 562488
rect 57054 562368 57060 562420
rect 57112 562408 57118 562420
rect 110506 562408 110512 562420
rect 57112 562380 110512 562408
rect 57112 562368 57118 562380
rect 110506 562368 110512 562380
rect 110564 562368 110570 562420
rect 138750 562368 138756 562420
rect 138808 562408 138814 562420
rect 138808 562380 142154 562408
rect 138808 562368 138814 562380
rect 63586 562300 63592 562352
rect 63644 562340 63650 562352
rect 122926 562340 122932 562352
rect 63644 562312 122932 562340
rect 63644 562300 63650 562312
rect 122926 562300 122932 562312
rect 122984 562300 122990 562352
rect 139394 562300 139400 562352
rect 139452 562340 139458 562352
rect 139946 562340 139952 562352
rect 139452 562312 139952 562340
rect 139452 562300 139458 562312
rect 139946 562300 139952 562312
rect 140004 562300 140010 562352
rect 142126 562340 142154 562380
rect 184934 562368 184940 562420
rect 184992 562408 184998 562420
rect 274634 562408 274640 562420
rect 184992 562380 274640 562408
rect 184992 562368 184998 562380
rect 274634 562368 274640 562380
rect 274692 562368 274698 562420
rect 173894 562340 173900 562352
rect 142126 562312 173900 562340
rect 173894 562300 173900 562312
rect 173952 562300 173958 562352
rect 186314 562300 186320 562352
rect 186372 562340 186378 562352
rect 281994 562340 282000 562352
rect 186372 562312 282000 562340
rect 186372 562300 186378 562312
rect 281994 562300 282000 562312
rect 282052 562300 282058 562352
rect 285030 562340 285036 562352
rect 282886 562312 285036 562340
rect 281534 562232 281540 562284
rect 281592 562272 281598 562284
rect 282886 562272 282914 562312
rect 285030 562300 285036 562312
rect 285088 562300 285094 562352
rect 281592 562244 282914 562272
rect 281592 562232 281598 562244
rect 190546 561144 190552 561196
rect 190604 561184 190610 561196
rect 204990 561184 204996 561196
rect 190604 561156 204996 561184
rect 190604 561144 190610 561156
rect 204990 561144 204996 561156
rect 205048 561144 205054 561196
rect 88610 561076 88616 561128
rect 88668 561116 88674 561128
rect 103514 561116 103520 561128
rect 88668 561088 103520 561116
rect 88668 561076 88674 561088
rect 103514 561076 103520 561088
rect 103572 561076 103578 561128
rect 193214 561076 193220 561128
rect 193272 561116 193278 561128
rect 218790 561116 218796 561128
rect 193272 561088 218796 561116
rect 193272 561076 193278 561088
rect 218790 561076 218796 561088
rect 218848 561076 218854 561128
rect 59170 561008 59176 561060
rect 59228 561048 59234 561060
rect 92566 561048 92572 561060
rect 59228 561020 92572 561048
rect 59228 561008 59234 561020
rect 92566 561008 92572 561020
rect 92624 561008 92630 561060
rect 142246 561008 142252 561060
rect 142304 561048 142310 561060
rect 203242 561048 203248 561060
rect 142304 561020 203248 561048
rect 142304 561008 142310 561020
rect 203242 561008 203248 561020
rect 203300 561008 203306 561060
rect 217594 561008 217600 561060
rect 217652 561048 217658 561060
rect 231946 561048 231952 561060
rect 217652 561020 231952 561048
rect 217652 561008 217658 561020
rect 231946 561008 231952 561020
rect 232004 561008 232010 561060
rect 263594 561008 263600 561060
rect 263652 561048 263658 561060
rect 311250 561048 311256 561060
rect 263652 561020 311256 561048
rect 263652 561008 263658 561020
rect 311250 561008 311256 561020
rect 311308 561008 311314 561060
rect 70394 560940 70400 560992
rect 70452 560980 70458 560992
rect 120810 560980 120816 560992
rect 70452 560952 120816 560980
rect 70452 560940 70458 560952
rect 120810 560940 120816 560952
rect 120868 560940 120874 560992
rect 138934 560940 138940 560992
rect 138992 560980 138998 560992
rect 165706 560980 165712 560992
rect 138992 560952 165712 560980
rect 138992 560940 138998 560952
rect 165706 560940 165712 560952
rect 165764 560940 165770 560992
rect 201494 560940 201500 560992
rect 201552 560980 201558 560992
rect 283006 560980 283012 560992
rect 201552 560952 283012 560980
rect 201552 560940 201558 560952
rect 283006 560940 283012 560952
rect 283064 560940 283070 560992
rect 21358 560260 21364 560312
rect 21416 560300 21422 560312
rect 317966 560300 317972 560312
rect 21416 560272 317972 560300
rect 21416 560260 21422 560272
rect 317966 560260 317972 560272
rect 318024 560260 318030 560312
rect 266446 559784 266452 559836
rect 266504 559824 266510 559836
rect 287698 559824 287704 559836
rect 266504 559796 287704 559824
rect 266504 559784 266510 559796
rect 287698 559784 287704 559796
rect 287756 559784 287762 559836
rect 88426 559716 88432 559768
rect 88484 559756 88490 559768
rect 104894 559756 104900 559768
rect 88484 559728 104900 559756
rect 88484 559716 88490 559728
rect 104894 559716 104900 559728
rect 104952 559716 104958 559768
rect 176654 559716 176660 559768
rect 176712 559756 176718 559768
rect 213270 559756 213276 559768
rect 176712 559728 213276 559756
rect 176712 559716 176718 559728
rect 213270 559716 213276 559728
rect 213328 559716 213334 559768
rect 273254 559716 273260 559768
rect 273312 559756 273318 559768
rect 318150 559756 318156 559768
rect 273312 559728 318156 559756
rect 273312 559716 273318 559728
rect 318150 559716 318156 559728
rect 318208 559716 318214 559768
rect 129826 559648 129832 559700
rect 129884 559688 129890 559700
rect 202874 559688 202880 559700
rect 129884 559660 202880 559688
rect 129884 559648 129890 559660
rect 202874 559648 202880 559660
rect 202932 559648 202938 559700
rect 240134 559648 240140 559700
rect 240192 559688 240198 559700
rect 314010 559688 314016 559700
rect 240192 559660 314016 559688
rect 240192 559648 240198 559660
rect 314010 559648 314016 559660
rect 314068 559648 314074 559700
rect 62574 559580 62580 559632
rect 62632 559620 62638 559632
rect 104986 559620 104992 559632
rect 62632 559592 104992 559620
rect 62632 559580 62638 559592
rect 104986 559580 104992 559592
rect 105044 559580 105050 559632
rect 122926 559580 122932 559632
rect 122984 559620 122990 559632
rect 201862 559620 201868 559632
rect 122984 559592 201868 559620
rect 122984 559580 122990 559592
rect 201862 559580 201868 559592
rect 201920 559580 201926 559632
rect 233326 559580 233332 559632
rect 233384 559620 233390 559632
rect 319622 559620 319628 559632
rect 233384 559592 319628 559620
rect 233384 559580 233390 559592
rect 319622 559580 319628 559592
rect 319680 559580 319686 559632
rect 65058 559512 65064 559564
rect 65116 559552 65122 559564
rect 123110 559552 123116 559564
rect 65116 559524 123116 559552
rect 65116 559512 65122 559524
rect 123110 559512 123116 559524
rect 123168 559512 123174 559564
rect 138658 559512 138664 559564
rect 138716 559552 138722 559564
rect 168466 559552 168472 559564
rect 138716 559524 168472 559552
rect 138716 559512 138722 559524
rect 168466 559512 168472 559524
rect 168524 559512 168530 559564
rect 196066 559512 196072 559564
rect 196124 559552 196130 559564
rect 283374 559552 283380 559564
rect 196124 559524 283380 559552
rect 196124 559512 196130 559524
rect 283374 559512 283380 559524
rect 283432 559512 283438 559564
rect 219618 558424 219624 558476
rect 219676 558464 219682 558476
rect 247126 558464 247132 558476
rect 219676 558436 247132 558464
rect 219676 558424 219682 558436
rect 247126 558424 247132 558436
rect 247184 558424 247190 558476
rect 279510 558424 279516 558476
rect 279568 558464 279574 558476
rect 294598 558464 294604 558476
rect 279568 558436 294604 558464
rect 279568 558424 279574 558436
rect 294598 558424 294604 558436
rect 294656 558424 294662 558476
rect 176746 558356 176752 558408
rect 176804 558396 176810 558408
rect 225046 558396 225052 558408
rect 176804 558368 225052 558396
rect 176804 558356 176810 558368
rect 225046 558356 225052 558368
rect 225104 558356 225110 558408
rect 256694 558356 256700 558408
rect 256752 558396 256758 558408
rect 309778 558396 309784 558408
rect 256752 558368 309784 558396
rect 256752 558356 256758 558368
rect 309778 558356 309784 558368
rect 309836 558356 309842 558408
rect 57606 558288 57612 558340
rect 57664 558328 57670 558340
rect 107746 558328 107752 558340
rect 57664 558300 107752 558328
rect 57664 558288 57670 558300
rect 107746 558288 107752 558300
rect 107804 558288 107810 558340
rect 134518 558288 134524 558340
rect 134576 558328 134582 558340
rect 187878 558328 187884 558340
rect 134576 558300 187884 558328
rect 134576 558288 134582 558300
rect 187878 558288 187884 558300
rect 187936 558288 187942 558340
rect 197354 558288 197360 558340
rect 197412 558328 197418 558340
rect 209038 558328 209044 558340
rect 197412 558300 209044 558328
rect 197412 558288 197418 558300
rect 209038 558288 209044 558300
rect 209096 558288 209102 558340
rect 227806 558288 227812 558340
rect 227864 558328 227870 558340
rect 282914 558328 282920 558340
rect 227864 558300 282920 558328
rect 227864 558288 227870 558300
rect 282914 558288 282920 558300
rect 282972 558288 282978 558340
rect 70486 558220 70492 558272
rect 70544 558260 70550 558272
rect 121730 558260 121736 558272
rect 70544 558232 121736 558260
rect 70544 558220 70550 558232
rect 121730 558220 121736 558232
rect 121788 558220 121794 558272
rect 124306 558220 124312 558272
rect 124364 558260 124370 558272
rect 201218 558260 201224 558272
rect 124364 558232 201224 558260
rect 124364 558220 124370 558232
rect 201218 558220 201224 558232
rect 201276 558220 201282 558272
rect 245654 558220 245660 558272
rect 245712 558260 245718 558272
rect 307018 558260 307024 558272
rect 245712 558232 307024 558260
rect 245712 558220 245718 558232
rect 307018 558220 307024 558232
rect 307076 558220 307082 558272
rect 66346 558152 66352 558204
rect 66404 558192 66410 558204
rect 123570 558192 123576 558204
rect 66404 558164 123576 558192
rect 66404 558152 66410 558164
rect 123570 558152 123576 558164
rect 123628 558152 123634 558204
rect 137922 558152 137928 558204
rect 137980 558192 137986 558204
rect 149146 558192 149152 558204
rect 137980 558164 149152 558192
rect 137980 558152 137986 558164
rect 149146 558152 149152 558164
rect 149204 558152 149210 558204
rect 186406 558152 186412 558204
rect 186464 558192 186470 558204
rect 283098 558192 283104 558204
rect 186464 558164 283104 558192
rect 186464 558152 186470 558164
rect 283098 558152 283104 558164
rect 283156 558152 283162 558204
rect 40034 557472 40040 557524
rect 40092 557512 40098 557524
rect 317414 557512 317420 557524
rect 40092 557484 317420 557512
rect 40092 557472 40098 557484
rect 317414 557472 317420 557484
rect 317472 557472 317478 557524
rect 192110 556996 192116 557048
rect 192168 557036 192174 557048
rect 210418 557036 210424 557048
rect 192168 557008 210424 557036
rect 192168 556996 192174 557008
rect 210418 556996 210424 557008
rect 210476 556996 210482 557048
rect 188522 556928 188528 556980
rect 188580 556968 188586 556980
rect 233234 556968 233240 556980
rect 188580 556940 233240 556968
rect 188580 556928 188586 556940
rect 233234 556928 233240 556940
rect 233292 556928 233298 556980
rect 260190 556928 260196 556980
rect 260248 556968 260254 556980
rect 287882 556968 287888 556980
rect 260248 556940 287888 556968
rect 260248 556928 260254 556940
rect 287882 556928 287888 556940
rect 287940 556928 287946 556980
rect 78858 556860 78864 556912
rect 78916 556900 78922 556912
rect 115382 556900 115388 556912
rect 78916 556872 115388 556900
rect 78916 556860 78922 556872
rect 115382 556860 115388 556872
rect 115440 556860 115446 556912
rect 152642 556860 152648 556912
rect 152700 556900 152706 556912
rect 202046 556900 202052 556912
rect 152700 556872 202052 556900
rect 152700 556860 152706 556872
rect 202046 556860 202052 556872
rect 202104 556860 202110 556912
rect 229278 556860 229284 556912
rect 229336 556900 229342 556912
rect 281258 556900 281264 556912
rect 229336 556872 281264 556900
rect 229336 556860 229342 556872
rect 281258 556860 281264 556872
rect 281316 556860 281322 556912
rect 58894 556792 58900 556844
rect 58952 556832 58958 556844
rect 102502 556832 102508 556844
rect 58952 556804 102508 556832
rect 58952 556792 58958 556804
rect 102502 556792 102508 556804
rect 102560 556792 102566 556844
rect 140498 556792 140504 556844
rect 140556 556832 140562 556844
rect 197998 556832 198004 556844
rect 140556 556804 198004 556832
rect 140556 556792 140562 556804
rect 197998 556792 198004 556804
rect 198056 556792 198062 556844
rect 245102 556792 245108 556844
rect 245160 556832 245166 556844
rect 315298 556832 315304 556844
rect 245160 556804 315304 556832
rect 245160 556792 245166 556804
rect 315298 556792 315304 556804
rect 315356 556792 315362 556844
rect 124214 556452 124220 556504
rect 124272 556492 124278 556504
rect 125410 556492 125416 556504
rect 124272 556464 125416 556492
rect 124272 556452 124278 556464
rect 125410 556452 125416 556464
rect 125468 556452 125474 556504
rect 126974 556316 126980 556368
rect 127032 556356 127038 556368
rect 128262 556356 128268 556368
rect 127032 556328 128268 556356
rect 127032 556316 127038 556328
rect 128262 556316 128268 556328
rect 128320 556316 128326 556368
rect 217778 556180 217784 556232
rect 217836 556220 217842 556232
rect 218606 556220 218612 556232
rect 217836 556192 218612 556220
rect 217836 556180 217842 556192
rect 218606 556180 218612 556192
rect 218664 556180 218670 556232
rect 219618 556044 219624 556096
rect 219676 556084 219682 556096
rect 220722 556084 220728 556096
rect 219676 556056 220728 556084
rect 219676 556044 219682 556056
rect 220722 556044 220728 556056
rect 220780 556044 220786 556096
rect 222194 555772 222200 555824
rect 222252 555812 222258 555824
rect 222838 555812 222844 555824
rect 222252 555784 222844 555812
rect 222252 555772 222258 555784
rect 222838 555772 222844 555784
rect 222896 555772 222902 555824
rect 193490 555636 193496 555688
rect 193548 555676 193554 555688
rect 215938 555676 215944 555688
rect 193548 555648 215944 555676
rect 193548 555636 193554 555648
rect 215938 555636 215944 555648
rect 215996 555636 216002 555688
rect 217870 555636 217876 555688
rect 217928 555676 217934 555688
rect 260098 555676 260104 555688
rect 217928 555648 260104 555676
rect 217928 555636 217934 555648
rect 260098 555636 260104 555648
rect 260156 555636 260162 555688
rect 94590 555568 94596 555620
rect 94648 555608 94654 555620
rect 122006 555608 122012 555620
rect 94648 555580 122012 555608
rect 94648 555568 94654 555580
rect 122006 555568 122012 555580
rect 122064 555568 122070 555620
rect 142338 555568 142344 555620
rect 142396 555608 142402 555620
rect 167730 555608 167736 555620
rect 142396 555580 167736 555608
rect 142396 555568 142402 555580
rect 167730 555568 167736 555580
rect 167788 555568 167794 555620
rect 178494 555568 178500 555620
rect 178552 555608 178558 555620
rect 206554 555608 206560 555620
rect 178552 555580 206560 555608
rect 178552 555568 178558 555580
rect 206554 555568 206560 555580
rect 206612 555568 206618 555620
rect 250070 555568 250076 555620
rect 250128 555608 250134 555620
rect 295978 555608 295984 555620
rect 250128 555580 295984 555608
rect 250128 555568 250134 555580
rect 295978 555568 295984 555580
rect 296036 555568 296042 555620
rect 58434 555500 58440 555552
rect 58492 555540 58498 555552
rect 103238 555540 103244 555552
rect 58492 555512 103244 555540
rect 58492 555500 58498 555512
rect 103238 555500 103244 555512
rect 103296 555500 103302 555552
rect 144086 555500 144092 555552
rect 144144 555540 144150 555552
rect 202230 555540 202236 555552
rect 144144 555512 202236 555540
rect 144144 555500 144150 555512
rect 202230 555500 202236 555512
rect 202288 555500 202294 555552
rect 208486 555500 208492 555552
rect 208544 555540 208550 555552
rect 235994 555540 236000 555552
rect 208544 555512 236000 555540
rect 208544 555500 208550 555512
rect 235994 555500 236000 555512
rect 236052 555500 236058 555552
rect 236086 555500 236092 555552
rect 236144 555540 236150 555552
rect 283190 555540 283196 555552
rect 236144 555512 283196 555540
rect 236144 555500 236150 555512
rect 283190 555500 283196 555512
rect 283248 555500 283254 555552
rect 63126 555432 63132 555484
rect 63184 555472 63190 555484
rect 110598 555472 110604 555484
rect 63184 555444 110604 555472
rect 63184 555432 63190 555444
rect 110598 555432 110604 555444
rect 110656 555432 110662 555484
rect 121822 555432 121828 555484
rect 121880 555472 121886 555484
rect 201126 555472 201132 555484
rect 121880 555444 201132 555472
rect 121880 555432 121886 555444
rect 201126 555432 201132 555444
rect 201184 555432 201190 555484
rect 205634 555432 205640 555484
rect 205692 555472 205698 555484
rect 264238 555472 264244 555484
rect 205692 555444 264244 555472
rect 205692 555432 205698 555444
rect 264238 555432 264244 555444
rect 264296 555432 264302 555484
rect 270126 555432 270132 555484
rect 270184 555472 270190 555484
rect 286318 555472 286324 555484
rect 270184 555444 286324 555472
rect 270184 555432 270190 555444
rect 286318 555432 286324 555444
rect 286376 555432 286382 555484
rect 58618 554208 58624 554260
rect 58676 554248 58682 554260
rect 74534 554248 74540 554260
rect 58676 554220 74540 554248
rect 58676 554208 58682 554220
rect 74534 554208 74540 554220
rect 74592 554208 74598 554260
rect 189902 554208 189908 554260
rect 189960 554248 189966 554260
rect 217318 554248 217324 554260
rect 189960 554220 217324 554248
rect 189960 554208 189966 554220
rect 217318 554208 217324 554220
rect 217376 554208 217382 554260
rect 73154 554140 73160 554192
rect 73212 554180 73218 554192
rect 106918 554180 106924 554192
rect 73212 554152 106924 554180
rect 73212 554140 73218 554152
rect 106918 554140 106924 554152
rect 106976 554140 106982 554192
rect 157242 554140 157248 554192
rect 157300 554180 157306 554192
rect 203058 554180 203064 554192
rect 157300 554152 203064 554180
rect 157300 554140 157306 554152
rect 203058 554140 203064 554152
rect 203116 554140 203122 554192
rect 250806 554140 250812 554192
rect 250864 554180 250870 554192
rect 319530 554180 319536 554192
rect 250864 554152 319536 554180
rect 250864 554140 250870 554152
rect 319530 554140 319536 554152
rect 319588 554140 319594 554192
rect 72418 554072 72424 554124
rect 72476 554112 72482 554124
rect 109678 554112 109684 554124
rect 72476 554084 109684 554112
rect 72476 554072 72482 554084
rect 109678 554072 109684 554084
rect 109736 554072 109742 554124
rect 136910 554072 136916 554124
rect 136968 554112 136974 554124
rect 202322 554112 202328 554124
rect 136968 554084 202328 554112
rect 136968 554072 136974 554084
rect 202322 554072 202328 554084
rect 202380 554072 202386 554124
rect 206370 554072 206376 554124
rect 206428 554112 206434 554124
rect 241514 554112 241520 554124
rect 206428 554084 241520 554112
rect 206428 554072 206434 554084
rect 241514 554072 241520 554084
rect 241572 554072 241578 554124
rect 242894 554072 242900 554124
rect 242952 554112 242958 554124
rect 316862 554112 316868 554124
rect 242952 554084 316868 554112
rect 242952 554072 242958 554084
rect 316862 554072 316868 554084
rect 316920 554072 316926 554124
rect 69566 554004 69572 554056
rect 69624 554044 69630 554056
rect 114554 554044 114560 554056
rect 69624 554016 114560 554044
rect 69624 554004 69630 554016
rect 114554 554004 114560 554016
rect 114612 554004 114618 554056
rect 179138 554004 179144 554056
rect 179196 554044 179202 554056
rect 269758 554044 269764 554056
rect 179196 554016 269764 554044
rect 179196 554004 179202 554016
rect 269758 554004 269764 554016
rect 269816 554004 269822 554056
rect 57330 552916 57336 552968
rect 57388 552956 57394 552968
rect 123202 552956 123208 552968
rect 57388 552928 64874 552956
rect 57388 552916 57394 552928
rect 59538 552848 59544 552900
rect 59596 552848 59602 552900
rect 59556 552684 59584 552848
rect 64846 552820 64874 552928
rect 122806 552928 123208 552956
rect 70486 552848 70492 552900
rect 70544 552888 70550 552900
rect 71682 552888 71688 552900
rect 70544 552860 71688 552888
rect 70544 552848 70550 552860
rect 71682 552848 71688 552860
rect 71740 552848 71746 552900
rect 81710 552820 81716 552832
rect 64846 552792 81716 552820
rect 81710 552780 81716 552792
rect 81768 552780 81774 552832
rect 86954 552780 86960 552832
rect 87012 552820 87018 552832
rect 88150 552820 88156 552832
rect 87012 552792 88156 552820
rect 87012 552780 87018 552792
rect 88150 552780 88156 552792
rect 88208 552780 88214 552832
rect 88426 552780 88432 552832
rect 88484 552820 88490 552832
rect 89622 552820 89628 552832
rect 88484 552792 89628 552820
rect 88484 552780 88490 552792
rect 89622 552780 89628 552792
rect 89680 552780 89686 552832
rect 98086 552780 98092 552832
rect 98144 552820 98150 552832
rect 122806 552820 122834 552928
rect 123202 552916 123208 552928
rect 123260 552916 123266 552968
rect 216030 552956 216036 552968
rect 200086 552928 216036 552956
rect 122926 552848 122932 552900
rect 122984 552888 122990 552900
rect 124030 552888 124036 552900
rect 122984 552860 124036 552888
rect 122984 552848 122990 552860
rect 124030 552848 124036 552860
rect 124088 552848 124094 552900
rect 184934 552848 184940 552900
rect 184992 552888 184998 552900
rect 200086 552888 200114 552928
rect 216030 552916 216036 552928
rect 216088 552916 216094 552968
rect 251542 552916 251548 552968
rect 251600 552956 251606 552968
rect 251600 552928 258074 552956
rect 251600 552916 251606 552928
rect 184992 552860 200114 552888
rect 184992 552848 184998 552860
rect 202138 552848 202144 552900
rect 202196 552848 202202 552900
rect 210694 552848 210700 552900
rect 210752 552888 210758 552900
rect 210752 552860 219434 552888
rect 210752 552848 210758 552860
rect 98144 552792 122834 552820
rect 98144 552780 98150 552792
rect 139026 552780 139032 552832
rect 139084 552820 139090 552832
rect 202156 552820 202184 552848
rect 139084 552792 202184 552820
rect 139084 552780 139090 552792
rect 208394 552780 208400 552832
rect 208452 552820 208458 552832
rect 209222 552820 209228 552832
rect 208452 552792 209228 552820
rect 208452 552780 208458 552792
rect 209222 552780 209228 552792
rect 209280 552780 209286 552832
rect 212534 552780 212540 552832
rect 212592 552820 212598 552832
rect 213546 552820 213552 552832
rect 212592 552792 213552 552820
rect 212592 552780 212598 552792
rect 213546 552780 213552 552792
rect 213604 552780 213610 552832
rect 213914 552780 213920 552832
rect 213972 552820 213978 552832
rect 215018 552820 215024 552832
rect 213972 552792 215024 552820
rect 213972 552780 213978 552792
rect 215018 552780 215024 552792
rect 215076 552780 215082 552832
rect 219406 552820 219434 552860
rect 255314 552848 255320 552900
rect 255372 552888 255378 552900
rect 256510 552888 256516 552900
rect 255372 552860 256516 552888
rect 255372 552848 255378 552860
rect 256510 552848 256516 552860
rect 256568 552848 256574 552900
rect 258046 552888 258074 552928
rect 259454 552916 259460 552968
rect 259512 552956 259518 552968
rect 311158 552956 311164 552968
rect 259512 552928 311164 552956
rect 259512 552916 259518 552928
rect 311158 552916 311164 552928
rect 311216 552916 311222 552968
rect 316678 552888 316684 552900
rect 258046 552860 316684 552888
rect 316678 552848 316684 552860
rect 316736 552848 316742 552900
rect 280982 552820 280988 552832
rect 219406 552792 280988 552820
rect 280982 552780 280988 552792
rect 281040 552780 281046 552832
rect 67634 552712 67640 552764
rect 67692 552752 67698 552764
rect 68830 552752 68836 552764
rect 67692 552724 68836 552752
rect 67692 552712 67698 552724
rect 68830 552712 68836 552724
rect 68888 552712 68894 552764
rect 69014 552712 69020 552764
rect 69072 552752 69078 552764
rect 70302 552752 70308 552764
rect 69072 552724 70308 552752
rect 69072 552712 69078 552724
rect 70302 552712 70308 552724
rect 70360 552712 70366 552764
rect 75914 552712 75920 552764
rect 75972 552752 75978 552764
rect 76742 552752 76748 552764
rect 75972 552724 76748 552752
rect 75972 552712 75978 552724
rect 76742 552712 76748 552724
rect 76800 552712 76806 552764
rect 82446 552712 82452 552764
rect 82504 552752 82510 552764
rect 116578 552752 116584 552764
rect 82504 552724 116584 552752
rect 82504 552712 82510 552724
rect 116578 552712 116584 552724
rect 116636 552712 116642 552764
rect 125594 552712 125600 552764
rect 125652 552752 125658 552764
rect 126882 552752 126888 552764
rect 125652 552724 126888 552752
rect 125652 552712 125658 552724
rect 126882 552712 126888 552724
rect 126940 552712 126946 552764
rect 129734 552712 129740 552764
rect 129792 552752 129798 552764
rect 130470 552752 130476 552764
rect 129792 552724 130476 552752
rect 129792 552712 129798 552724
rect 130470 552712 130476 552724
rect 130528 552712 130534 552764
rect 142154 552712 142160 552764
rect 142212 552752 142218 552764
rect 143350 552752 143356 552764
rect 142212 552724 143356 552752
rect 142212 552712 142218 552724
rect 143350 552712 143356 552724
rect 143408 552712 143414 552764
rect 143534 552712 143540 552764
rect 143592 552752 143598 552764
rect 144730 552752 144736 552764
rect 143592 552724 144736 552752
rect 143592 552712 143598 552724
rect 144730 552712 144736 552724
rect 144788 552712 144794 552764
rect 154574 552712 154580 552764
rect 154632 552752 154638 552764
rect 155494 552752 155500 552764
rect 154632 552724 155500 552752
rect 154632 552712 154638 552724
rect 155494 552712 155500 552724
rect 155552 552712 155558 552764
rect 160094 552712 160100 552764
rect 160152 552752 160158 552764
rect 161290 552752 161296 552764
rect 160152 552724 161296 552752
rect 160152 552712 160158 552724
rect 161290 552712 161296 552724
rect 161348 552712 161354 552764
rect 164326 552712 164332 552764
rect 164384 552752 164390 552764
rect 165522 552752 165528 552764
rect 164384 552724 165528 552752
rect 164384 552712 164390 552724
rect 165522 552712 165528 552724
rect 165580 552712 165586 552764
rect 180794 552712 180800 552764
rect 180852 552752 180858 552764
rect 181990 552752 181996 552764
rect 180852 552724 181996 552752
rect 180852 552712 180858 552724
rect 181990 552712 181996 552724
rect 182048 552712 182054 552764
rect 189166 552712 189172 552764
rect 189224 552752 189230 552764
rect 266998 552752 267004 552764
rect 189224 552724 267004 552752
rect 189224 552712 189230 552724
rect 266998 552712 267004 552724
rect 267056 552712 267062 552764
rect 273254 552712 273260 552764
rect 273312 552752 273318 552764
rect 274450 552752 274456 552764
rect 273312 552724 274456 552752
rect 273312 552712 273318 552724
rect 274450 552712 274456 552724
rect 274508 552712 274514 552764
rect 293954 552712 293960 552764
rect 294012 552752 294018 552764
rect 295242 552752 295248 552764
rect 294012 552724 295248 552752
rect 294012 552712 294018 552724
rect 295242 552712 295248 552724
rect 295300 552712 295306 552764
rect 101030 552684 101036 552696
rect 59556 552656 101036 552684
rect 101030 552644 101036 552656
rect 101088 552644 101094 552696
rect 106274 552644 106280 552696
rect 106332 552684 106338 552696
rect 107562 552684 107568 552696
rect 106332 552656 107568 552684
rect 106332 552644 106338 552656
rect 107562 552644 107568 552656
rect 107620 552644 107626 552696
rect 127618 552644 127624 552696
rect 127676 552684 127682 552696
rect 194686 552684 194692 552696
rect 127676 552656 194692 552684
rect 127676 552644 127682 552656
rect 194686 552644 194692 552656
rect 194744 552644 194750 552696
rect 198550 552644 198556 552696
rect 198608 552684 198614 552696
rect 278038 552684 278044 552696
rect 198608 552656 278044 552684
rect 198608 552644 198614 552656
rect 278038 552644 278044 552656
rect 278096 552644 278102 552696
rect 238662 552576 238668 552628
rect 238720 552616 238726 552628
rect 318518 552616 318524 552628
rect 238720 552588 318524 552616
rect 238720 552576 238726 552588
rect 318518 552576 318524 552588
rect 318576 552576 318582 552628
rect 256694 552508 256700 552560
rect 256752 552548 256758 552560
rect 257982 552548 257988 552560
rect 256752 552520 257988 552548
rect 256752 552508 256758 552520
rect 257982 552508 257988 552520
rect 258040 552508 258046 552560
rect 293126 552508 293132 552560
rect 293184 552548 293190 552560
rect 312906 552548 312912 552560
rect 293184 552520 312912 552548
rect 293184 552508 293190 552520
rect 312906 552508 312912 552520
rect 312964 552508 312970 552560
rect 289538 552440 289544 552492
rect 289596 552480 289602 552492
rect 312722 552480 312728 552492
rect 289596 552452 312728 552480
rect 289596 552440 289602 552452
rect 312722 552440 312728 552452
rect 312780 552440 312786 552492
rect 285950 552372 285956 552424
rect 286008 552412 286014 552424
rect 312998 552412 313004 552424
rect 286008 552384 313004 552412
rect 286008 552372 286014 552384
rect 312998 552372 313004 552384
rect 313056 552372 313062 552424
rect 283098 552304 283104 552356
rect 283156 552344 283162 552356
rect 315390 552344 315396 552356
rect 283156 552316 315396 552344
rect 283156 552304 283162 552316
rect 315390 552304 315396 552316
rect 315448 552304 315454 552356
rect 284110 552236 284116 552288
rect 284168 552276 284174 552288
rect 316862 552276 316868 552288
rect 284168 552248 316868 552276
rect 284168 552236 284174 552248
rect 316862 552236 316868 552248
rect 316920 552236 316926 552288
rect 242250 552168 242256 552220
rect 242308 552208 242314 552220
rect 315298 552208 315304 552220
rect 242308 552180 315304 552208
rect 242308 552168 242314 552180
rect 315298 552168 315304 552180
rect 315356 552168 315362 552220
rect 237926 552100 237932 552152
rect 237984 552140 237990 552152
rect 318426 552140 318432 552152
rect 237984 552112 318432 552140
rect 237984 552100 237990 552112
rect 318426 552100 318432 552112
rect 318484 552100 318490 552152
rect 283742 552032 283748 552084
rect 283800 552072 283806 552084
rect 287790 552072 287796 552084
rect 283800 552044 287796 552072
rect 283800 552032 283806 552044
rect 287790 552032 287796 552044
rect 287848 552032 287854 552084
rect 293770 552032 293776 552084
rect 293828 552072 293834 552084
rect 312630 552072 312636 552084
rect 293828 552044 312636 552072
rect 293828 552032 293834 552044
rect 312630 552032 312636 552044
rect 312688 552032 312694 552084
rect 137738 551964 137744 552016
rect 137796 552004 137802 552016
rect 139762 552004 139768 552016
rect 137796 551976 139768 552004
rect 137796 551964 137802 551976
rect 139762 551964 139768 551976
rect 139820 551964 139826 552016
rect 171318 551420 171324 551472
rect 171376 551460 171382 551472
rect 203426 551460 203432 551472
rect 171376 551432 203432 551460
rect 171376 551420 171382 551432
rect 203426 551420 203432 551432
rect 203484 551420 203490 551472
rect 252278 551420 252284 551472
rect 252336 551460 252342 551472
rect 318058 551460 318064 551472
rect 252336 551432 318064 551460
rect 252336 551420 252342 551432
rect 318058 551420 318064 551432
rect 318116 551420 318122 551472
rect 137830 551352 137836 551404
rect 137888 551392 137894 551404
rect 149054 551392 149060 551404
rect 137888 551364 149060 551392
rect 137888 551352 137894 551364
rect 149054 551352 149060 551364
rect 149112 551352 149118 551404
rect 168374 551352 168380 551404
rect 168432 551392 168438 551404
rect 200758 551392 200764 551404
rect 168432 551364 200764 551392
rect 168432 551352 168438 551364
rect 200758 551352 200764 551364
rect 200816 551352 200822 551404
rect 219158 551352 219164 551404
rect 219216 551392 219222 551404
rect 227162 551392 227168 551404
rect 219216 551364 227168 551392
rect 219216 551352 219222 551364
rect 227162 551352 227168 551364
rect 227220 551352 227226 551404
rect 271598 551352 271604 551404
rect 271656 551392 271662 551404
rect 317966 551392 317972 551404
rect 271656 551364 317972 551392
rect 271656 551352 271662 551364
rect 317966 551352 317972 551364
rect 318024 551352 318030 551404
rect 57698 551284 57704 551336
rect 57756 551324 57762 551336
rect 89714 551324 89720 551336
rect 57756 551296 89720 551324
rect 57756 551284 57762 551296
rect 89714 551284 89720 551296
rect 89772 551284 89778 551336
rect 120442 551284 120448 551336
rect 120500 551324 120506 551336
rect 129090 551324 129096 551336
rect 120500 551296 129096 551324
rect 120500 551284 120506 551296
rect 129090 551284 129096 551296
rect 129148 551284 129154 551336
rect 139394 551284 139400 551336
rect 139452 551324 139458 551336
rect 163406 551324 163412 551336
rect 139452 551296 163412 551324
rect 139452 551284 139458 551296
rect 163406 551284 163412 551296
rect 163464 551284 163470 551336
rect 184198 551284 184204 551336
rect 184256 551324 184262 551336
rect 281626 551324 281632 551336
rect 184256 551296 281632 551324
rect 184256 551284 184262 551296
rect 281626 551284 281632 551296
rect 281684 551284 281690 551336
rect 285214 551284 285220 551336
rect 285272 551324 285278 551336
rect 292482 551324 292488 551336
rect 285272 551296 292488 551324
rect 285272 551284 285278 551296
rect 292482 551284 292488 551296
rect 292540 551284 292546 551336
rect 244366 551216 244372 551268
rect 244424 551256 244430 551268
rect 318242 551256 318248 551268
rect 244424 551228 318248 551256
rect 244424 551216 244430 551228
rect 318242 551216 318248 551228
rect 318300 551216 318306 551268
rect 287330 551148 287336 551200
rect 287388 551188 287394 551200
rect 313090 551188 313096 551200
rect 287388 551160 313096 551188
rect 287388 551148 287394 551160
rect 313090 551148 313096 551160
rect 313148 551148 313154 551200
rect 207106 551080 207112 551132
rect 207164 551120 207170 551132
rect 210510 551120 210516 551132
rect 207164 551092 210516 551120
rect 207164 551080 207170 551092
rect 210510 551080 210516 551092
rect 210568 551080 210574 551132
rect 291654 551080 291660 551132
rect 291712 551120 291718 551132
rect 292390 551120 292396 551132
rect 291712 551092 292396 551120
rect 291712 551080 291718 551092
rect 292390 551080 292396 551092
rect 292448 551080 292454 551132
rect 292482 551080 292488 551132
rect 292540 551120 292546 551132
rect 312814 551120 312820 551132
rect 292540 551092 312820 551120
rect 292540 551080 292546 551092
rect 312814 551080 312820 551092
rect 312872 551080 312878 551132
rect 273070 551012 273076 551064
rect 273128 551052 273134 551064
rect 302878 551052 302884 551064
rect 273128 551024 302884 551052
rect 273128 551012 273134 551024
rect 302878 551012 302884 551024
rect 302936 551012 302942 551064
rect 272334 550944 272340 550996
rect 272392 550984 272398 550996
rect 318334 550984 318340 550996
rect 272392 550956 318340 550984
rect 272392 550944 272398 550956
rect 318334 550944 318340 550956
rect 318392 550944 318398 550996
rect 263042 550876 263048 550928
rect 263100 550916 263106 550928
rect 314010 550916 314016 550928
rect 263100 550888 314016 550916
rect 263100 550876 263106 550888
rect 314010 550876 314016 550888
rect 314068 550876 314074 550928
rect 264422 550808 264428 550860
rect 264480 550848 264486 550860
rect 318150 550848 318156 550860
rect 264480 550820 318156 550848
rect 264480 550808 264486 550820
rect 318150 550808 318156 550820
rect 318208 550808 318214 550860
rect 255866 550740 255872 550792
rect 255924 550780 255930 550792
rect 316678 550780 316684 550792
rect 255924 550752 316684 550780
rect 255924 550740 255930 550752
rect 316678 550740 316684 550752
rect 316736 550740 316742 550792
rect 291194 550672 291200 550724
rect 291252 550712 291258 550724
rect 292390 550712 292396 550724
rect 291252 550684 292396 550712
rect 291252 550672 291258 550684
rect 292390 550672 292396 550684
rect 292448 550672 292454 550724
rect 292482 550672 292488 550724
rect 292540 550712 292546 550724
rect 309778 550712 309784 550724
rect 292540 550684 309784 550712
rect 292540 550672 292546 550684
rect 309778 550672 309784 550684
rect 309836 550672 309842 550724
rect 278774 550604 278780 550656
rect 278832 550644 278838 550656
rect 301406 550644 301412 550656
rect 278832 550616 301412 550644
rect 278832 550604 278838 550616
rect 301406 550604 301412 550616
rect 301464 550604 301470 550656
rect 84838 550536 84844 550588
rect 84896 550576 84902 550588
rect 86770 550576 86776 550588
rect 84896 550548 86776 550576
rect 84896 550536 84902 550548
rect 86770 550536 86776 550548
rect 86828 550536 86834 550588
rect 87598 550536 87604 550588
rect 87656 550576 87662 550588
rect 91002 550576 91008 550588
rect 87656 550548 91008 550576
rect 87656 550536 87662 550548
rect 91002 550536 91008 550548
rect 91060 550536 91066 550588
rect 108298 550536 108304 550588
rect 108356 550576 108362 550588
rect 111794 550576 111800 550588
rect 108356 550548 111800 550576
rect 108356 550536 108362 550548
rect 111794 550536 111800 550548
rect 111852 550536 111858 550588
rect 115198 550536 115204 550588
rect 115256 550576 115262 550588
rect 116118 550576 116124 550588
rect 115256 550548 116124 550576
rect 115256 550536 115262 550548
rect 116118 550536 116124 550548
rect 116176 550536 116182 550588
rect 135438 550536 135444 550588
rect 135496 550576 135502 550588
rect 137278 550576 137284 550588
rect 135496 550548 137284 550576
rect 135496 550536 135502 550548
rect 137278 550536 137284 550548
rect 137336 550536 137342 550588
rect 154114 550536 154120 550588
rect 154172 550576 154178 550588
rect 157242 550576 157248 550588
rect 154172 550548 157248 550576
rect 154172 550536 154178 550548
rect 157242 550536 157248 550548
rect 157300 550536 157306 550588
rect 165614 550536 165620 550588
rect 165672 550576 165678 550588
rect 169846 550576 169852 550588
rect 165672 550548 169852 550576
rect 165672 550536 165678 550548
rect 169846 550536 169852 550548
rect 169904 550536 169910 550588
rect 174170 550536 174176 550588
rect 174228 550576 174234 550588
rect 179506 550576 179512 550588
rect 174228 550548 179512 550576
rect 174228 550536 174234 550548
rect 179506 550536 179512 550548
rect 179564 550536 179570 550588
rect 201402 550536 201408 550588
rect 201460 550576 201466 550588
rect 206278 550576 206284 550588
rect 201460 550548 206284 550576
rect 201460 550536 201466 550548
rect 206278 550536 206284 550548
rect 206336 550536 206342 550588
rect 217502 550536 217508 550588
rect 217560 550576 217566 550588
rect 219250 550576 219256 550588
rect 217560 550548 219256 550576
rect 217560 550536 217566 550548
rect 219250 550536 219256 550548
rect 219308 550536 219314 550588
rect 219526 550536 219532 550588
rect 219584 550576 219590 550588
rect 221458 550576 221464 550588
rect 219584 550548 221464 550576
rect 219584 550536 219590 550548
rect 221458 550536 221464 550548
rect 221516 550536 221522 550588
rect 222286 550536 222292 550588
rect 222344 550576 222350 550588
rect 225782 550576 225788 550588
rect 222344 550548 225788 550576
rect 222344 550536 222350 550548
rect 225782 550536 225788 550548
rect 225840 550536 225846 550588
rect 105538 550468 105544 550520
rect 105596 550508 105602 550520
rect 108942 550508 108948 550520
rect 105596 550480 108948 550508
rect 105596 550468 105602 550480
rect 108942 550468 108948 550480
rect 109000 550468 109006 550520
rect 134978 550468 134984 550520
rect 135036 550508 135042 550520
rect 146938 550508 146944 550520
rect 135036 550480 146944 550508
rect 135036 550468 135042 550480
rect 146938 550468 146944 550480
rect 146996 550468 147002 550520
rect 162670 550468 162676 550520
rect 162728 550508 162734 550520
rect 168466 550508 168472 550520
rect 162728 550480 168472 550508
rect 162728 550468 162734 550480
rect 168466 550468 168472 550480
rect 168524 550468 168530 550520
rect 202782 550468 202788 550520
rect 202840 550508 202846 550520
rect 208486 550508 208492 550520
rect 202840 550480 208492 550508
rect 202840 550468 202846 550480
rect 208486 550468 208492 550480
rect 208544 550468 208550 550520
rect 55122 550400 55128 550452
rect 55180 550440 55186 550452
rect 67358 550440 67364 550452
rect 55180 550412 67364 550440
rect 55180 550400 55186 550412
rect 67358 550400 67364 550412
rect 67416 550400 67422 550452
rect 91186 550400 91192 550452
rect 91244 550440 91250 550452
rect 96798 550440 96804 550452
rect 91244 550412 96804 550440
rect 91244 550400 91250 550412
rect 96798 550400 96804 550412
rect 96856 550400 96862 550452
rect 139854 550400 139860 550452
rect 139912 550440 139918 550452
rect 153378 550440 153384 550452
rect 139912 550412 153384 550440
rect 139912 550400 139918 550412
rect 153378 550400 153384 550412
rect 153436 550400 153442 550452
rect 164878 550400 164884 550452
rect 164936 550440 164942 550452
rect 173434 550440 173440 550452
rect 164936 550412 173440 550440
rect 164936 550400 164942 550412
rect 173434 550400 173440 550412
rect 173492 550400 173498 550452
rect 55030 550332 55036 550384
rect 55088 550372 55094 550384
rect 88886 550372 88892 550384
rect 55088 550344 88892 550372
rect 55088 550332 55094 550344
rect 88886 550332 88892 550344
rect 88944 550332 88950 550384
rect 89714 550332 89720 550384
rect 89772 550372 89778 550384
rect 117590 550372 117596 550384
rect 89772 550344 117596 550372
rect 89772 550332 89778 550344
rect 117590 550332 117596 550344
rect 117648 550332 117654 550384
rect 135162 550332 135168 550384
rect 135220 550372 135226 550384
rect 151262 550372 151268 550384
rect 135220 550344 151268 550372
rect 135220 550332 135226 550344
rect 151262 550332 151268 550344
rect 151320 550332 151326 550384
rect 159358 550332 159364 550384
rect 159416 550372 159422 550384
rect 166994 550372 167000 550384
rect 159416 550344 167000 550372
rect 159416 550332 159422 550344
rect 166994 550332 167000 550344
rect 167052 550332 167058 550384
rect 57790 550264 57796 550316
rect 57848 550304 57854 550316
rect 93210 550304 93216 550316
rect 57848 550276 93216 550304
rect 57848 550264 57854 550276
rect 93210 550264 93216 550276
rect 93268 550264 93274 550316
rect 96062 550264 96068 550316
rect 96120 550304 96126 550316
rect 98086 550304 98092 550316
rect 96120 550276 98092 550304
rect 96120 550264 96126 550276
rect 98086 550264 98092 550276
rect 98144 550264 98150 550316
rect 118970 550264 118976 550316
rect 119028 550304 119034 550316
rect 126238 550304 126244 550316
rect 119028 550276 126244 550304
rect 119028 550264 119034 550276
rect 126238 550264 126244 550276
rect 126296 550264 126302 550316
rect 135070 550264 135076 550316
rect 135128 550304 135134 550316
rect 157702 550304 157708 550316
rect 135128 550276 157708 550304
rect 135128 550264 135134 550276
rect 157702 550264 157708 550276
rect 157760 550264 157766 550316
rect 164142 550264 164148 550316
rect 164200 550304 164206 550316
rect 173158 550304 173164 550316
rect 164200 550276 173164 550304
rect 164200 550264 164206 550276
rect 173158 550264 173164 550276
rect 173216 550264 173222 550316
rect 199930 550264 199936 550316
rect 199988 550304 199994 550316
rect 205082 550304 205088 550316
rect 199988 550276 205088 550304
rect 199988 550264 199994 550276
rect 205082 550264 205088 550276
rect 205140 550264 205146 550316
rect 262306 550264 262312 550316
rect 262364 550304 262370 550316
rect 300486 550304 300492 550316
rect 262364 550276 300492 550304
rect 262364 550264 262370 550276
rect 300486 550264 300492 550276
rect 300544 550264 300550 550316
rect 60366 550196 60372 550248
rect 60424 550236 60430 550248
rect 95326 550236 95332 550248
rect 60424 550208 95332 550236
rect 60424 550196 60430 550208
rect 95326 550196 95332 550208
rect 95384 550196 95390 550248
rect 114002 550196 114008 550248
rect 114060 550236 114066 550248
rect 127066 550236 127072 550248
rect 114060 550208 127072 550236
rect 114060 550196 114066 550208
rect 127066 550196 127072 550208
rect 127124 550196 127130 550248
rect 138290 550196 138296 550248
rect 138348 550236 138354 550248
rect 157978 550236 157984 550248
rect 138348 550208 157984 550236
rect 138348 550196 138354 550208
rect 157978 550196 157984 550208
rect 158036 550196 158042 550248
rect 160738 550196 160744 550248
rect 160796 550236 160802 550248
rect 172698 550236 172704 550248
rect 160796 550208 172704 550236
rect 160796 550196 160802 550208
rect 172698 550196 172704 550208
rect 172756 550196 172762 550248
rect 257246 550196 257252 550248
rect 257304 550236 257310 550248
rect 301958 550236 301964 550248
rect 257304 550208 301964 550236
rect 257304 550196 257310 550208
rect 301958 550196 301964 550208
rect 302016 550196 302022 550248
rect 56502 550128 56508 550180
rect 56560 550168 56566 550180
rect 83918 550168 83924 550180
rect 56560 550140 83924 550168
rect 56560 550128 56566 550140
rect 83918 550128 83924 550140
rect 83976 550128 83982 550180
rect 85298 550128 85304 550180
rect 85356 550168 85362 550180
rect 120902 550168 120908 550180
rect 85356 550140 120908 550168
rect 85356 550128 85362 550140
rect 120902 550128 120908 550140
rect 120960 550128 120966 550180
rect 137922 550128 137928 550180
rect 137980 550168 137986 550180
rect 156966 550168 156972 550180
rect 137980 550140 156972 550168
rect 137980 550128 137986 550140
rect 156966 550128 156972 550140
rect 157024 550128 157030 550180
rect 158346 550128 158352 550180
rect 158404 550168 158410 550180
rect 182818 550168 182824 550180
rect 158404 550140 182824 550168
rect 158404 550128 158410 550140
rect 182818 550128 182824 550140
rect 182876 550128 182882 550180
rect 195606 550128 195612 550180
rect 195664 550168 195670 550180
rect 206462 550168 206468 550180
rect 195664 550140 206468 550168
rect 195664 550128 195670 550140
rect 206462 550128 206468 550140
rect 206520 550128 206526 550180
rect 270862 550128 270868 550180
rect 270920 550168 270926 550180
rect 319714 550168 319720 550180
rect 270920 550140 319720 550168
rect 270920 550128 270926 550140
rect 319714 550128 319720 550140
rect 319772 550128 319778 550180
rect 59262 550060 59268 550112
rect 59320 550100 59326 550112
rect 98914 550100 98920 550112
rect 59320 550072 98920 550100
rect 59320 550060 59326 550072
rect 98914 550060 98920 550072
rect 98972 550060 98978 550112
rect 106826 550060 106832 550112
rect 106884 550100 106890 550112
rect 124398 550100 124404 550112
rect 106884 550072 124404 550100
rect 106884 550060 106890 550072
rect 124398 550060 124404 550072
rect 124456 550060 124462 550112
rect 136542 550060 136548 550112
rect 136600 550100 136606 550112
rect 164878 550100 164884 550112
rect 136600 550072 164884 550100
rect 136600 550060 136606 550072
rect 164878 550060 164884 550072
rect 164936 550060 164942 550112
rect 170582 550060 170588 550112
rect 170640 550100 170646 550112
rect 200942 550100 200948 550112
rect 170640 550072 200948 550100
rect 170640 550060 170646 550072
rect 200942 550060 200948 550072
rect 201000 550060 201006 550112
rect 212166 550060 212172 550112
rect 212224 550100 212230 550112
rect 236086 550100 236092 550112
rect 212224 550072 236092 550100
rect 212224 550060 212230 550072
rect 236086 550060 236092 550072
rect 236144 550060 236150 550112
rect 252922 550060 252928 550112
rect 252980 550100 252986 550112
rect 319806 550100 319812 550112
rect 252980 550072 319812 550100
rect 252980 550060 252986 550072
rect 319806 550060 319812 550072
rect 319864 550060 319870 550112
rect 56410 549992 56416 550044
rect 56468 550032 56474 550044
rect 73798 550032 73804 550044
rect 56468 550004 73804 550032
rect 56468 549992 56474 550004
rect 73798 549992 73804 550004
rect 73856 549992 73862 550044
rect 78122 549992 78128 550044
rect 78180 550032 78186 550044
rect 121638 550032 121644 550044
rect 78180 550004 121644 550032
rect 78180 549992 78186 550004
rect 121638 549992 121644 550004
rect 121696 549992 121702 550044
rect 136450 549992 136456 550044
rect 136508 550032 136514 550044
rect 171962 550032 171968 550044
rect 136508 550004 171968 550032
rect 136508 549992 136514 550004
rect 171962 549992 171968 550004
rect 172020 549992 172026 550044
rect 176286 549992 176292 550044
rect 176344 550032 176350 550044
rect 213178 550032 213184 550044
rect 176344 550004 213184 550032
rect 176344 549992 176350 550004
rect 213178 549992 213184 550004
rect 213236 549992 213242 550044
rect 217962 549992 217968 550044
rect 218020 550032 218026 550044
rect 230014 550032 230020 550044
rect 218020 550004 230020 550032
rect 218020 549992 218026 550004
rect 230014 549992 230020 550004
rect 230072 549992 230078 550044
rect 231486 549992 231492 550044
rect 231544 550032 231550 550044
rect 238754 550032 238760 550044
rect 231544 550004 238760 550032
rect 231544 549992 231550 550004
rect 238754 549992 238760 550004
rect 238812 549992 238818 550044
rect 239398 549992 239404 550044
rect 239456 550032 239462 550044
rect 284938 550032 284944 550044
rect 239456 550004 284944 550032
rect 239456 549992 239462 550004
rect 284938 549992 284944 550004
rect 284996 549992 285002 550044
rect 54938 549924 54944 549976
rect 54996 549964 55002 549976
rect 99650 549964 99656 549976
rect 54996 549936 99656 549964
rect 54996 549924 55002 549936
rect 99650 549924 99656 549936
rect 99708 549924 99714 549976
rect 103974 549924 103980 549976
rect 104032 549964 104038 549976
rect 124490 549964 124496 549976
rect 104032 549936 124496 549964
rect 104032 549924 104038 549936
rect 124490 549924 124496 549936
rect 124548 549924 124554 549976
rect 146202 549924 146208 549976
rect 146260 549964 146266 549976
rect 201586 549964 201592 549976
rect 146260 549936 201592 549964
rect 146260 549924 146266 549936
rect 201586 549924 201592 549936
rect 201644 549924 201650 549976
rect 220078 549924 220084 549976
rect 220136 549964 220142 549976
rect 233602 549964 233608 549976
rect 220136 549936 233608 549964
rect 220136 549924 220142 549936
rect 233602 549924 233608 549936
rect 233660 549924 233666 549976
rect 237190 549924 237196 549976
rect 237248 549964 237254 549976
rect 284110 549964 284116 549976
rect 237248 549936 284116 549964
rect 237248 549924 237254 549936
rect 284110 549924 284116 549936
rect 284168 549924 284174 549976
rect 299566 549924 299572 549976
rect 299624 549964 299630 549976
rect 319438 549964 319444 549976
rect 299624 549936 319444 549964
rect 299624 549924 299630 549936
rect 319438 549924 319444 549936
rect 319496 549924 319502 549976
rect 61378 549856 61384 549908
rect 61436 549896 61442 549908
rect 116854 549896 116860 549908
rect 61436 549868 116860 549896
rect 61436 549856 61442 549868
rect 116854 549856 116860 549868
rect 116912 549856 116918 549908
rect 139302 549856 139308 549908
rect 139360 549896 139366 549908
rect 175550 549896 175556 549908
rect 139360 549868 175556 549896
rect 139360 549856 139366 549868
rect 175550 549856 175556 549868
rect 175608 549856 175614 549908
rect 182726 549856 182732 549908
rect 182784 549896 182790 549908
rect 242158 549896 242164 549908
rect 182784 549868 242164 549896
rect 182784 549856 182790 549868
rect 242158 549856 242164 549868
rect 242216 549856 242222 549908
rect 245838 549856 245844 549908
rect 245896 549896 245902 549908
rect 281166 549896 281172 549908
rect 245896 549868 281172 549896
rect 245896 549856 245902 549868
rect 281166 549856 281172 549868
rect 281224 549856 281230 549908
rect 281626 549856 281632 549908
rect 281684 549896 281690 549908
rect 303154 549896 303160 549908
rect 281684 549868 303160 549896
rect 281684 549856 281690 549868
rect 303154 549856 303160 549868
rect 303212 549856 303218 549908
rect 278038 549788 278044 549840
rect 278096 549828 278102 549840
rect 300670 549828 300676 549840
rect 278096 549800 300676 549828
rect 278096 549788 278102 549800
rect 300670 549788 300676 549800
rect 300728 549788 300734 549840
rect 277302 549720 277308 549772
rect 277360 549760 277366 549772
rect 300394 549760 300400 549772
rect 277360 549732 300400 549760
rect 277360 549720 277366 549732
rect 300394 549720 300400 549732
rect 300452 549720 300458 549772
rect 276566 549652 276572 549704
rect 276624 549692 276630 549704
rect 301682 549692 301688 549704
rect 276624 549664 301688 549692
rect 276624 549652 276630 549664
rect 301682 549652 301688 549664
rect 301740 549652 301746 549704
rect 273714 549584 273720 549636
rect 273772 549624 273778 549636
rect 301866 549624 301872 549636
rect 273772 549596 301872 549624
rect 273772 549584 273778 549596
rect 301866 549584 301872 549596
rect 301924 549584 301930 549636
rect 296714 549516 296720 549568
rect 296772 549556 296778 549568
rect 315482 549556 315488 549568
rect 296772 549528 315488 549556
rect 296772 549516 296778 549528
rect 315482 549516 315488 549528
rect 315540 549516 315546 549568
rect 240042 549448 240048 549500
rect 240100 549488 240106 549500
rect 266354 549488 266360 549500
rect 240100 549460 266360 549488
rect 240100 549448 240106 549460
rect 266354 549448 266360 549460
rect 266412 549448 266418 549500
rect 275922 549448 275928 549500
rect 275980 549488 275986 549500
rect 316954 549488 316960 549500
rect 275980 549460 316960 549488
rect 275980 549448 275986 549460
rect 316954 549448 316960 549460
rect 317012 549448 317018 549500
rect 280154 549380 280160 549432
rect 280212 549420 280218 549432
rect 280212 549392 282914 549420
rect 280212 549380 280218 549392
rect 61654 549312 61660 549364
rect 61712 549352 61718 549364
rect 64966 549352 64972 549364
rect 61712 549324 64972 549352
rect 61712 549312 61718 549324
rect 64966 549312 64972 549324
rect 65024 549312 65030 549364
rect 102778 549312 102784 549364
rect 102836 549352 102842 549364
rect 106090 549352 106096 549364
rect 102836 549324 106096 549352
rect 102836 549312 102842 549324
rect 106090 549312 106096 549324
rect 106148 549312 106154 549364
rect 108390 549312 108396 549364
rect 108448 549352 108454 549364
rect 114646 549352 114652 549364
rect 108448 549324 114652 549352
rect 108448 549312 108454 549324
rect 114646 549312 114652 549324
rect 114704 549312 114710 549364
rect 118234 549312 118240 549364
rect 118292 549352 118298 549364
rect 124858 549352 124864 549364
rect 118292 549324 124864 549352
rect 118292 549312 118298 549324
rect 124858 549312 124864 549324
rect 124916 549312 124922 549364
rect 131206 549312 131212 549364
rect 131264 549352 131270 549364
rect 134518 549352 134524 549364
rect 131264 549324 134524 549352
rect 131264 549312 131270 549324
rect 134518 549312 134524 549324
rect 134576 549312 134582 549364
rect 203518 549312 203524 549364
rect 203576 549352 203582 549364
rect 211798 549352 211804 549364
rect 203576 549324 211804 549352
rect 203576 549312 203582 549324
rect 211798 549312 211804 549324
rect 211856 549312 211862 549364
rect 243630 549312 243636 549364
rect 243688 549352 243694 549364
rect 273254 549352 273260 549364
rect 243688 549324 273260 549352
rect 243688 549312 243694 549324
rect 273254 549312 273260 549324
rect 273312 549312 273318 549364
rect 282886 549284 282914 549392
rect 298830 549380 298836 549432
rect 298888 549420 298894 549432
rect 319530 549420 319536 549432
rect 298888 549392 319536 549420
rect 298888 549380 298894 549392
rect 319530 549380 319536 549392
rect 319588 549380 319594 549432
rect 284478 549312 284484 549364
rect 284536 549352 284542 549364
rect 300210 549352 300216 549364
rect 284536 549324 300216 549352
rect 284536 549312 284542 549324
rect 300210 549312 300216 549324
rect 300268 549312 300274 549364
rect 302050 549284 302056 549296
rect 282886 549256 302056 549284
rect 302050 549244 302056 549256
rect 302108 549244 302114 549296
rect 295978 548768 295984 548820
rect 296036 548808 296042 548820
rect 315666 548808 315672 548820
rect 296036 548780 315672 548808
rect 296036 548768 296042 548780
rect 315666 548768 315672 548780
rect 315724 548768 315730 548820
rect 268746 548700 268752 548752
rect 268804 548740 268810 548752
rect 300118 548740 300124 548752
rect 268804 548712 300124 548740
rect 268804 548700 268810 548712
rect 300118 548700 300124 548712
rect 300176 548700 300182 548752
rect 265894 548632 265900 548684
rect 265952 548672 265958 548684
rect 301774 548672 301780 548684
rect 265952 548644 301780 548672
rect 265952 548632 265958 548644
rect 301774 548632 301780 548644
rect 301832 548632 301838 548684
rect 273254 548564 273260 548616
rect 273312 548604 273318 548616
rect 318702 548604 318708 548616
rect 273312 548576 318708 548604
rect 273312 548564 273318 548576
rect 318702 548564 318708 548576
rect 318760 548564 318766 548616
rect 266354 548496 266360 548548
rect 266412 548536 266418 548548
rect 318610 548536 318616 548548
rect 266412 548508 318616 548536
rect 266412 548496 266418 548508
rect 318610 548496 318616 548508
rect 318668 548496 318674 548548
rect 265158 548428 265164 548480
rect 265216 548468 265222 548480
rect 305638 548468 305644 548480
rect 265216 548440 305644 548468
rect 265216 548428 265222 548440
rect 305638 548428 305644 548440
rect 305696 548428 305702 548480
rect 260834 548360 260840 548412
rect 260892 548400 260898 548412
rect 304442 548400 304448 548412
rect 260892 548372 304448 548400
rect 260892 548360 260898 548372
rect 304442 548360 304448 548372
rect 304500 548360 304506 548412
rect 254394 548292 254400 548344
rect 254452 548332 254458 548344
rect 302970 548332 302976 548344
rect 254452 548304 302976 548332
rect 254452 548292 254458 548304
rect 302970 548292 302976 548304
rect 303028 548292 303034 548344
rect 236454 548224 236460 548276
rect 236512 548264 236518 548276
rect 301222 548264 301228 548276
rect 236512 548236 301228 548264
rect 236512 548224 236518 548236
rect 301222 548224 301228 548236
rect 301280 548224 301286 548276
rect 249426 548156 249432 548208
rect 249484 548196 249490 548208
rect 319622 548196 319628 548208
rect 249484 548168 319628 548196
rect 249484 548156 249490 548168
rect 319622 548156 319628 548168
rect 319680 548156 319686 548208
rect 235810 548088 235816 548140
rect 235868 548088 235874 548140
rect 247218 548088 247224 548140
rect 247276 548128 247282 548140
rect 319438 548128 319444 548140
rect 247276 548100 319444 548128
rect 247276 548088 247282 548100
rect 319438 548088 319444 548100
rect 319496 548088 319502 548140
rect 235828 548060 235856 548088
rect 319714 548060 319720 548072
rect 235828 548032 319720 548060
rect 319714 548020 319720 548032
rect 319772 548020 319778 548072
rect 301406 547816 301412 547868
rect 301464 547856 301470 547868
rect 317966 547856 317972 547868
rect 301464 547828 317972 547856
rect 301464 547816 301470 547828
rect 317966 547816 317972 547828
rect 318024 547816 318030 547868
rect 301222 542308 301228 542360
rect 301280 542348 301286 542360
rect 317966 542348 317972 542360
rect 301280 542320 317972 542348
rect 301280 542308 301286 542320
rect 317966 542308 317972 542320
rect 318024 542308 318030 542360
rect 302786 539588 302792 539640
rect 302844 539628 302850 539640
rect 311158 539628 311164 539640
rect 302844 539600 311164 539628
rect 302844 539588 302850 539600
rect 311158 539588 311164 539600
rect 311216 539588 311222 539640
rect 312998 528504 313004 528556
rect 313056 528544 313062 528556
rect 495434 528544 495440 528556
rect 313056 528516 495440 528544
rect 313056 528504 313062 528516
rect 495434 528504 495440 528516
rect 495492 528504 495498 528556
rect 313090 528436 313096 528488
rect 313148 528476 313154 528488
rect 476114 528476 476120 528488
rect 313148 528448 476120 528476
rect 313148 528436 313154 528448
rect 476114 528436 476120 528448
rect 476172 528436 476178 528488
rect 315666 528368 315672 528420
rect 315724 528408 315730 528420
rect 457438 528408 457444 528420
rect 315724 528380 457444 528408
rect 315724 528368 315730 528380
rect 457438 528368 457444 528380
rect 457496 528368 457502 528420
rect 300578 528300 300584 528352
rect 300636 528340 300642 528352
rect 430574 528340 430580 528352
rect 300636 528312 430580 528340
rect 300636 528300 300642 528312
rect 430574 528300 430580 528312
rect 430632 528300 430638 528352
rect 300670 528232 300676 528284
rect 300728 528272 300734 528284
rect 431218 528272 431224 528284
rect 300728 528244 431224 528272
rect 300728 528232 300734 528244
rect 431218 528232 431224 528244
rect 431276 528232 431282 528284
rect 301958 528164 301964 528216
rect 302016 528204 302022 528216
rect 431310 528204 431316 528216
rect 302016 528176 431316 528204
rect 302016 528164 302022 528176
rect 431310 528164 431316 528176
rect 431368 528164 431374 528216
rect 302050 528096 302056 528148
rect 302108 528136 302114 528148
rect 431402 528136 431408 528148
rect 302108 528108 431408 528136
rect 302108 528096 302114 528108
rect 431402 528096 431408 528108
rect 431460 528096 431466 528148
rect 318058 528028 318064 528080
rect 318116 528068 318122 528080
rect 430666 528068 430672 528080
rect 318116 528040 430672 528068
rect 318116 528028 318122 528040
rect 430666 528028 430672 528040
rect 430724 528028 430730 528080
rect 319898 527960 319904 528012
rect 319956 528000 319962 528012
rect 431126 528000 431132 528012
rect 319956 527972 431132 528000
rect 319956 527960 319962 527972
rect 431126 527960 431132 527972
rect 431184 527960 431190 528012
rect 319806 527892 319812 527944
rect 319864 527932 319870 527944
rect 430850 527932 430856 527944
rect 319864 527904 430856 527932
rect 319864 527892 319870 527904
rect 430850 527892 430856 527904
rect 430908 527892 430914 527944
rect 318518 527824 318524 527876
rect 318576 527864 318582 527876
rect 429562 527864 429568 527876
rect 318576 527836 429568 527864
rect 318576 527824 318582 527836
rect 429562 527824 429568 527836
rect 429620 527824 429626 527876
rect 318426 527756 318432 527808
rect 318484 527796 318490 527808
rect 428366 527796 428372 527808
rect 318484 527768 428372 527796
rect 318484 527756 318490 527768
rect 428366 527756 428372 527768
rect 428424 527756 428430 527808
rect 304258 527212 304264 527264
rect 304316 527252 304322 527264
rect 369302 527252 369308 527264
rect 304316 527224 369308 527252
rect 304316 527212 304322 527224
rect 369302 527212 369308 527224
rect 369360 527212 369366 527264
rect 301866 527144 301872 527196
rect 301924 527184 301930 527196
rect 396902 527184 396908 527196
rect 301924 527156 396908 527184
rect 301924 527144 301930 527156
rect 396902 527144 396908 527156
rect 396960 527144 396966 527196
rect 312906 527076 312912 527128
rect 312964 527116 312970 527128
rect 512270 527116 512276 527128
rect 312964 527088 512276 527116
rect 312964 527076 312970 527088
rect 512270 527076 512276 527088
rect 512328 527076 512334 527128
rect 315574 527008 315580 527060
rect 315632 527048 315638 527060
rect 500954 527048 500960 527060
rect 315632 527020 500960 527048
rect 315632 527008 315638 527020
rect 500954 527008 500960 527020
rect 501012 527008 501018 527060
rect 309778 526940 309784 526992
rect 309836 526980 309842 526992
rect 457806 526980 457812 526992
rect 309836 526952 457812 526980
rect 309836 526940 309842 526952
rect 457806 526940 457812 526952
rect 457864 526940 457870 526992
rect 315482 526872 315488 526924
rect 315540 526912 315546 526924
rect 459554 526912 459560 526924
rect 315540 526884 459560 526912
rect 315540 526872 315546 526884
rect 459554 526872 459560 526884
rect 459612 526872 459618 526924
rect 319530 526804 319536 526856
rect 319588 526844 319594 526856
rect 457622 526844 457628 526856
rect 319588 526816 457628 526844
rect 319588 526804 319594 526816
rect 457622 526804 457628 526816
rect 457680 526804 457686 526856
rect 300394 526736 300400 526788
rect 300452 526776 300458 526788
rect 430942 526776 430948 526788
rect 300452 526748 430948 526776
rect 300452 526736 300458 526748
rect 430942 526736 430948 526748
rect 431000 526736 431006 526788
rect 300210 526668 300216 526720
rect 300268 526708 300274 526720
rect 430758 526708 430764 526720
rect 300268 526680 430764 526708
rect 300268 526668 300274 526680
rect 430758 526668 430764 526680
rect 430816 526668 430822 526720
rect 303154 526600 303160 526652
rect 303212 526640 303218 526652
rect 431034 526640 431040 526652
rect 303212 526612 431040 526640
rect 303212 526600 303218 526612
rect 431034 526600 431040 526612
rect 431092 526600 431098 526652
rect 315390 526532 315396 526584
rect 315448 526572 315454 526584
rect 429470 526572 429476 526584
rect 315448 526544 429476 526572
rect 315448 526532 315454 526544
rect 429470 526532 429476 526544
rect 429528 526532 429534 526584
rect 301682 526464 301688 526516
rect 301740 526504 301746 526516
rect 414934 526504 414940 526516
rect 301740 526476 414940 526504
rect 301740 526464 301746 526476
rect 414934 526464 414940 526476
rect 414992 526464 414998 526516
rect 324866 526396 324872 526448
rect 324924 526436 324930 526448
rect 429194 526436 429200 526448
rect 324924 526408 429200 526436
rect 324924 526396 324930 526408
rect 429194 526396 429200 526408
rect 429252 526396 429258 526448
rect 316954 526328 316960 526380
rect 317012 526368 317018 526380
rect 351270 526368 351276 526380
rect 317012 526340 351276 526368
rect 317012 526328 317018 526340
rect 351270 526328 351276 526340
rect 351328 526328 351334 526380
rect 313918 526260 313924 526312
rect 313976 526300 313982 526312
rect 337654 526300 337660 526312
rect 313976 526272 337660 526300
rect 313976 526260 313982 526272
rect 337654 526260 337660 526272
rect 337712 526260 337718 526312
rect 300486 526192 300492 526244
rect 300544 526232 300550 526244
rect 328638 526232 328644 526244
rect 300544 526204 328644 526232
rect 300544 526192 300550 526204
rect 328638 526192 328644 526204
rect 328696 526192 328702 526244
rect 319622 525716 319628 525768
rect 319680 525756 319686 525768
rect 423950 525756 423956 525768
rect 319680 525728 423956 525756
rect 319680 525716 319686 525728
rect 423950 525716 423956 525728
rect 424008 525716 424014 525768
rect 319714 525648 319720 525700
rect 319772 525688 319778 525700
rect 319772 525660 320220 525688
rect 319772 525648 319778 525660
rect 305638 525580 305644 525632
rect 305696 525620 305702 525632
rect 320082 525620 320088 525632
rect 305696 525592 320088 525620
rect 305696 525580 305702 525592
rect 320082 525580 320088 525592
rect 320140 525580 320146 525632
rect 320192 525620 320220 525660
rect 320450 525648 320456 525700
rect 320508 525688 320514 525700
rect 419534 525688 419540 525700
rect 320508 525660 419540 525688
rect 320508 525648 320514 525660
rect 419534 525648 419540 525660
rect 419592 525648 419598 525700
rect 333238 525620 333244 525632
rect 320192 525592 333244 525620
rect 333238 525580 333244 525592
rect 333296 525580 333302 525632
rect 318242 525512 318248 525564
rect 318300 525552 318306 525564
rect 320266 525552 320272 525564
rect 318300 525524 320272 525552
rect 318300 525512 318306 525524
rect 320266 525512 320272 525524
rect 320324 525512 320330 525564
rect 320542 525512 320548 525564
rect 320600 525552 320606 525564
rect 405918 525552 405924 525564
rect 320600 525524 405924 525552
rect 320600 525512 320606 525524
rect 405918 525512 405924 525524
rect 405976 525512 405982 525564
rect 300118 525444 300124 525496
rect 300176 525484 300182 525496
rect 387886 525484 387892 525496
rect 300176 525456 387892 525484
rect 300176 525444 300182 525456
rect 387886 525444 387892 525456
rect 387944 525444 387950 525496
rect 316678 525376 316684 525428
rect 316736 525416 316742 525428
rect 320358 525416 320364 525428
rect 316736 525388 320364 525416
rect 316736 525376 316742 525388
rect 320358 525376 320364 525388
rect 320416 525376 320422 525428
rect 320634 525376 320640 525428
rect 320692 525416 320698 525428
rect 401594 525416 401600 525428
rect 320692 525388 401600 525416
rect 320692 525376 320698 525388
rect 401594 525376 401600 525388
rect 401652 525376 401658 525428
rect 301774 525308 301780 525360
rect 301832 525348 301838 525360
rect 383654 525348 383660 525360
rect 301832 525320 383660 525348
rect 301832 525308 301838 525320
rect 383654 525308 383660 525320
rect 383712 525308 383718 525360
rect 302878 525240 302884 525292
rect 302936 525280 302942 525292
rect 364702 525280 364708 525292
rect 302936 525252 364708 525280
rect 302936 525240 302942 525252
rect 364702 525240 364708 525252
rect 364760 525240 364766 525292
rect 318150 525172 318156 525224
rect 318208 525212 318214 525224
rect 374454 525212 374460 525224
rect 318208 525184 374460 525212
rect 318208 525172 318214 525184
rect 374454 525172 374460 525184
rect 374512 525172 374518 525224
rect 301590 525104 301596 525156
rect 301648 525144 301654 525156
rect 356238 525144 356244 525156
rect 301648 525116 356244 525144
rect 301648 525104 301654 525116
rect 356238 525104 356244 525116
rect 356296 525104 356302 525156
rect 319438 525036 319444 525088
rect 319496 525076 319502 525088
rect 360286 525076 360292 525088
rect 319496 525048 360292 525076
rect 319496 525036 319502 525048
rect 360286 525036 360292 525048
rect 360344 525036 360350 525088
rect 302970 524968 302976 525020
rect 303028 525008 303034 525020
rect 346670 525008 346676 525020
rect 303028 524980 346676 525008
rect 303028 524968 303034 524980
rect 346670 524968 346676 524980
rect 346728 524968 346734 525020
rect 304442 524900 304448 524952
rect 304500 524940 304506 524952
rect 342254 524940 342260 524952
rect 304500 524912 342260 524940
rect 304500 524900 304506 524912
rect 342254 524900 342260 524912
rect 342312 524900 342318 524952
rect 318334 524832 318340 524884
rect 318392 524872 318398 524884
rect 410518 524872 410524 524884
rect 318392 524844 410524 524872
rect 318392 524832 318398 524844
rect 410518 524832 410524 524844
rect 410576 524832 410582 524884
rect 314010 524764 314016 524816
rect 314068 524804 314074 524816
rect 320634 524804 320640 524816
rect 314068 524776 320640 524804
rect 314068 524764 314074 524776
rect 320634 524764 320640 524776
rect 320692 524764 320698 524816
rect 304350 524356 304356 524408
rect 304408 524396 304414 524408
rect 512178 524396 512184 524408
rect 304408 524368 512184 524396
rect 304408 524356 304414 524368
rect 512178 524356 512184 524368
rect 512236 524356 512242 524408
rect 301498 524288 301504 524340
rect 301556 524328 301562 524340
rect 488534 524328 488540 524340
rect 301556 524300 488540 524328
rect 301556 524288 301562 524300
rect 488534 524288 488540 524300
rect 488592 524288 488598 524340
rect 312814 524220 312820 524272
rect 312872 524260 312878 524272
rect 470594 524260 470600 524272
rect 312872 524232 470600 524260
rect 312872 524220 312878 524232
rect 470594 524220 470600 524232
rect 470652 524220 470658 524272
rect 302326 523676 302332 523728
rect 302384 523716 302390 523728
rect 578878 523716 578884 523728
rect 302384 523688 578884 523716
rect 302384 523676 302390 523688
rect 578878 523676 578884 523688
rect 578936 523676 578942 523728
rect 312630 522928 312636 522980
rect 312688 522968 312694 522980
rect 465074 522968 465080 522980
rect 312688 522940 465080 522968
rect 312688 522928 312694 522940
rect 465074 522928 465080 522940
rect 465132 522928 465138 522980
rect 312722 522860 312728 522912
rect 312780 522900 312786 522912
rect 457714 522900 457720 522912
rect 312780 522872 457720 522900
rect 312780 522860 312786 522872
rect 457714 522860 457720 522872
rect 457772 522860 457778 522912
rect 315298 522792 315304 522844
rect 315356 522832 315362 522844
rect 429654 522832 429660 522844
rect 315356 522804 429660 522832
rect 315356 522792 315362 522804
rect 429654 522792 429660 522804
rect 429712 522792 429718 522844
rect 316862 522724 316868 522776
rect 316920 522764 316926 522776
rect 427814 522764 427820 522776
rect 316920 522736 427820 522764
rect 316920 522724 316926 522736
rect 427814 522724 427820 522736
rect 427872 522724 427878 522776
rect 44082 518168 44088 518220
rect 44140 518208 44146 518220
rect 57882 518208 57888 518220
rect 44140 518180 57888 518208
rect 44140 518168 44146 518180
rect 57882 518168 57888 518180
rect 57940 518168 57946 518220
rect 311158 515380 311164 515432
rect 311216 515420 311222 515432
rect 580258 515420 580264 515432
rect 311216 515392 580264 515420
rect 311216 515380 311222 515392
rect 580258 515380 580264 515392
rect 580316 515380 580322 515432
rect 560938 511912 560944 511964
rect 560996 511952 561002 511964
rect 580166 511952 580172 511964
rect 560996 511924 580172 511952
rect 560996 511912 561002 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 302234 495456 302240 495508
rect 302292 495496 302298 495508
rect 520918 495496 520924 495508
rect 302292 495468 520924 495496
rect 302292 495456 302298 495468
rect 520918 495456 520924 495468
rect 520976 495456 520982 495508
rect 201510 487772 201516 487824
rect 201568 487812 201574 487824
rect 201770 487812 201776 487824
rect 201568 487784 201776 487812
rect 201568 487772 201574 487784
rect 201770 487772 201776 487784
rect 201828 487772 201834 487824
rect 274650 487772 274656 487824
rect 274708 487812 274714 487824
rect 274818 487812 274824 487824
rect 274708 487784 274824 487812
rect 274708 487772 274714 487784
rect 274818 487772 274824 487784
rect 274876 487772 274882 487824
rect 128354 487024 128360 487076
rect 128412 487064 128418 487076
rect 128630 487064 128636 487076
rect 128412 487036 128636 487064
rect 128412 487024 128418 487036
rect 128630 487024 128636 487036
rect 128688 487024 128694 487076
rect 178034 487024 178040 487076
rect 178092 487064 178098 487076
rect 178310 487064 178316 487076
rect 178092 487036 178316 487064
rect 178092 487024 178098 487036
rect 178310 487024 178316 487036
rect 178368 487024 178374 487076
rect 248506 487024 248512 487076
rect 248564 487064 248570 487076
rect 248782 487064 248788 487076
rect 248564 487036 248788 487064
rect 248564 487024 248570 487036
rect 248782 487024 248788 487036
rect 248840 487024 248846 487076
rect 140866 486480 140872 486532
rect 140924 486520 140930 486532
rect 199010 486520 199016 486532
rect 140924 486492 199016 486520
rect 140924 486480 140930 486492
rect 199010 486480 199016 486492
rect 199068 486480 199074 486532
rect 14458 486412 14464 486464
rect 14516 486452 14522 486464
rect 378134 486452 378140 486464
rect 14516 486424 378140 486452
rect 14516 486412 14522 486424
rect 378134 486412 378140 486424
rect 378192 486412 378198 486464
rect 53742 485732 53748 485784
rect 53800 485772 53806 485784
rect 74258 485772 74264 485784
rect 53800 485744 74264 485772
rect 53800 485732 53806 485744
rect 74258 485732 74264 485744
rect 74316 485732 74322 485784
rect 74350 485732 74356 485784
rect 74408 485772 74414 485784
rect 102870 485772 102876 485784
rect 74408 485744 102876 485772
rect 74408 485732 74414 485744
rect 102870 485732 102876 485744
rect 102928 485732 102934 485784
rect 152182 485732 152188 485784
rect 152240 485772 152246 485784
rect 209774 485772 209780 485784
rect 152240 485744 209780 485772
rect 152240 485732 152246 485744
rect 209774 485732 209780 485744
rect 209832 485732 209838 485784
rect 209866 485732 209872 485784
rect 209924 485772 209930 485784
rect 219894 485772 219900 485784
rect 209924 485744 219900 485772
rect 209924 485732 209930 485744
rect 219894 485732 219900 485744
rect 219952 485732 219958 485784
rect 56502 485664 56508 485716
rect 56560 485704 56566 485716
rect 89162 485704 89168 485716
rect 56560 485676 89168 485704
rect 56560 485664 56566 485676
rect 89162 485664 89168 485676
rect 89220 485664 89226 485716
rect 150434 485664 150440 485716
rect 150492 485704 150498 485716
rect 150492 485676 205772 485704
rect 150492 485664 150498 485676
rect 59998 485596 60004 485648
rect 60056 485636 60062 485648
rect 91830 485636 91836 485648
rect 60056 485608 91836 485636
rect 60056 485596 60062 485608
rect 91830 485596 91836 485608
rect 91888 485596 91894 485648
rect 149514 485596 149520 485648
rect 149572 485636 149578 485648
rect 205634 485636 205640 485648
rect 149572 485608 205640 485636
rect 149572 485596 149578 485608
rect 205634 485596 205640 485608
rect 205692 485596 205698 485648
rect 205744 485636 205772 485676
rect 208210 485664 208216 485716
rect 208268 485704 208274 485716
rect 217778 485704 217784 485716
rect 208268 485676 217784 485704
rect 208268 485664 208274 485676
rect 217778 485664 217784 485676
rect 217836 485664 217842 485716
rect 208394 485636 208400 485648
rect 205744 485608 208400 485636
rect 208394 485596 208400 485608
rect 208452 485596 208458 485648
rect 209774 485596 209780 485648
rect 209832 485636 209838 485648
rect 211246 485636 211252 485648
rect 209832 485608 211252 485636
rect 209832 485596 209838 485608
rect 211246 485596 211252 485608
rect 211304 485596 211310 485648
rect 56318 485528 56324 485580
rect 56376 485568 56382 485580
rect 88334 485568 88340 485580
rect 56376 485540 88340 485568
rect 56376 485528 56382 485540
rect 88334 485528 88340 485540
rect 88392 485528 88398 485580
rect 151262 485528 151268 485580
rect 151320 485568 151326 485580
rect 205726 485568 205732 485580
rect 151320 485540 205732 485568
rect 151320 485528 151326 485540
rect 205726 485528 205732 485540
rect 205784 485528 205790 485580
rect 211154 485568 211160 485580
rect 209746 485540 211160 485568
rect 50890 485460 50896 485512
rect 50948 485500 50954 485512
rect 79318 485500 79324 485512
rect 50948 485472 79324 485500
rect 50948 485460 50954 485472
rect 79318 485460 79324 485472
rect 79376 485460 79382 485512
rect 157702 485460 157708 485512
rect 157760 485500 157766 485512
rect 209746 485500 209774 485540
rect 211154 485528 211160 485540
rect 211212 485528 211218 485580
rect 244550 485528 244556 485580
rect 244608 485568 244614 485580
rect 356790 485568 356796 485580
rect 244608 485540 356796 485568
rect 244608 485528 244614 485540
rect 356790 485528 356796 485540
rect 356848 485528 356854 485580
rect 157760 485472 209774 485500
rect 157760 485460 157766 485472
rect 239674 485460 239680 485512
rect 239732 485500 239738 485512
rect 358262 485500 358268 485512
rect 239732 485472 358268 485500
rect 239732 485460 239738 485472
rect 358262 485460 358268 485472
rect 358320 485460 358326 485512
rect 56226 485392 56232 485444
rect 56284 485432 56290 485444
rect 90542 485432 90548 485444
rect 56284 485404 90548 485432
rect 56284 485392 56290 485404
rect 90542 485392 90548 485404
rect 90600 485392 90606 485444
rect 149422 485392 149428 485444
rect 149480 485432 149486 485444
rect 149480 485404 191144 485432
rect 149480 485392 149486 485404
rect 79226 485324 79232 485376
rect 79284 485364 79290 485376
rect 104158 485364 104164 485376
rect 79284 485336 104164 485364
rect 79284 485324 79290 485336
rect 104158 485324 104164 485336
rect 104216 485324 104222 485376
rect 157426 485324 157432 485376
rect 157484 485364 157490 485376
rect 188338 485364 188344 485376
rect 157484 485336 188344 485364
rect 157484 485324 157490 485336
rect 188338 485324 188344 485336
rect 188396 485324 188402 485376
rect 191116 485364 191144 485404
rect 191190 485392 191196 485444
rect 191248 485432 191254 485444
rect 205634 485432 205640 485444
rect 191248 485404 205640 485432
rect 191248 485392 191254 485404
rect 205634 485392 205640 485404
rect 205692 485392 205698 485444
rect 209314 485392 209320 485444
rect 209372 485432 209378 485444
rect 219066 485432 219072 485444
rect 209372 485404 219072 485432
rect 209372 485392 209378 485404
rect 219066 485392 219072 485404
rect 219124 485392 219130 485444
rect 240042 485392 240048 485444
rect 240100 485432 240106 485444
rect 358354 485432 358360 485444
rect 240100 485404 358360 485432
rect 240100 485392 240106 485404
rect 358354 485392 358360 485404
rect 358412 485392 358418 485444
rect 191116 485336 193214 485364
rect 68278 485256 68284 485308
rect 68336 485296 68342 485308
rect 105538 485296 105544 485308
rect 68336 485268 105544 485296
rect 68336 485256 68342 485268
rect 105538 485256 105544 485268
rect 105596 485256 105602 485308
rect 156690 485256 156696 485308
rect 156748 485296 156754 485308
rect 157702 485296 157708 485308
rect 156748 485268 157708 485296
rect 156748 485256 156754 485268
rect 157702 485256 157708 485268
rect 157760 485256 157766 485308
rect 157794 485256 157800 485308
rect 157852 485296 157858 485308
rect 189258 485296 189264 485308
rect 157852 485268 189264 485296
rect 157852 485256 157858 485268
rect 189258 485256 189264 485268
rect 189316 485256 189322 485308
rect 193186 485296 193214 485336
rect 206922 485324 206928 485376
rect 206980 485364 206986 485376
rect 219158 485364 219164 485376
rect 206980 485336 219164 485364
rect 206980 485324 206986 485336
rect 219158 485324 219164 485336
rect 219216 485324 219222 485376
rect 234522 485324 234528 485376
rect 234580 485364 234586 485376
rect 364978 485364 364984 485376
rect 234580 485336 364984 485364
rect 234580 485324 234586 485336
rect 364978 485324 364984 485336
rect 365036 485324 365042 485376
rect 200298 485296 200304 485308
rect 193186 485268 200304 485296
rect 200298 485256 200304 485268
rect 200356 485256 200362 485308
rect 200390 485256 200396 485308
rect 200448 485296 200454 485308
rect 200448 485268 208992 485296
rect 200448 485256 200454 485268
rect 55950 485188 55956 485240
rect 56008 485228 56014 485240
rect 103330 485228 103336 485240
rect 56008 485200 103336 485228
rect 56008 485188 56014 485200
rect 103330 485188 103336 485200
rect 103388 485188 103394 485240
rect 154298 485188 154304 485240
rect 154356 485228 154362 485240
rect 200482 485228 200488 485240
rect 154356 485200 200488 485228
rect 154356 485188 154362 485200
rect 200482 485188 200488 485200
rect 200540 485188 200546 485240
rect 208964 485228 208992 485268
rect 209498 485256 209504 485308
rect 209556 485296 209562 485308
rect 221734 485296 221740 485308
rect 209556 485268 221740 485296
rect 209556 485256 209562 485268
rect 221734 485256 221740 485268
rect 221792 485256 221798 485308
rect 226058 485256 226064 485308
rect 226116 485296 226122 485308
rect 356698 485296 356704 485308
rect 226116 485268 356704 485296
rect 226116 485256 226122 485268
rect 356698 485256 356704 485268
rect 356756 485256 356762 485308
rect 217502 485228 217508 485240
rect 208964 485200 217508 485228
rect 217502 485188 217508 485200
rect 217560 485188 217566 485240
rect 224218 485188 224224 485240
rect 224276 485228 224282 485240
rect 358170 485228 358176 485240
rect 224276 485200 358176 485228
rect 224276 485188 224282 485200
rect 358170 485188 358176 485200
rect 358228 485188 358234 485240
rect 61010 485120 61016 485172
rect 61068 485160 61074 485172
rect 116578 485160 116584 485172
rect 61068 485132 116584 485160
rect 61068 485120 61074 485132
rect 116578 485120 116584 485132
rect 116636 485120 116642 485172
rect 139210 485120 139216 485172
rect 139268 485160 139274 485172
rect 139268 485132 186314 485160
rect 139268 485120 139274 485132
rect 51626 485052 51632 485104
rect 51684 485092 51690 485104
rect 100662 485092 100668 485104
rect 51684 485064 100668 485092
rect 51684 485052 51690 485064
rect 100662 485052 100668 485064
rect 100720 485052 100726 485104
rect 110322 485052 110328 485104
rect 110380 485092 110386 485104
rect 180058 485092 180064 485104
rect 110380 485064 180064 485092
rect 110380 485052 110386 485064
rect 180058 485052 180064 485064
rect 180116 485052 180122 485104
rect 186286 485092 186314 485132
rect 188338 485120 188344 485172
rect 188396 485160 188402 485172
rect 191190 485160 191196 485172
rect 188396 485132 191196 485160
rect 188396 485120 188402 485132
rect 191190 485120 191196 485132
rect 191248 485120 191254 485172
rect 212350 485160 212356 485172
rect 197740 485132 212356 485160
rect 193858 485092 193864 485104
rect 186286 485064 193864 485092
rect 193858 485052 193864 485064
rect 193916 485052 193922 485104
rect 195330 485052 195336 485104
rect 195388 485092 195394 485104
rect 197740 485092 197768 485132
rect 212350 485120 212356 485132
rect 212408 485120 212414 485172
rect 230658 485120 230664 485172
rect 230716 485160 230722 485172
rect 366358 485160 366364 485172
rect 230716 485132 366364 485160
rect 230716 485120 230722 485132
rect 366358 485120 366364 485132
rect 366416 485120 366422 485172
rect 195388 485064 197768 485092
rect 195388 485052 195394 485064
rect 199930 485052 199936 485104
rect 199988 485092 199994 485104
rect 217410 485092 217416 485104
rect 199988 485064 217416 485092
rect 199988 485052 199994 485064
rect 217410 485052 217416 485064
rect 217468 485052 217474 485104
rect 225598 485052 225604 485104
rect 225656 485092 225662 485104
rect 362218 485092 362224 485104
rect 225656 485064 362224 485092
rect 225656 485052 225662 485064
rect 362218 485052 362224 485064
rect 362276 485052 362282 485104
rect 56410 484984 56416 485036
rect 56468 485024 56474 485036
rect 56468 484996 78168 485024
rect 56468 484984 56474 484996
rect 64138 484916 64144 484968
rect 64196 484956 64202 484968
rect 72418 484956 72424 484968
rect 64196 484928 72424 484956
rect 64196 484916 64202 484928
rect 72418 484916 72424 484928
rect 72476 484916 72482 484968
rect 73798 484916 73804 484968
rect 73856 484956 73862 484968
rect 78030 484956 78036 484968
rect 73856 484928 78036 484956
rect 73856 484916 73862 484928
rect 78030 484916 78036 484928
rect 78088 484916 78094 484968
rect 58526 484848 58532 484900
rect 58584 484888 58590 484900
rect 78140 484888 78168 484996
rect 79318 484984 79324 485036
rect 79376 485024 79382 485036
rect 84378 485024 84384 485036
rect 79376 484996 84384 485024
rect 79376 484984 79382 484996
rect 84378 484984 84384 484996
rect 84436 484984 84442 485036
rect 139394 484984 139400 485036
rect 139452 485024 139458 485036
rect 185578 485024 185584 485036
rect 139452 484996 185584 485024
rect 139452 484984 139458 484996
rect 185578 484984 185584 484996
rect 185636 484984 185642 485036
rect 189258 484984 189264 485036
rect 189316 485024 189322 485036
rect 201494 485024 201500 485036
rect 189316 484996 201500 485024
rect 189316 484984 189322 484996
rect 201494 484984 201500 484996
rect 201552 484984 201558 485036
rect 78214 484916 78220 484968
rect 78272 484956 78278 484968
rect 100202 484956 100208 484968
rect 78272 484928 100208 484956
rect 78272 484916 78278 484928
rect 100202 484916 100208 484928
rect 100260 484916 100266 484968
rect 158622 484916 158628 484968
rect 158680 484956 158686 484968
rect 197446 484956 197452 484968
rect 158680 484928 197452 484956
rect 158680 484916 158686 484928
rect 197446 484916 197452 484928
rect 197504 484916 197510 484968
rect 81710 484888 81716 484900
rect 58584 484860 64874 484888
rect 78140 484860 81716 484888
rect 58584 484848 58590 484860
rect 64846 484820 64874 484860
rect 81710 484848 81716 484860
rect 81768 484848 81774 484900
rect 204898 484888 204904 484900
rect 171106 484860 204904 484888
rect 81250 484820 81256 484832
rect 64846 484792 81256 484820
rect 81250 484780 81256 484792
rect 81308 484780 81314 484832
rect 155310 484780 155316 484832
rect 155368 484820 155374 484832
rect 157794 484820 157800 484832
rect 155368 484792 157800 484820
rect 155368 484780 155374 484792
rect 157794 484780 157800 484792
rect 157852 484780 157858 484832
rect 68370 484712 68376 484764
rect 68428 484752 68434 484764
rect 79226 484752 79232 484764
rect 68428 484724 79232 484752
rect 68428 484712 68434 484724
rect 79226 484712 79232 484724
rect 79284 484712 79290 484764
rect 166074 484712 166080 484764
rect 166132 484752 166138 484764
rect 171106 484752 171134 484860
rect 204898 484848 204904 484860
rect 204956 484848 204962 484900
rect 166132 484724 171134 484752
rect 166132 484712 166138 484724
rect 291028 484452 292160 484480
rect 50982 484372 50988 484424
rect 51040 484412 51046 484424
rect 68462 484412 68468 484424
rect 51040 484384 68468 484412
rect 51040 484372 51046 484384
rect 68462 484372 68468 484384
rect 68520 484372 68526 484424
rect 195146 484372 195152 484424
rect 195204 484412 195210 484424
rect 197078 484412 197084 484424
rect 195204 484384 197084 484412
rect 195204 484372 195210 484384
rect 197078 484372 197084 484384
rect 197136 484372 197142 484424
rect 205910 484372 205916 484424
rect 205968 484412 205974 484424
rect 207658 484412 207664 484424
rect 205968 484384 207664 484412
rect 205968 484372 205974 484384
rect 207658 484372 207664 484384
rect 207716 484372 207722 484424
rect 211706 484372 211712 484424
rect 211764 484412 211770 484424
rect 212810 484412 212816 484424
rect 211764 484384 212816 484412
rect 211764 484372 211770 484384
rect 212810 484372 212816 484384
rect 212868 484372 212874 484424
rect 213362 484372 213368 484424
rect 213420 484412 213426 484424
rect 215018 484412 215024 484424
rect 213420 484384 215024 484412
rect 213420 484372 213426 484384
rect 215018 484372 215024 484384
rect 215076 484372 215082 484424
rect 217042 484372 217048 484424
rect 217100 484412 217106 484424
rect 218146 484412 218152 484424
rect 217100 484384 218152 484412
rect 217100 484372 217106 484384
rect 218146 484372 218152 484384
rect 218204 484372 218210 484424
rect 220170 484372 220176 484424
rect 220228 484412 220234 484424
rect 222654 484412 222660 484424
rect 220228 484384 222660 484412
rect 220228 484372 220234 484384
rect 222654 484372 222660 484384
rect 222712 484372 222718 484424
rect 285490 484304 285496 484356
rect 285548 484344 285554 484356
rect 291028 484344 291056 484452
rect 285548 484316 291056 484344
rect 291120 484384 292068 484412
rect 285548 484304 285554 484316
rect 285858 484236 285864 484288
rect 285916 484276 285922 484288
rect 286134 484276 286140 484288
rect 285916 484248 286140 484276
rect 285916 484236 285922 484248
rect 286134 484236 286140 484248
rect 286192 484236 286198 484288
rect 289722 484236 289728 484288
rect 289780 484276 289786 484288
rect 291120 484276 291148 484384
rect 289780 484248 291148 484276
rect 289780 484236 289786 484248
rect 291194 484236 291200 484288
rect 291252 484276 291258 484288
rect 291930 484276 291936 484288
rect 291252 484248 291936 484276
rect 291252 484236 291258 484248
rect 291930 484236 291936 484248
rect 291988 484236 291994 484288
rect 292040 484276 292068 484384
rect 292132 484344 292160 484452
rect 358078 484344 358084 484356
rect 292132 484316 358084 484344
rect 358078 484304 358084 484316
rect 358136 484304 358142 484356
rect 371142 484276 371148 484288
rect 292040 484248 371148 484276
rect 371142 484236 371148 484248
rect 371200 484236 371206 484288
rect 62114 484168 62120 484220
rect 62172 484208 62178 484220
rect 62942 484208 62948 484220
rect 62172 484180 62948 484208
rect 62172 484168 62178 484180
rect 62942 484168 62948 484180
rect 63000 484168 63006 484220
rect 78674 484168 78680 484220
rect 78732 484208 78738 484220
rect 79686 484208 79692 484220
rect 78732 484180 79692 484208
rect 78732 484168 78738 484180
rect 79686 484168 79692 484180
rect 79744 484168 79750 484220
rect 92566 484168 92572 484220
rect 92624 484208 92630 484220
rect 93302 484208 93308 484220
rect 92624 484180 93308 484208
rect 92624 484168 92630 484180
rect 93302 484168 93308 484180
rect 93360 484168 93366 484220
rect 140774 484168 140780 484220
rect 140832 484208 140838 484220
rect 141694 484208 141700 484220
rect 140832 484180 141700 484208
rect 140832 484168 140838 484180
rect 141694 484168 141700 484180
rect 141752 484168 141758 484220
rect 142246 484168 142252 484220
rect 142304 484208 142310 484220
rect 142982 484208 142988 484220
rect 142304 484180 142988 484208
rect 142304 484168 142310 484180
rect 142982 484168 142988 484180
rect 143040 484168 143046 484220
rect 207106 484168 207112 484220
rect 207164 484208 207170 484220
rect 207750 484208 207756 484220
rect 207164 484180 207756 484208
rect 207164 484168 207170 484180
rect 207750 484168 207756 484180
rect 207808 484168 207814 484220
rect 280062 484168 280068 484220
rect 280120 484208 280126 484220
rect 366910 484208 366916 484220
rect 280120 484180 366916 484208
rect 280120 484168 280126 484180
rect 366910 484168 366916 484180
rect 366968 484168 366974 484220
rect 62206 484100 62212 484152
rect 62264 484140 62270 484152
rect 62390 484140 62396 484152
rect 62264 484112 62396 484140
rect 62264 484100 62270 484112
rect 62390 484100 62396 484112
rect 62448 484100 62454 484152
rect 67726 484100 67732 484152
rect 67784 484140 67790 484152
rect 68186 484140 68192 484152
rect 67784 484112 68192 484140
rect 67784 484100 67790 484112
rect 68186 484100 68192 484112
rect 68244 484100 68250 484152
rect 69014 484100 69020 484152
rect 69072 484140 69078 484152
rect 69566 484140 69572 484152
rect 69072 484112 69572 484140
rect 69072 484100 69078 484112
rect 69566 484100 69572 484112
rect 69624 484100 69630 484152
rect 70394 484100 70400 484152
rect 70452 484140 70458 484152
rect 70854 484140 70860 484152
rect 70452 484112 70860 484140
rect 70452 484100 70458 484112
rect 70854 484100 70860 484112
rect 70912 484100 70918 484152
rect 71866 484100 71872 484152
rect 71924 484140 71930 484152
rect 72602 484140 72608 484152
rect 71924 484112 72608 484140
rect 71924 484100 71930 484112
rect 72602 484100 72608 484112
rect 72660 484100 72666 484152
rect 74534 484100 74540 484152
rect 74592 484140 74598 484152
rect 74718 484140 74724 484152
rect 74592 484112 74724 484140
rect 74592 484100 74598 484112
rect 74718 484100 74724 484112
rect 74776 484100 74782 484152
rect 75914 484100 75920 484152
rect 75972 484140 75978 484152
rect 76558 484140 76564 484152
rect 75972 484112 76564 484140
rect 75972 484100 75978 484112
rect 76558 484100 76564 484112
rect 76616 484100 76622 484152
rect 78766 484100 78772 484152
rect 78824 484140 78830 484152
rect 78950 484140 78956 484152
rect 78824 484112 78956 484140
rect 78824 484100 78830 484112
rect 78950 484100 78956 484112
rect 79008 484100 79014 484152
rect 92474 484100 92480 484152
rect 92532 484140 92538 484152
rect 92934 484140 92940 484152
rect 92532 484112 92940 484140
rect 92532 484100 92538 484112
rect 92934 484100 92940 484112
rect 92992 484100 92998 484152
rect 93854 484100 93860 484152
rect 93912 484140 93918 484152
rect 94590 484140 94596 484152
rect 93912 484112 94596 484140
rect 93912 484100 93918 484112
rect 94590 484100 94596 484112
rect 94648 484100 94654 484152
rect 100754 484100 100760 484152
rect 100812 484140 100818 484152
rect 101582 484140 101588 484152
rect 100812 484112 101588 484140
rect 100812 484100 100818 484112
rect 101582 484100 101588 484112
rect 101640 484100 101646 484152
rect 106274 484100 106280 484152
rect 106332 484140 106338 484152
rect 106918 484140 106924 484152
rect 106332 484112 106924 484140
rect 106332 484100 106338 484112
rect 106918 484100 106924 484112
rect 106976 484100 106982 484152
rect 107654 484100 107660 484152
rect 107712 484140 107718 484152
rect 108206 484140 108212 484152
rect 107712 484112 108212 484140
rect 107712 484100 107718 484112
rect 108206 484100 108212 484112
rect 108264 484100 108270 484152
rect 109034 484100 109040 484152
rect 109092 484140 109098 484152
rect 109586 484140 109592 484152
rect 109092 484112 109592 484140
rect 109092 484100 109098 484112
rect 109586 484100 109592 484112
rect 109644 484100 109650 484152
rect 116026 484100 116032 484152
rect 116084 484140 116090 484152
rect 116670 484140 116676 484152
rect 116084 484112 116676 484140
rect 116084 484100 116090 484112
rect 116670 484100 116676 484112
rect 116728 484100 116734 484152
rect 139394 484100 139400 484152
rect 139452 484140 139458 484152
rect 140038 484140 140044 484152
rect 139452 484112 140044 484140
rect 139452 484100 139458 484112
rect 140038 484100 140044 484112
rect 140096 484100 140102 484152
rect 140866 484100 140872 484152
rect 140924 484140 140930 484152
rect 141326 484140 141332 484152
rect 140924 484112 141332 484140
rect 140924 484100 140930 484112
rect 141326 484100 141332 484112
rect 141384 484100 141390 484152
rect 142154 484100 142160 484152
rect 142212 484140 142218 484152
rect 142614 484140 142620 484152
rect 142212 484112 142620 484140
rect 142212 484100 142218 484112
rect 142614 484100 142620 484112
rect 142672 484100 142678 484152
rect 143534 484100 143540 484152
rect 143592 484140 143598 484152
rect 143902 484140 143908 484152
rect 143592 484112 143908 484140
rect 143592 484100 143598 484112
rect 143902 484100 143908 484112
rect 143960 484100 143966 484152
rect 154574 484100 154580 484152
rect 154632 484140 154638 484152
rect 155402 484140 155408 484152
rect 154632 484112 155408 484140
rect 154632 484100 154638 484112
rect 155402 484100 155408 484112
rect 155460 484100 155466 484152
rect 167086 484100 167092 484152
rect 167144 484140 167150 484152
rect 167730 484140 167736 484152
rect 167144 484112 167736 484140
rect 167144 484100 167150 484112
rect 167730 484100 167736 484112
rect 167788 484100 167794 484152
rect 169846 484100 169852 484152
rect 169904 484140 169910 484152
rect 170398 484140 170404 484152
rect 169904 484112 170404 484140
rect 169904 484100 169910 484112
rect 170398 484100 170404 484112
rect 170456 484100 170462 484152
rect 171134 484100 171140 484152
rect 171192 484140 171198 484152
rect 171686 484140 171692 484152
rect 171192 484112 171692 484140
rect 171192 484100 171198 484112
rect 171686 484100 171692 484112
rect 171744 484100 171750 484152
rect 172514 484100 172520 484152
rect 172572 484140 172578 484152
rect 173526 484140 173532 484152
rect 172572 484112 173532 484140
rect 172572 484100 172578 484112
rect 173526 484100 173532 484112
rect 173584 484100 173590 484152
rect 175274 484100 175280 484152
rect 175332 484140 175338 484152
rect 176102 484140 176108 484152
rect 175332 484112 176108 484140
rect 175332 484100 175338 484112
rect 176102 484100 176108 484112
rect 176160 484100 176166 484152
rect 198734 484100 198740 484152
rect 198792 484140 198798 484152
rect 198918 484140 198924 484152
rect 198792 484112 198924 484140
rect 198792 484100 198798 484112
rect 198918 484100 198924 484112
rect 198976 484100 198982 484152
rect 200206 484100 200212 484152
rect 200264 484140 200270 484152
rect 201034 484140 201040 484152
rect 200264 484112 201040 484140
rect 200264 484100 200270 484112
rect 201034 484100 201040 484112
rect 201092 484100 201098 484152
rect 201494 484100 201500 484152
rect 201552 484140 201558 484152
rect 202046 484140 202052 484152
rect 201552 484112 202052 484140
rect 201552 484100 201558 484112
rect 202046 484100 202052 484112
rect 202104 484100 202110 484152
rect 202874 484100 202880 484152
rect 202932 484140 202938 484152
rect 203886 484140 203892 484152
rect 202932 484112 203892 484140
rect 202932 484100 202938 484112
rect 203886 484100 203892 484112
rect 203944 484100 203950 484152
rect 204346 484100 204352 484152
rect 204404 484140 204410 484152
rect 205174 484140 205180 484152
rect 204404 484112 205180 484140
rect 204404 484100 204410 484112
rect 205174 484100 205180 484112
rect 205232 484100 205238 484152
rect 205726 484100 205732 484152
rect 205784 484140 205790 484152
rect 206462 484140 206468 484152
rect 205784 484112 206468 484140
rect 205784 484100 205790 484112
rect 206462 484100 206468 484112
rect 206520 484100 206526 484152
rect 207198 484100 207204 484152
rect 207256 484140 207262 484152
rect 207566 484140 207572 484152
rect 207256 484112 207572 484140
rect 207256 484100 207262 484112
rect 207566 484100 207572 484112
rect 207624 484100 207630 484152
rect 208394 484100 208400 484152
rect 208452 484140 208458 484152
rect 209406 484140 209412 484152
rect 208452 484112 209412 484140
rect 208452 484100 208458 484112
rect 209406 484100 209412 484112
rect 209464 484100 209470 484152
rect 211246 484100 211252 484152
rect 211304 484140 211310 484152
rect 211798 484140 211804 484152
rect 211304 484112 211804 484140
rect 211304 484100 211310 484112
rect 211798 484100 211804 484112
rect 211856 484100 211862 484152
rect 212626 484100 212632 484152
rect 212684 484140 212690 484152
rect 213454 484140 213460 484152
rect 212684 484112 213460 484140
rect 212684 484100 212690 484112
rect 213454 484100 213460 484112
rect 213512 484100 213518 484152
rect 213914 484100 213920 484152
rect 213972 484140 213978 484152
rect 214926 484140 214932 484152
rect 213972 484112 214932 484140
rect 213972 484100 213978 484112
rect 214926 484100 214932 484112
rect 214984 484100 214990 484152
rect 226334 484100 226340 484152
rect 226392 484140 226398 484152
rect 226702 484140 226708 484152
rect 226392 484112 226708 484140
rect 226392 484100 226398 484112
rect 226702 484100 226708 484112
rect 226760 484100 226766 484152
rect 227806 484100 227812 484152
rect 227864 484140 227870 484152
rect 228542 484140 228548 484152
rect 227864 484112 228548 484140
rect 227864 484100 227870 484112
rect 228542 484100 228548 484112
rect 228600 484100 228606 484152
rect 231854 484100 231860 484152
rect 231912 484140 231918 484152
rect 232406 484140 232412 484152
rect 231912 484112 232412 484140
rect 231912 484100 231918 484112
rect 232406 484100 232412 484112
rect 232464 484100 232470 484152
rect 235994 484100 236000 484152
rect 236052 484140 236058 484152
rect 236822 484140 236828 484152
rect 236052 484112 236828 484140
rect 236052 484100 236058 484112
rect 236822 484100 236828 484112
rect 236880 484100 236886 484152
rect 240226 484100 240232 484152
rect 240284 484140 240290 484152
rect 240870 484140 240876 484152
rect 240284 484112 240876 484140
rect 240284 484100 240290 484112
rect 240870 484100 240876 484112
rect 240928 484100 240934 484152
rect 241514 484100 241520 484152
rect 241572 484140 241578 484152
rect 242158 484140 242164 484152
rect 241572 484112 242164 484140
rect 241572 484100 241578 484112
rect 242158 484100 242164 484112
rect 242216 484100 242222 484152
rect 263686 484100 263692 484152
rect 263744 484140 263750 484152
rect 264238 484140 264244 484152
rect 263744 484112 264244 484140
rect 263744 484100 263750 484112
rect 264238 484100 264244 484112
rect 264296 484100 264302 484152
rect 265066 484100 265072 484152
rect 265124 484140 265130 484152
rect 265894 484140 265900 484152
rect 265124 484112 265900 484140
rect 265124 484100 265130 484112
rect 265894 484100 265900 484112
rect 265952 484100 265958 484152
rect 266354 484100 266360 484152
rect 266412 484140 266418 484152
rect 266814 484140 266820 484152
rect 266412 484112 266820 484140
rect 266412 484100 266418 484112
rect 266814 484100 266820 484112
rect 266872 484100 266878 484152
rect 267734 484100 267740 484152
rect 267792 484140 267798 484152
rect 268654 484140 268660 484152
rect 267792 484112 268660 484140
rect 267792 484100 267798 484112
rect 268654 484100 268660 484112
rect 268712 484100 268718 484152
rect 269206 484100 269212 484152
rect 269264 484140 269270 484152
rect 269942 484140 269948 484152
rect 269264 484112 269948 484140
rect 269264 484100 269270 484112
rect 269942 484100 269948 484112
rect 270000 484100 270006 484152
rect 270494 484100 270500 484152
rect 270552 484140 270558 484152
rect 271230 484140 271236 484152
rect 270552 484112 271236 484140
rect 270552 484100 270558 484112
rect 271230 484100 271236 484112
rect 271288 484100 271294 484152
rect 271966 484100 271972 484152
rect 272024 484140 272030 484152
rect 272518 484140 272524 484152
rect 272024 484112 272524 484140
rect 272024 484100 272030 484112
rect 272518 484100 272524 484112
rect 272576 484100 272582 484152
rect 273254 484100 273260 484152
rect 273312 484140 273318 484152
rect 273806 484140 273812 484152
rect 273312 484112 273812 484140
rect 273312 484100 273318 484112
rect 273806 484100 273812 484112
rect 273864 484100 273870 484152
rect 274634 484100 274640 484152
rect 274692 484140 274698 484152
rect 275186 484140 275192 484152
rect 274692 484112 275192 484140
rect 274692 484100 274698 484112
rect 275186 484100 275192 484112
rect 275244 484100 275250 484152
rect 277394 484100 277400 484152
rect 277452 484140 277458 484152
rect 278222 484140 278228 484152
rect 277452 484112 278228 484140
rect 277452 484100 277458 484112
rect 278222 484100 278228 484112
rect 278280 484100 278286 484152
rect 278774 484100 278780 484152
rect 278832 484140 278838 484152
rect 279142 484140 279148 484152
rect 278832 484112 279148 484140
rect 278832 484100 278838 484112
rect 279142 484100 279148 484112
rect 279200 484100 279206 484152
rect 281626 484100 281632 484152
rect 281684 484140 281690 484152
rect 282270 484140 282276 484152
rect 281684 484112 282276 484140
rect 281684 484100 281690 484112
rect 282270 484100 282276 484112
rect 282328 484100 282334 484152
rect 282914 484100 282920 484152
rect 282972 484140 282978 484152
rect 283190 484140 283196 484152
rect 282972 484112 283196 484140
rect 282972 484100 282978 484112
rect 283190 484100 283196 484112
rect 283248 484100 283254 484152
rect 285766 484100 285772 484152
rect 285824 484140 285830 484152
rect 286686 484140 286692 484152
rect 285824 484112 286692 484140
rect 285824 484100 285830 484112
rect 286686 484100 286692 484112
rect 286744 484100 286750 484152
rect 287054 484100 287060 484152
rect 287112 484140 287118 484152
rect 287974 484140 287980 484152
rect 287112 484112 287980 484140
rect 287112 484100 287118 484112
rect 287974 484100 287980 484112
rect 288032 484100 288038 484152
rect 288434 484100 288440 484152
rect 288492 484140 288498 484152
rect 288894 484140 288900 484152
rect 288492 484112 288900 484140
rect 288492 484100 288498 484112
rect 288894 484100 288900 484112
rect 288952 484100 288958 484152
rect 289906 484100 289912 484152
rect 289964 484140 289970 484152
rect 290550 484140 290556 484152
rect 289964 484112 290556 484140
rect 289964 484100 289970 484112
rect 290550 484100 290556 484112
rect 290608 484100 290614 484152
rect 291286 484100 291292 484152
rect 291344 484140 291350 484152
rect 291470 484140 291476 484152
rect 291344 484112 291476 484140
rect 291344 484100 291350 484112
rect 291470 484100 291476 484112
rect 291528 484100 291534 484152
rect 297358 484100 297364 484152
rect 297416 484140 297422 484152
rect 379974 484140 379980 484152
rect 297416 484112 379980 484140
rect 297416 484100 297422 484112
rect 379974 484100 379980 484112
rect 380032 484100 380038 484152
rect 203794 484032 203800 484084
rect 203852 484072 203858 484084
rect 209590 484072 209596 484084
rect 203852 484044 209596 484072
rect 203852 484032 203858 484044
rect 209590 484032 209596 484044
rect 209648 484032 209654 484084
rect 257982 484032 257988 484084
rect 258040 484072 258046 484084
rect 363966 484072 363972 484084
rect 258040 484044 363972 484072
rect 258040 484032 258046 484044
rect 363966 484032 363972 484044
rect 364024 484032 364030 484084
rect 226426 483964 226432 484016
rect 226484 484004 226490 484016
rect 227254 484004 227260 484016
rect 226484 483976 227260 484004
rect 226484 483964 226490 483976
rect 227254 483964 227260 483976
rect 227312 483964 227318 484016
rect 262122 483964 262128 484016
rect 262180 484004 262186 484016
rect 376202 484004 376208 484016
rect 262180 483976 376208 484004
rect 262180 483964 262186 483976
rect 376202 483964 376208 483976
rect 376260 483964 376266 484016
rect 245194 483896 245200 483948
rect 245252 483936 245258 483948
rect 369118 483936 369124 483948
rect 245252 483908 369124 483936
rect 245252 483896 245258 483908
rect 369118 483896 369124 483908
rect 369176 483896 369182 483948
rect 248322 483828 248328 483880
rect 248380 483868 248386 483880
rect 378778 483868 378784 483880
rect 248380 483840 378784 483868
rect 248380 483828 248386 483840
rect 378778 483828 378784 483840
rect 378836 483828 378842 483880
rect 60642 483760 60648 483812
rect 60700 483800 60706 483812
rect 80698 483800 80704 483812
rect 60700 483772 80704 483800
rect 60700 483760 60706 483772
rect 80698 483760 80704 483772
rect 80756 483760 80762 483812
rect 229738 483760 229744 483812
rect 229796 483800 229802 483812
rect 363598 483800 363604 483812
rect 229796 483772 363604 483800
rect 229796 483760 229802 483772
rect 363598 483760 363604 483772
rect 363656 483760 363662 483812
rect 54754 483692 54760 483744
rect 54812 483732 54818 483744
rect 117314 483732 117320 483744
rect 54812 483704 117320 483732
rect 54812 483692 54818 483704
rect 117314 483692 117320 483704
rect 117372 483692 117378 483744
rect 176930 483692 176936 483744
rect 176988 483732 176994 483744
rect 206554 483732 206560 483744
rect 176988 483704 206560 483732
rect 176988 483692 176994 483704
rect 206554 483692 206560 483704
rect 206612 483692 206618 483744
rect 224770 483692 224776 483744
rect 224828 483732 224834 483744
rect 370498 483732 370504 483744
rect 224828 483704 370504 483732
rect 224828 483692 224834 483704
rect 370498 483692 370504 483704
rect 370556 483692 370562 483744
rect 3418 483624 3424 483676
rect 3476 483664 3482 483676
rect 316770 483664 316776 483676
rect 3476 483636 316776 483664
rect 3476 483624 3482 483636
rect 316770 483624 316776 483636
rect 316828 483624 316834 483676
rect 287422 483556 287428 483608
rect 287480 483596 287486 483608
rect 297358 483596 297364 483608
rect 287480 483568 297364 483596
rect 287480 483556 287486 483568
rect 297358 483556 297364 483568
rect 297416 483556 297422 483608
rect 113266 483352 113272 483404
rect 113324 483392 113330 483404
rect 113542 483392 113548 483404
rect 113324 483364 113548 483392
rect 113324 483352 113330 483364
rect 113542 483352 113548 483364
rect 113600 483352 113606 483404
rect 51902 482944 51908 482996
rect 51960 482984 51966 482996
rect 98454 482984 98460 482996
rect 51960 482956 98460 482984
rect 51960 482944 51966 482956
rect 98454 482944 98460 482956
rect 98512 482944 98518 482996
rect 47854 482876 47860 482928
rect 47912 482916 47918 482928
rect 97534 482916 97540 482928
rect 47912 482888 97540 482916
rect 47912 482876 47918 482888
rect 97534 482876 97540 482888
rect 97592 482876 97598 482928
rect 49234 482808 49240 482860
rect 49292 482848 49298 482860
rect 97994 482848 98000 482860
rect 49292 482820 98000 482848
rect 49292 482808 49298 482820
rect 97994 482808 98000 482820
rect 98052 482808 98058 482860
rect 46658 482740 46664 482792
rect 46716 482780 46722 482792
rect 111242 482780 111248 482792
rect 46716 482752 111248 482780
rect 46716 482740 46722 482752
rect 111242 482740 111248 482752
rect 111300 482740 111306 482792
rect 46566 482672 46572 482724
rect 46624 482712 46630 482724
rect 111702 482712 111708 482724
rect 46624 482684 111708 482712
rect 46624 482672 46630 482684
rect 111702 482672 111708 482684
rect 111760 482672 111766 482724
rect 176010 482672 176016 482724
rect 176068 482712 176074 482724
rect 210694 482712 210700 482724
rect 176068 482684 210700 482712
rect 176068 482672 176074 482684
rect 210694 482672 210700 482684
rect 210752 482672 210758 482724
rect 285122 482672 285128 482724
rect 285180 482712 285186 482724
rect 359826 482712 359832 482724
rect 285180 482684 359832 482712
rect 285180 482672 285186 482684
rect 359826 482672 359832 482684
rect 359884 482672 359890 482724
rect 49326 482604 49332 482656
rect 49384 482644 49390 482656
rect 115198 482644 115204 482656
rect 49384 482616 115204 482644
rect 49384 482604 49390 482616
rect 115198 482604 115204 482616
rect 115256 482604 115262 482656
rect 173434 482604 173440 482656
rect 173492 482644 173498 482656
rect 209038 482644 209044 482656
rect 173492 482616 209044 482644
rect 173492 482604 173498 482616
rect 209038 482604 209044 482616
rect 209096 482604 209102 482656
rect 274818 482604 274824 482656
rect 274876 482644 274882 482656
rect 361298 482644 361304 482656
rect 274876 482616 361304 482644
rect 274876 482604 274882 482616
rect 361298 482604 361304 482616
rect 361356 482604 361362 482656
rect 46382 482536 46388 482588
rect 46440 482576 46446 482588
rect 112070 482576 112076 482588
rect 46440 482548 112076 482576
rect 46440 482536 46446 482548
rect 112070 482536 112076 482548
rect 112128 482536 112134 482588
rect 138474 482536 138480 482588
rect 138532 482576 138538 482588
rect 196986 482576 196992 482588
rect 138532 482548 196992 482576
rect 138532 482536 138538 482548
rect 196986 482536 196992 482548
rect 197044 482536 197050 482588
rect 278130 482536 278136 482588
rect 278188 482576 278194 482588
rect 369578 482576 369584 482588
rect 278188 482548 369584 482576
rect 278188 482536 278194 482548
rect 369578 482536 369584 482548
rect 369636 482536 369642 482588
rect 46290 482468 46296 482520
rect 46348 482508 46354 482520
rect 112530 482508 112536 482520
rect 46348 482480 112536 482508
rect 46348 482468 46354 482480
rect 112530 482468 112536 482480
rect 112588 482468 112594 482520
rect 137186 482468 137192 482520
rect 137244 482508 137250 482520
rect 198090 482508 198096 482520
rect 137244 482480 198096 482508
rect 137244 482468 137250 482480
rect 198090 482468 198096 482480
rect 198148 482468 198154 482520
rect 277302 482468 277308 482520
rect 277360 482508 277366 482520
rect 368290 482508 368296 482520
rect 277360 482480 368296 482508
rect 277360 482468 277366 482480
rect 368290 482468 368296 482480
rect 368348 482468 368354 482520
rect 46842 482400 46848 482452
rect 46900 482440 46906 482452
rect 115658 482440 115664 482452
rect 46900 482412 115664 482440
rect 46900 482400 46906 482412
rect 115658 482400 115664 482412
rect 115716 482400 115722 482452
rect 138842 482400 138848 482452
rect 138900 482440 138906 482452
rect 200390 482440 200396 482452
rect 138900 482412 200396 482440
rect 138900 482400 138906 482412
rect 200390 482400 200396 482412
rect 200448 482400 200454 482452
rect 257706 482400 257712 482452
rect 257764 482440 257770 482452
rect 362586 482440 362592 482452
rect 257764 482412 362592 482440
rect 257764 482400 257770 482412
rect 362586 482400 362592 482412
rect 362644 482400 362650 482452
rect 45922 482332 45928 482384
rect 45980 482372 45986 482384
rect 119614 482372 119620 482384
rect 45980 482344 119620 482372
rect 45980 482332 45986 482344
rect 119614 482332 119620 482344
rect 119672 482332 119678 482384
rect 136542 482332 136548 482384
rect 136600 482372 136606 482384
rect 203150 482372 203156 482384
rect 136600 482344 203156 482372
rect 136600 482332 136606 482344
rect 203150 482332 203156 482344
rect 203208 482332 203214 482384
rect 261754 482332 261760 482384
rect 261812 482372 261818 482384
rect 373534 482372 373540 482384
rect 261812 482344 373540 482372
rect 261812 482332 261818 482344
rect 373534 482332 373540 482344
rect 373592 482332 373598 482384
rect 50154 482264 50160 482316
rect 50212 482304 50218 482316
rect 131114 482304 131120 482316
rect 50212 482276 131120 482304
rect 50212 482264 50218 482276
rect 131114 482264 131120 482276
rect 131172 482264 131178 482316
rect 136266 482264 136272 482316
rect 136324 482304 136330 482316
rect 204530 482304 204536 482316
rect 136324 482276 204536 482304
rect 136324 482264 136330 482276
rect 204530 482264 204536 482276
rect 204588 482264 204594 482316
rect 245010 482264 245016 482316
rect 245068 482304 245074 482316
rect 360930 482304 360936 482316
rect 245068 482276 360936 482304
rect 245068 482264 245074 482276
rect 360930 482264 360936 482276
rect 360988 482264 360994 482316
rect 50430 482196 50436 482248
rect 50488 482236 50494 482248
rect 97166 482236 97172 482248
rect 50488 482208 97172 482236
rect 50488 482196 50494 482208
rect 97166 482196 97172 482208
rect 97224 482196 97230 482248
rect 54662 482128 54668 482180
rect 54720 482168 54726 482180
rect 96706 482168 96712 482180
rect 54720 482140 96712 482168
rect 54720 482128 54726 482140
rect 96706 482128 96712 482140
rect 96764 482128 96770 482180
rect 58802 482060 58808 482112
rect 58860 482100 58866 482112
rect 96246 482100 96252 482112
rect 58860 482072 96252 482100
rect 58860 482060 58866 482072
rect 96246 482060 96252 482072
rect 96304 482060 96310 482112
rect 127158 482060 127164 482112
rect 127216 482100 127222 482112
rect 127342 482100 127348 482112
rect 127216 482072 127348 482100
rect 127216 482060 127222 482072
rect 127342 482060 127348 482072
rect 127400 482060 127406 482112
rect 182358 481312 182364 481364
rect 182416 481312 182422 481364
rect 283006 481312 283012 481364
rect 283064 481352 283070 481364
rect 283558 481352 283564 481364
rect 283064 481324 283564 481352
rect 283064 481312 283070 481324
rect 283558 481312 283564 481324
rect 283616 481312 283622 481364
rect 294046 481312 294052 481364
rect 294104 481352 294110 481364
rect 294230 481352 294236 481364
rect 294104 481324 294236 481352
rect 294104 481312 294110 481324
rect 294230 481312 294236 481324
rect 294288 481312 294294 481364
rect 182376 481160 182404 481312
rect 281442 481244 281448 481296
rect 281500 481284 281506 481296
rect 370406 481284 370412 481296
rect 281500 481256 370412 481284
rect 281500 481244 281506 481256
rect 370406 481244 370412 481256
rect 370464 481244 370470 481296
rect 192110 481176 192116 481228
rect 192168 481216 192174 481228
rect 192294 481216 192300 481228
rect 192168 481188 192300 481216
rect 192168 481176 192174 481188
rect 192294 481176 192300 481188
rect 192352 481176 192358 481228
rect 281074 481176 281080 481228
rect 281132 481216 281138 481228
rect 376478 481216 376484 481228
rect 281132 481188 376484 481216
rect 281132 481176 281138 481188
rect 376478 481176 376484 481188
rect 376536 481176 376542 481228
rect 180886 481108 180892 481160
rect 180944 481148 180950 481160
rect 181070 481148 181076 481160
rect 180944 481120 181076 481148
rect 180944 481108 180950 481120
rect 181070 481108 181076 481120
rect 181128 481108 181134 481160
rect 182358 481108 182364 481160
rect 182416 481108 182422 481160
rect 189350 481108 189356 481160
rect 189408 481148 189414 481160
rect 203886 481148 203892 481160
rect 189408 481120 203892 481148
rect 189408 481108 189414 481120
rect 203886 481108 203892 481120
rect 203944 481108 203950 481160
rect 251174 481108 251180 481160
rect 251232 481148 251238 481160
rect 251358 481148 251364 481160
rect 251232 481120 251364 481148
rect 251232 481108 251238 481120
rect 251358 481108 251364 481120
rect 251416 481108 251422 481160
rect 261202 481108 261208 481160
rect 261260 481148 261266 481160
rect 366726 481148 366732 481160
rect 261260 481120 366732 481148
rect 261260 481108 261266 481120
rect 366726 481108 366732 481120
rect 366784 481108 366790 481160
rect 180518 481040 180524 481092
rect 180576 481080 180582 481092
rect 214834 481080 214840 481092
rect 180576 481052 214840 481080
rect 180576 481040 180582 481052
rect 214834 481040 214840 481052
rect 214892 481040 214898 481092
rect 243078 481040 243084 481092
rect 243136 481080 243142 481092
rect 365070 481080 365076 481092
rect 243136 481052 365076 481080
rect 243136 481040 243142 481052
rect 365070 481040 365076 481052
rect 365128 481040 365134 481092
rect 56870 480972 56876 481024
rect 56928 481012 56934 481024
rect 114278 481012 114284 481024
rect 56928 480984 114284 481012
rect 56928 480972 56934 480984
rect 114278 480972 114284 480984
rect 114336 480972 114342 481024
rect 158714 480972 158720 481024
rect 158772 481012 158778 481024
rect 159358 481012 159364 481024
rect 158772 480984 159364 481012
rect 158772 480972 158778 480984
rect 159358 480972 159364 480984
rect 159416 480972 159422 481024
rect 160278 480972 160284 481024
rect 160336 481012 160342 481024
rect 210418 481012 210424 481024
rect 160336 480984 210424 481012
rect 160336 480972 160342 480984
rect 210418 480972 210424 480984
rect 210476 480972 210482 481024
rect 229554 480972 229560 481024
rect 229612 481012 229618 481024
rect 360838 481012 360844 481024
rect 229612 480984 360844 481012
rect 229612 480972 229618 480984
rect 360838 480972 360844 480984
rect 360896 480972 360902 481024
rect 3602 480904 3608 480956
rect 3660 480944 3666 480956
rect 429286 480944 429292 480956
rect 3660 480916 429292 480944
rect 3660 480904 3666 480916
rect 429286 480904 429292 480916
rect 429344 480904 429350 480956
rect 82814 480836 82820 480888
rect 82872 480876 82878 480888
rect 83550 480876 83556 480888
rect 82872 480848 83556 480876
rect 82872 480836 82878 480848
rect 83550 480836 83556 480848
rect 83608 480836 83614 480888
rect 85574 480836 85580 480888
rect 85632 480876 85638 480888
rect 86310 480876 86316 480888
rect 85632 480848 86316 480876
rect 85632 480836 85638 480848
rect 86310 480836 86316 480848
rect 86368 480836 86374 480888
rect 126974 480836 126980 480888
rect 127032 480876 127038 480888
rect 127710 480876 127716 480888
rect 127032 480848 127716 480876
rect 127032 480836 127038 480848
rect 127710 480836 127716 480848
rect 127768 480836 127774 480888
rect 158806 480836 158812 480888
rect 158864 480876 158870 480888
rect 158990 480876 158996 480888
rect 158864 480848 158996 480876
rect 158864 480836 158870 480848
rect 158990 480836 158996 480848
rect 159048 480836 159054 480888
rect 160094 480836 160100 480888
rect 160152 480876 160158 480888
rect 160646 480876 160652 480888
rect 160152 480848 160652 480876
rect 160152 480836 160158 480848
rect 160646 480836 160652 480848
rect 160704 480836 160710 480888
rect 161566 480836 161572 480888
rect 161624 480876 161630 480888
rect 162486 480876 162492 480888
rect 161624 480848 162492 480876
rect 161624 480836 161630 480848
rect 162486 480836 162492 480848
rect 162544 480836 162550 480888
rect 179414 480836 179420 480888
rect 179472 480876 179478 480888
rect 179598 480876 179604 480888
rect 179472 480848 179604 480876
rect 179472 480836 179478 480848
rect 179598 480836 179604 480848
rect 179656 480836 179662 480888
rect 182266 480836 182272 480888
rect 182324 480876 182330 480888
rect 183094 480876 183100 480888
rect 182324 480848 183100 480876
rect 182324 480836 182330 480848
rect 183094 480836 183100 480848
rect 183152 480836 183158 480888
rect 183646 480836 183652 480888
rect 183704 480876 183710 480888
rect 184014 480876 184020 480888
rect 183704 480848 184020 480876
rect 183704 480836 183710 480848
rect 184014 480836 184020 480848
rect 184072 480836 184078 480888
rect 184934 480836 184940 480888
rect 184992 480876 184998 480888
rect 185854 480876 185860 480888
rect 184992 480848 185860 480876
rect 184992 480836 184998 480848
rect 185854 480836 185860 480848
rect 185912 480836 185918 480888
rect 187694 480836 187700 480888
rect 187752 480876 187758 480888
rect 188430 480876 188436 480888
rect 187752 480848 188436 480876
rect 187752 480836 187758 480848
rect 188430 480836 188436 480848
rect 188488 480836 188494 480888
rect 191926 480836 191932 480888
rect 191984 480876 191990 480888
rect 192386 480876 192392 480888
rect 191984 480848 192392 480876
rect 191984 480836 191990 480848
rect 192386 480836 192392 480848
rect 192444 480836 192450 480888
rect 193306 480836 193312 480888
rect 193364 480876 193370 480888
rect 193766 480876 193772 480888
rect 193364 480848 193772 480876
rect 193364 480836 193370 480848
rect 193766 480836 193772 480848
rect 193824 480836 193830 480888
rect 245654 480836 245660 480888
rect 245712 480876 245718 480888
rect 246574 480876 246580 480888
rect 245712 480848 246580 480876
rect 245712 480836 245718 480848
rect 246574 480836 246580 480848
rect 246632 480836 246638 480888
rect 248414 480836 248420 480888
rect 248472 480876 248478 480888
rect 249150 480876 249156 480888
rect 248472 480848 249156 480876
rect 248472 480836 248478 480848
rect 249150 480836 249156 480848
rect 249208 480836 249214 480888
rect 251266 480836 251272 480888
rect 251324 480876 251330 480888
rect 251910 480876 251916 480888
rect 251324 480848 251916 480876
rect 251324 480836 251330 480848
rect 251910 480836 251916 480848
rect 251968 480836 251974 480888
rect 252646 480836 252652 480888
rect 252704 480876 252710 480888
rect 253198 480876 253204 480888
rect 252704 480848 253204 480876
rect 252704 480836 252710 480848
rect 253198 480836 253204 480848
rect 253256 480836 253262 480888
rect 253934 480836 253940 480888
rect 253992 480876 253998 480888
rect 254486 480876 254492 480888
rect 253992 480848 254492 480876
rect 253992 480836 253998 480848
rect 254486 480836 254492 480848
rect 254544 480836 254550 480888
rect 259454 480836 259460 480888
rect 259512 480876 259518 480888
rect 259638 480876 259644 480888
rect 259512 480848 259644 480876
rect 259512 480836 259518 480848
rect 259638 480836 259644 480848
rect 259696 480836 259702 480888
rect 262214 480836 262220 480888
rect 262272 480876 262278 480888
rect 262398 480876 262404 480888
rect 262272 480848 262404 480876
rect 262272 480836 262278 480848
rect 262398 480836 262404 480848
rect 262456 480836 262462 480888
rect 295426 480836 295432 480888
rect 295484 480876 295490 480888
rect 295886 480876 295892 480888
rect 295484 480848 295892 480876
rect 295484 480836 295490 480848
rect 295886 480836 295892 480848
rect 295944 480836 295950 480888
rect 296714 480836 296720 480888
rect 296772 480876 296778 480888
rect 297726 480876 297732 480888
rect 296772 480848 297732 480876
rect 296772 480836 296778 480848
rect 297726 480836 297732 480848
rect 297784 480836 297790 480888
rect 298094 480836 298100 480888
rect 298152 480876 298158 480888
rect 298462 480876 298468 480888
rect 298152 480848 298468 480876
rect 298152 480836 298158 480848
rect 298462 480836 298468 480848
rect 298520 480836 298526 480888
rect 183554 480768 183560 480820
rect 183612 480808 183618 480820
rect 184382 480808 184388 480820
rect 183612 480780 184388 480808
rect 183612 480768 183618 480780
rect 184382 480768 184388 480780
rect 184440 480768 184446 480820
rect 192018 480768 192024 480820
rect 192076 480808 192082 480820
rect 192846 480808 192852 480820
rect 192076 480780 192852 480808
rect 192076 480768 192082 480780
rect 192846 480768 192852 480780
rect 192904 480768 192910 480820
rect 193214 480768 193220 480820
rect 193272 480808 193278 480820
rect 194134 480808 194140 480820
rect 193272 480780 194140 480808
rect 193272 480768 193278 480780
rect 194134 480768 194140 480780
rect 194192 480768 194198 480820
rect 88426 480564 88432 480616
rect 88484 480604 88490 480616
rect 89254 480604 89260 480616
rect 88484 480576 89260 480604
rect 88484 480564 88490 480576
rect 89254 480564 89260 480576
rect 89312 480564 89318 480616
rect 70486 480360 70492 480412
rect 70544 480400 70550 480412
rect 71222 480400 71228 480412
rect 70544 480372 71228 480400
rect 70544 480360 70550 480372
rect 71222 480360 71228 480372
rect 71280 480360 71286 480412
rect 292666 480292 292672 480344
rect 292724 480332 292730 480344
rect 293310 480332 293316 480344
rect 292724 480304 293316 480332
rect 292724 480292 292730 480304
rect 293310 480292 293316 480304
rect 293368 480292 293374 480344
rect 220814 480224 220820 480276
rect 220872 480264 220878 480276
rect 220998 480264 221004 480276
rect 220872 480236 221004 480264
rect 220872 480224 220878 480236
rect 220998 480224 221004 480236
rect 221056 480224 221062 480276
rect 59722 480156 59728 480208
rect 59780 480196 59786 480208
rect 130286 480196 130292 480208
rect 59780 480168 130292 480196
rect 59780 480156 59786 480168
rect 130286 480156 130292 480168
rect 130344 480156 130350 480208
rect 45462 480088 45468 480140
rect 45520 480128 45526 480140
rect 118878 480128 118884 480140
rect 45520 480100 118884 480128
rect 45520 480088 45526 480100
rect 118878 480088 118884 480100
rect 118936 480088 118942 480140
rect 43898 480020 43904 480072
rect 43956 480060 43962 480072
rect 117958 480060 117964 480072
rect 43956 480032 117964 480060
rect 43956 480020 43962 480032
rect 117958 480020 117964 480032
rect 118016 480020 118022 480072
rect 294598 480020 294604 480072
rect 294656 480060 294662 480072
rect 371694 480060 371700 480072
rect 294656 480032 371700 480060
rect 294656 480020 294662 480032
rect 371694 480020 371700 480032
rect 371752 480020 371758 480072
rect 43806 479952 43812 480004
rect 43864 479992 43870 480004
rect 117406 479992 117412 480004
rect 43864 479964 117412 479992
rect 43864 479952 43870 479964
rect 117406 479952 117412 479964
rect 117464 479952 117470 480004
rect 278866 479952 278872 480004
rect 278924 479992 278930 480004
rect 361390 479992 361396 480004
rect 278924 479964 361396 479992
rect 278924 479952 278930 479964
rect 361390 479952 361396 479964
rect 361448 479952 361454 480004
rect 58618 479884 58624 479936
rect 58676 479924 58682 479936
rect 132770 479924 132776 479936
rect 58676 479896 132776 479924
rect 58676 479884 58682 479896
rect 132770 479884 132776 479896
rect 132828 479884 132834 479936
rect 275646 479884 275652 479936
rect 275704 479924 275710 479936
rect 372430 479924 372436 479936
rect 275704 479896 372436 479924
rect 275704 479884 275710 479896
rect 372430 479884 372436 479896
rect 372488 479884 372494 479936
rect 53558 479816 53564 479868
rect 53616 479856 53622 479868
rect 131574 479856 131580 479868
rect 53616 479828 131580 479856
rect 53616 479816 53622 479828
rect 131574 479816 131580 479828
rect 131632 479816 131638 479868
rect 272058 479816 272064 479868
rect 272116 479856 272122 479868
rect 370314 479856 370320 479868
rect 272116 479828 370320 479856
rect 272116 479816 272122 479828
rect 370314 479816 370320 479828
rect 370372 479816 370378 479868
rect 57330 479748 57336 479800
rect 57388 479788 57394 479800
rect 135254 479788 135260 479800
rect 57388 479760 135260 479788
rect 57388 479748 57394 479760
rect 135254 479748 135260 479760
rect 135312 479748 135318 479800
rect 161658 479748 161664 479800
rect 161716 479788 161722 479800
rect 161934 479788 161940 479800
rect 161716 479760 161940 479788
rect 161716 479748 161722 479760
rect 161934 479748 161940 479760
rect 161992 479748 161998 479800
rect 255774 479748 255780 479800
rect 255832 479788 255838 479800
rect 356882 479788 356888 479800
rect 255832 479760 356888 479788
rect 255832 479748 255838 479760
rect 356882 479748 356888 479760
rect 356940 479748 356946 479800
rect 42518 479680 42524 479732
rect 42576 479720 42582 479732
rect 123018 479720 123024 479732
rect 42576 479692 123024 479720
rect 42576 479680 42582 479692
rect 123018 479680 123024 479692
rect 123076 479680 123082 479732
rect 190546 479680 190552 479732
rect 190604 479720 190610 479732
rect 191006 479720 191012 479732
rect 190604 479692 191012 479720
rect 190604 479680 190610 479692
rect 191006 479680 191012 479692
rect 191064 479680 191070 479732
rect 256694 479680 256700 479732
rect 256752 479720 256758 479732
rect 361022 479720 361028 479732
rect 256752 479692 361028 479720
rect 256752 479680 256758 479692
rect 361022 479680 361028 479692
rect 361080 479680 361086 479732
rect 49050 479612 49056 479664
rect 49108 479652 49114 479664
rect 130654 479652 130660 479664
rect 49108 479624 130660 479652
rect 49108 479612 49114 479624
rect 130654 479612 130660 479624
rect 130712 479612 130718 479664
rect 258442 479612 258448 479664
rect 258500 479652 258506 479664
rect 370866 479652 370872 479664
rect 258500 479624 370872 479652
rect 258500 479612 258506 479624
rect 370866 479612 370872 479624
rect 370924 479612 370930 479664
rect 47762 479544 47768 479596
rect 47820 479584 47826 479596
rect 129918 479584 129924 479596
rect 47820 479556 129924 479584
rect 47820 479544 47826 479556
rect 129918 479544 129924 479556
rect 129976 479544 129982 479596
rect 178310 479544 178316 479596
rect 178368 479584 178374 479596
rect 200758 479584 200764 479596
rect 178368 479556 200764 479584
rect 178368 479544 178374 479556
rect 200758 479544 200764 479556
rect 200816 479544 200822 479596
rect 245930 479544 245936 479596
rect 245988 479584 245994 479596
rect 371970 479584 371976 479596
rect 245988 479556 371976 479584
rect 245988 479544 245994 479556
rect 371970 479544 371976 479556
rect 372028 479544 372034 479596
rect 46106 479476 46112 479528
rect 46164 479516 46170 479528
rect 128906 479516 128912 479528
rect 46164 479488 128912 479516
rect 46164 479476 46170 479488
rect 128906 479476 128912 479488
rect 128964 479476 128970 479528
rect 163038 479476 163044 479528
rect 163096 479516 163102 479528
rect 206370 479516 206376 479528
rect 163096 479488 206376 479516
rect 163096 479476 163102 479488
rect 206370 479476 206376 479488
rect 206428 479476 206434 479528
rect 236454 479476 236460 479528
rect 236512 479516 236518 479528
rect 363782 479516 363788 479528
rect 236512 479488 363788 479516
rect 236512 479476 236518 479488
rect 363782 479476 363788 479488
rect 363840 479476 363846 479528
rect 46474 479408 46480 479460
rect 46532 479448 46538 479460
rect 116026 479448 116032 479460
rect 46532 479420 116032 479448
rect 46532 479408 46538 479420
rect 116026 479408 116032 479420
rect 116084 479408 116090 479460
rect 259454 479408 259460 479460
rect 259512 479448 259518 479460
rect 260190 479448 260196 479460
rect 259512 479420 260196 479448
rect 259512 479408 259518 479420
rect 260190 479408 260196 479420
rect 260248 479408 260254 479460
rect 47946 479340 47952 479392
rect 48004 479380 48010 479392
rect 116118 479380 116124 479392
rect 48004 479352 116124 479380
rect 48004 479340 48010 479352
rect 116118 479340 116124 479352
rect 116176 479340 116182 479392
rect 50338 479272 50344 479324
rect 50396 479312 50402 479324
rect 115934 479312 115940 479324
rect 50396 479284 115940 479312
rect 50396 479272 50402 479284
rect 115934 479272 115940 479284
rect 115992 479272 115998 479324
rect 269206 478456 269212 478508
rect 269264 478496 269270 478508
rect 357066 478496 357072 478508
rect 269264 478468 357072 478496
rect 269264 478456 269270 478468
rect 357066 478456 357072 478468
rect 357124 478456 357130 478508
rect 269390 478388 269396 478440
rect 269448 478428 269454 478440
rect 359458 478428 359464 478440
rect 269448 478400 359464 478428
rect 269448 478388 269454 478400
rect 359458 478388 359464 478400
rect 359516 478388 359522 478440
rect 186406 478320 186412 478372
rect 186464 478360 186470 478372
rect 216030 478360 216036 478372
rect 186464 478332 216036 478360
rect 186464 478320 186470 478332
rect 216030 478320 216036 478332
rect 216088 478320 216094 478372
rect 270862 478320 270868 478372
rect 270920 478360 270926 478372
rect 373166 478360 373172 478372
rect 270920 478332 373172 478360
rect 270920 478320 270926 478332
rect 373166 478320 373172 478332
rect 373224 478320 373230 478372
rect 177022 478252 177028 478304
rect 177080 478292 177086 478304
rect 209222 478292 209228 478304
rect 177080 478264 209228 478292
rect 177080 478252 177086 478264
rect 209222 478252 209228 478264
rect 209280 478252 209286 478304
rect 270586 478252 270592 478304
rect 270644 478292 270650 478304
rect 377306 478292 377312 478304
rect 270644 478264 377312 478292
rect 270644 478252 270650 478264
rect 377306 478252 377312 478264
rect 377364 478252 377370 478304
rect 85666 478184 85672 478236
rect 85724 478224 85730 478236
rect 85850 478224 85856 478236
rect 85724 478196 85856 478224
rect 85724 478184 85730 478196
rect 85850 478184 85856 478196
rect 85908 478184 85914 478236
rect 165062 478184 165068 478236
rect 165120 478224 165126 478236
rect 211890 478224 211896 478236
rect 165120 478196 211896 478224
rect 165120 478184 165126 478196
rect 211890 478184 211896 478196
rect 211948 478184 211954 478236
rect 247402 478184 247408 478236
rect 247460 478224 247466 478236
rect 376018 478224 376024 478236
rect 247460 478196 376024 478224
rect 247460 478184 247466 478196
rect 376018 478184 376024 478196
rect 376076 478184 376082 478236
rect 62298 478116 62304 478168
rect 62356 478156 62362 478168
rect 199286 478156 199292 478168
rect 62356 478128 199292 478156
rect 62356 478116 62362 478128
rect 199286 478116 199292 478128
rect 199344 478116 199350 478168
rect 238202 478116 238208 478168
rect 238260 478156 238266 478168
rect 378870 478156 378876 478168
rect 238260 478128 378876 478156
rect 238260 478116 238266 478128
rect 378870 478116 378876 478128
rect 378928 478116 378934 478168
rect 49142 477436 49148 477488
rect 49200 477476 49206 477488
rect 125594 477476 125600 477488
rect 49200 477448 125600 477476
rect 49200 477436 49206 477448
rect 125594 477436 125600 477448
rect 125652 477436 125658 477488
rect 291286 477436 291292 477488
rect 291344 477476 291350 477488
rect 362770 477476 362776 477488
rect 291344 477448 362776 477476
rect 291344 477436 291350 477448
rect 362770 477436 362776 477448
rect 362828 477436 362834 477488
rect 56594 477368 56600 477420
rect 56652 477408 56658 477420
rect 134702 477408 134708 477420
rect 56652 477380 134708 477408
rect 56652 477368 56658 477380
rect 134702 477368 134708 477380
rect 134760 477368 134766 477420
rect 291378 477368 291384 477420
rect 291436 477408 291442 477420
rect 368382 477408 368388 477420
rect 291436 477380 368388 477408
rect 291436 477368 291442 477380
rect 368382 477368 368388 477380
rect 368440 477368 368446 477420
rect 42610 477300 42616 477352
rect 42668 477340 42674 477352
rect 120534 477340 120540 477352
rect 42668 477312 120540 477340
rect 42668 477300 42674 477312
rect 120534 477300 120540 477312
rect 120592 477300 120598 477352
rect 278774 477300 278780 477352
rect 278832 477340 278838 477352
rect 364150 477340 364156 477352
rect 278832 477312 364156 477340
rect 278832 477300 278838 477312
rect 364150 477300 364156 477312
rect 364208 477300 364214 477352
rect 43990 477232 43996 477284
rect 44048 477272 44054 477284
rect 123294 477272 123300 477284
rect 44048 477244 123300 477272
rect 44048 477232 44054 477244
rect 123294 477232 123300 477244
rect 123352 477232 123358 477284
rect 274726 477232 274732 477284
rect 274784 477272 274790 477284
rect 364242 477272 364248 477284
rect 274784 477244 364248 477272
rect 274784 477232 274790 477244
rect 364242 477232 364248 477244
rect 364300 477232 364306 477284
rect 42426 477164 42432 477216
rect 42484 477204 42490 477216
rect 121546 477204 121552 477216
rect 42484 477176 121552 477204
rect 42484 477164 42490 477176
rect 121546 477164 121552 477176
rect 121604 477164 121610 477216
rect 263686 477164 263692 477216
rect 263744 477204 263750 477216
rect 366818 477204 366824 477216
rect 263744 477176 366824 477204
rect 263744 477164 263750 477176
rect 366818 477164 366824 477176
rect 366876 477164 366882 477216
rect 43622 477096 43628 477148
rect 43680 477136 43686 477148
rect 124950 477136 124956 477148
rect 43680 477108 124956 477136
rect 43680 477096 43686 477108
rect 124950 477096 124956 477108
rect 125008 477096 125014 477148
rect 258902 477096 258908 477148
rect 258960 477136 258966 477148
rect 365346 477136 365352 477148
rect 258960 477108 365352 477136
rect 258960 477096 258966 477108
rect 365346 477096 365352 477108
rect 365404 477096 365410 477148
rect 43714 477028 43720 477080
rect 43772 477068 43778 477080
rect 125870 477068 125876 477080
rect 43772 477040 125876 477068
rect 43772 477028 43778 477040
rect 125870 477028 125876 477040
rect 125928 477028 125934 477080
rect 254854 477028 254860 477080
rect 254912 477068 254918 477080
rect 365438 477068 365444 477080
rect 254912 477040 365444 477068
rect 254912 477028 254918 477040
rect 365438 477028 365444 477040
rect 365496 477028 365502 477080
rect 48958 476960 48964 477012
rect 49016 477000 49022 477012
rect 133414 477000 133420 477012
rect 49016 476972 133420 477000
rect 49016 476960 49022 476972
rect 133414 476960 133420 476972
rect 133472 476960 133478 477012
rect 263778 476960 263784 477012
rect 263836 477000 263842 477012
rect 376294 477000 376300 477012
rect 263836 476972 376300 477000
rect 263836 476960 263842 476972
rect 376294 476960 376300 476972
rect 376352 476960 376358 477012
rect 47670 476892 47676 476944
rect 47728 476932 47734 476944
rect 132862 476932 132868 476944
rect 47728 476904 132868 476932
rect 47728 476892 47734 476904
rect 132862 476892 132868 476904
rect 132920 476892 132926 476944
rect 185026 476892 185032 476944
rect 185084 476932 185090 476944
rect 212074 476932 212080 476944
rect 185084 476904 212080 476932
rect 185084 476892 185090 476904
rect 212074 476892 212080 476904
rect 212132 476892 212138 476944
rect 241698 476892 241704 476944
rect 241756 476932 241762 476944
rect 367830 476932 367836 476944
rect 241756 476904 367836 476932
rect 241756 476892 241762 476904
rect 367830 476892 367836 476904
rect 367888 476892 367894 476944
rect 43254 476824 43260 476876
rect 43312 476864 43318 476876
rect 143626 476864 143632 476876
rect 43312 476836 143632 476864
rect 43312 476824 43318 476836
rect 143626 476824 143632 476836
rect 143684 476824 143690 476876
rect 150434 476824 150440 476876
rect 150492 476864 150498 476876
rect 211798 476864 211804 476876
rect 150492 476836 211804 476864
rect 150492 476824 150498 476836
rect 211798 476824 211804 476836
rect 211856 476824 211862 476876
rect 238754 476824 238760 476876
rect 238812 476864 238818 476876
rect 373258 476864 373264 476876
rect 238812 476836 373264 476864
rect 238812 476824 238818 476836
rect 373258 476824 373264 476836
rect 373316 476824 373322 476876
rect 62206 476756 62212 476808
rect 62264 476796 62270 476808
rect 199378 476796 199384 476808
rect 62264 476768 199384 476796
rect 62264 476756 62270 476768
rect 199378 476756 199384 476768
rect 199436 476756 199442 476808
rect 204438 476756 204444 476808
rect 204496 476796 204502 476808
rect 217318 476796 217324 476808
rect 204496 476768 217324 476796
rect 204496 476756 204502 476768
rect 217318 476756 217324 476768
rect 217376 476756 217382 476808
rect 237466 476756 237472 476808
rect 237524 476796 237530 476808
rect 376110 476796 376116 476808
rect 237524 476768 376116 476796
rect 237524 476756 237530 476768
rect 376110 476756 376116 476768
rect 376168 476756 376174 476808
rect 57054 476688 57060 476740
rect 57112 476728 57118 476740
rect 128630 476728 128636 476740
rect 57112 476700 128636 476728
rect 57112 476688 57118 476700
rect 128630 476688 128636 476700
rect 128688 476688 128694 476740
rect 58434 476620 58440 476672
rect 58492 476660 58498 476672
rect 128354 476660 128360 476672
rect 58492 476632 128360 476660
rect 58492 476620 58498 476632
rect 128354 476620 128360 476632
rect 128412 476620 128418 476672
rect 290182 475600 290188 475652
rect 290240 475640 290246 475652
rect 363506 475640 363512 475652
rect 290240 475612 363512 475640
rect 290240 475600 290246 475612
rect 363506 475600 363512 475612
rect 363564 475600 363570 475652
rect 292758 475532 292764 475584
rect 292816 475572 292822 475584
rect 376754 475572 376760 475584
rect 292816 475544 376760 475572
rect 292816 475532 292822 475544
rect 376754 475532 376760 475544
rect 376812 475532 376818 475584
rect 270494 475464 270500 475516
rect 270552 475504 270558 475516
rect 375282 475504 375288 475516
rect 270552 475476 375288 475504
rect 270552 475464 270558 475476
rect 375282 475464 375288 475476
rect 375340 475464 375346 475516
rect 176654 475396 176660 475448
rect 176712 475436 176718 475448
rect 205082 475436 205088 475448
rect 176712 475408 205088 475436
rect 176712 475396 176718 475408
rect 205082 475396 205088 475408
rect 205140 475396 205146 475448
rect 207658 475396 207664 475448
rect 207716 475436 207722 475448
rect 217686 475436 217692 475448
rect 207716 475408 217692 475436
rect 207716 475396 207722 475408
rect 217686 475396 217692 475408
rect 217744 475396 217750 475448
rect 259638 475396 259644 475448
rect 259696 475436 259702 475448
rect 372154 475436 372160 475448
rect 259696 475408 372160 475436
rect 259696 475396 259702 475408
rect 372154 475396 372160 475408
rect 372212 475396 372218 475448
rect 164234 475328 164240 475380
rect 164292 475368 164298 475380
rect 218790 475368 218796 475380
rect 164292 475340 218796 475368
rect 164292 475328 164298 475340
rect 218790 475328 218796 475340
rect 218848 475328 218854 475380
rect 245746 475328 245752 475380
rect 245804 475368 245810 475380
rect 362402 475368 362408 475380
rect 245804 475340 362408 475368
rect 245804 475328 245810 475340
rect 362402 475328 362408 475340
rect 362460 475328 362466 475380
rect 182174 474784 182180 474836
rect 182232 474824 182238 474836
rect 182450 474824 182456 474836
rect 182232 474796 182456 474824
rect 182232 474784 182238 474796
rect 182450 474784 182456 474796
rect 182508 474784 182514 474836
rect 276014 474648 276020 474700
rect 276072 474688 276078 474700
rect 357250 474688 357256 474700
rect 276072 474660 357256 474688
rect 276072 474648 276078 474660
rect 357250 474648 357256 474660
rect 357308 474648 357314 474700
rect 47578 474580 47584 474632
rect 47636 474620 47642 474632
rect 65518 474620 65524 474632
rect 47636 474592 65524 474620
rect 47636 474580 47642 474592
rect 65518 474580 65524 474592
rect 65576 474580 65582 474632
rect 271966 474580 271972 474632
rect 272024 474620 272030 474632
rect 367554 474620 367560 474632
rect 272024 474592 367560 474620
rect 272024 474580 272030 474592
rect 367554 474580 367560 474592
rect 367612 474580 367618 474632
rect 45094 474512 45100 474564
rect 45152 474552 45158 474564
rect 68278 474552 68284 474564
rect 45152 474524 68284 474552
rect 45152 474512 45158 474524
rect 68278 474512 68284 474524
rect 68336 474512 68342 474564
rect 263594 474512 263600 474564
rect 263652 474552 263658 474564
rect 364058 474552 364064 474564
rect 263652 474524 364064 474552
rect 263652 474512 263658 474524
rect 364058 474512 364064 474524
rect 364116 474512 364122 474564
rect 43530 474444 43536 474496
rect 43588 474484 43594 474496
rect 68370 474484 68376 474496
rect 43588 474456 68376 474484
rect 43588 474444 43594 474456
rect 68370 474444 68376 474456
rect 68428 474444 68434 474496
rect 268102 474444 268108 474496
rect 268160 474484 268166 474496
rect 375098 474484 375104 474496
rect 268160 474456 375104 474484
rect 268160 474444 268166 474456
rect 375098 474444 375104 474456
rect 375156 474444 375162 474496
rect 57422 474376 57428 474428
rect 57480 474416 57486 474428
rect 103606 474416 103612 474428
rect 57480 474388 103612 474416
rect 57480 474376 57486 474388
rect 103606 474376 103612 474388
rect 103664 474376 103670 474428
rect 251358 474376 251364 474428
rect 251416 474416 251422 474428
rect 366634 474416 366640 474428
rect 251416 474388 366640 474416
rect 251416 474376 251422 474388
rect 366634 474376 366640 474388
rect 366692 474376 366698 474428
rect 51810 474308 51816 474360
rect 51868 474348 51874 474360
rect 99558 474348 99564 474360
rect 51868 474320 99564 474348
rect 51868 474308 51874 474320
rect 99558 474308 99564 474320
rect 99616 474308 99622 474360
rect 188062 474308 188068 474360
rect 188120 474348 188126 474360
rect 207750 474348 207756 474360
rect 188120 474320 207756 474348
rect 188120 474308 188126 474320
rect 207750 474308 207756 474320
rect 207808 474308 207814 474360
rect 245654 474308 245660 474360
rect 245712 474348 245718 474360
rect 366542 474348 366548 474360
rect 245712 474320 366548 474348
rect 245712 474308 245718 474320
rect 366542 474308 366548 474320
rect 366600 474308 366606 474360
rect 50246 474240 50252 474292
rect 50304 474280 50310 474292
rect 98638 474280 98644 474292
rect 50304 474252 98644 474280
rect 50304 474240 50310 474252
rect 98638 474240 98644 474252
rect 98696 474240 98702 474292
rect 179506 474240 179512 474292
rect 179564 474280 179570 474292
rect 214926 474280 214932 474292
rect 179564 474252 214932 474280
rect 179564 474240 179570 474252
rect 214926 474240 214932 474252
rect 214984 474240 214990 474292
rect 252738 474240 252744 474292
rect 252796 474280 252802 474292
rect 374822 474280 374828 474292
rect 252796 474252 374828 474280
rect 252796 474240 252802 474252
rect 374822 474240 374828 474252
rect 374880 474240 374886 474292
rect 51718 474172 51724 474224
rect 51776 474212 51782 474224
rect 99466 474212 99472 474224
rect 51776 474184 99472 474212
rect 51776 474172 51782 474184
rect 99466 474172 99472 474184
rect 99524 474172 99530 474224
rect 158898 474172 158904 474224
rect 158956 474212 158962 474224
rect 202230 474212 202236 474224
rect 158956 474184 202236 474212
rect 158956 474172 158962 474184
rect 202230 474172 202236 474184
rect 202288 474172 202294 474224
rect 243446 474172 243452 474224
rect 243504 474212 243510 474224
rect 366450 474212 366456 474224
rect 243504 474184 366456 474212
rect 243504 474172 243510 474184
rect 366450 474172 366456 474184
rect 366508 474172 366514 474224
rect 57790 474104 57796 474156
rect 57848 474144 57854 474156
rect 113266 474144 113272 474156
rect 57848 474116 113272 474144
rect 57848 474104 57854 474116
rect 113266 474104 113272 474116
rect 113324 474104 113330 474156
rect 168466 474104 168472 474156
rect 168524 474144 168530 474156
rect 214558 474144 214564 474156
rect 168524 474116 214564 474144
rect 168524 474104 168530 474116
rect 214558 474104 214564 474116
rect 214616 474104 214622 474156
rect 254026 474104 254032 474156
rect 254084 474144 254090 474156
rect 379054 474144 379060 474156
rect 254084 474116 379060 474144
rect 254084 474104 254090 474116
rect 379054 474104 379060 474116
rect 379112 474104 379118 474156
rect 45186 474036 45192 474088
rect 45244 474076 45250 474088
rect 104986 474076 104992 474088
rect 45244 474048 104992 474076
rect 45244 474036 45250 474048
rect 104986 474036 104992 474048
rect 105044 474036 105050 474088
rect 139486 474036 139492 474088
rect 139544 474076 139550 474088
rect 207290 474076 207296 474088
rect 139544 474048 207296 474076
rect 139544 474036 139550 474048
rect 207290 474036 207296 474048
rect 207348 474036 207354 474088
rect 231854 474036 231860 474088
rect 231912 474076 231918 474088
rect 363690 474076 363696 474088
rect 231912 474048 363696 474076
rect 231912 474036 231918 474048
rect 363690 474036 363696 474048
rect 363748 474036 363754 474088
rect 59354 473968 59360 474020
rect 59412 474008 59418 474020
rect 180150 474008 180156 474020
rect 59412 473980 180156 474008
rect 59412 473968 59418 473980
rect 180150 473968 180156 473980
rect 180208 473968 180214 474020
rect 185578 473968 185584 474020
rect 185636 474008 185642 474020
rect 205818 474008 205824 474020
rect 185636 473980 205824 474008
rect 185636 473968 185642 473980
rect 205818 473968 205824 473980
rect 205876 473968 205882 474020
rect 227806 473968 227812 474020
rect 227864 474008 227870 474020
rect 362310 474008 362316 474020
rect 227864 473980 362316 474008
rect 227864 473968 227870 473980
rect 362310 473968 362316 473980
rect 362368 473968 362374 474020
rect 288526 473900 288532 473952
rect 288584 473940 288590 473952
rect 369026 473940 369032 473952
rect 288584 473912 369032 473940
rect 288584 473900 288590 473912
rect 369026 473900 369032 473912
rect 369084 473900 369090 473952
rect 289906 473832 289912 473884
rect 289964 473872 289970 473884
rect 365530 473872 365536 473884
rect 289964 473844 365536 473872
rect 289964 473832 289970 473844
rect 365530 473832 365536 473844
rect 365588 473832 365594 473884
rect 299014 473220 299020 473272
rect 299072 473260 299078 473272
rect 367646 473260 367652 473272
rect 299072 473232 367652 473260
rect 299072 473220 299078 473232
rect 367646 473220 367652 473232
rect 367704 473220 367710 473272
rect 285950 473152 285956 473204
rect 286008 473192 286014 473204
rect 361482 473192 361488 473204
rect 286008 473164 361488 473192
rect 286008 473152 286014 473164
rect 361482 473152 361488 473164
rect 361540 473152 361546 473204
rect 262858 473084 262864 473136
rect 262916 473124 262922 473136
rect 370958 473124 370964 473136
rect 262916 473096 370964 473124
rect 262916 473084 262922 473096
rect 370958 473084 370964 473096
rect 371016 473084 371022 473136
rect 240134 473016 240140 473068
rect 240192 473056 240198 473068
rect 362494 473056 362500 473068
rect 240192 473028 362500 473056
rect 240192 473016 240198 473028
rect 362494 473016 362500 473028
rect 362552 473016 362558 473068
rect 241606 472948 241612 473000
rect 241664 472988 241670 473000
rect 374638 472988 374644 473000
rect 241664 472960 374644 472988
rect 241664 472948 241670 472960
rect 374638 472948 374644 472960
rect 374696 472948 374702 473000
rect 240226 472880 240232 472932
rect 240284 472920 240290 472932
rect 373350 472920 373356 472932
rect 240284 472892 373356 472920
rect 240284 472880 240290 472892
rect 373350 472880 373356 472892
rect 373408 472880 373414 472932
rect 58710 472812 58716 472864
rect 58768 472852 58774 472864
rect 110598 472852 110604 472864
rect 58768 472824 110604 472852
rect 58768 472812 58774 472824
rect 110598 472812 110604 472824
rect 110656 472812 110662 472864
rect 226426 472812 226432 472864
rect 226484 472852 226490 472864
rect 367738 472852 367744 472864
rect 226484 472824 367744 472852
rect 226484 472812 226490 472824
rect 367738 472812 367744 472824
rect 367796 472812 367802 472864
rect 45002 472744 45008 472796
rect 45060 472784 45066 472796
rect 105630 472784 105636 472796
rect 45060 472756 105636 472784
rect 45060 472744 45066 472756
rect 105630 472744 105636 472756
rect 105688 472744 105694 472796
rect 175366 472744 175372 472796
rect 175424 472784 175430 472796
rect 202414 472784 202420 472796
rect 175424 472756 202420 472784
rect 175424 472744 175430 472756
rect 202414 472744 202420 472756
rect 202472 472744 202478 472796
rect 237374 472744 237380 472796
rect 237432 472784 237438 472796
rect 378962 472784 378968 472796
rect 237432 472756 378968 472784
rect 237432 472744 237438 472756
rect 378962 472744 378968 472756
rect 379020 472744 379026 472796
rect 45278 472676 45284 472728
rect 45336 472716 45342 472728
rect 106366 472716 106372 472728
rect 45336 472688 106372 472716
rect 45336 472676 45342 472688
rect 106366 472676 106372 472688
rect 106424 472676 106430 472728
rect 169938 472676 169944 472728
rect 169996 472716 170002 472728
rect 214650 472716 214656 472728
rect 169996 472688 214656 472716
rect 169996 472676 170002 472688
rect 214650 472676 214656 472688
rect 214708 472676 214714 472728
rect 227714 472676 227720 472728
rect 227772 472716 227778 472728
rect 371878 472716 371884 472728
rect 227772 472688 371884 472716
rect 227772 472676 227778 472688
rect 371878 472676 371884 472688
rect 371936 472676 371942 472728
rect 45370 472608 45376 472660
rect 45428 472648 45434 472660
rect 106458 472648 106464 472660
rect 45428 472620 106464 472648
rect 45428 472608 45434 472620
rect 106458 472608 106464 472620
rect 106516 472608 106522 472660
rect 160370 472608 160376 472660
rect 160428 472648 160434 472660
rect 210510 472648 210516 472660
rect 160428 472620 210516 472648
rect 160428 472608 160434 472620
rect 210510 472608 210516 472620
rect 210568 472608 210574 472660
rect 226334 472608 226340 472660
rect 226392 472648 226398 472660
rect 370590 472648 370596 472660
rect 226392 472620 370596 472648
rect 226392 472608 226398 472620
rect 370590 472608 370596 472620
rect 370648 472608 370654 472660
rect 52270 471928 52276 471980
rect 52328 471968 52334 471980
rect 82814 471968 82820 471980
rect 52328 471940 82820 471968
rect 52328 471928 52334 471940
rect 82814 471928 82820 471940
rect 82872 471928 82878 471980
rect 182266 471928 182272 471980
rect 182324 471968 182330 471980
rect 205174 471968 205180 471980
rect 182324 471940 205180 471968
rect 182324 471928 182330 471940
rect 205174 471928 205180 471940
rect 205232 471928 205238 471980
rect 285766 471928 285772 471980
rect 285824 471968 285830 471980
rect 357158 471968 357164 471980
rect 285824 471940 357164 471968
rect 285824 471928 285830 471940
rect 357158 471928 357164 471940
rect 357216 471928 357222 471980
rect 42334 471860 42340 471912
rect 42392 471900 42398 471912
rect 74350 471900 74356 471912
rect 42392 471872 74356 471900
rect 42392 471860 42398 471872
rect 74350 471860 74356 471872
rect 74408 471860 74414 471912
rect 190638 471860 190644 471912
rect 190696 471900 190702 471912
rect 216214 471900 216220 471912
rect 190696 471872 216220 471900
rect 190696 471860 190702 471872
rect 216214 471860 216220 471872
rect 216272 471860 216278 471912
rect 287514 471860 287520 471912
rect 287572 471900 287578 471912
rect 359550 471900 359556 471912
rect 287572 471872 359556 471900
rect 287572 471860 287578 471872
rect 359550 471860 359556 471872
rect 359608 471860 359614 471912
rect 49602 471792 49608 471844
rect 49660 471832 49666 471844
rect 82262 471832 82268 471844
rect 49660 471804 82268 471832
rect 49660 471792 49666 471804
rect 82262 471792 82268 471804
rect 82320 471792 82326 471844
rect 174814 471792 174820 471844
rect 174872 471832 174878 471844
rect 200850 471832 200856 471844
rect 174872 471804 200856 471832
rect 174872 471792 174878 471804
rect 200850 471792 200856 471804
rect 200908 471792 200914 471844
rect 295518 471792 295524 471844
rect 295576 471832 295582 471844
rect 368934 471832 368940 471844
rect 295576 471804 368940 471832
rect 295576 471792 295582 471804
rect 368934 471792 368940 471804
rect 368992 471792 368998 471844
rect 52178 471724 52184 471776
rect 52236 471764 52242 471776
rect 84286 471764 84292 471776
rect 52236 471736 84292 471764
rect 52236 471724 52242 471736
rect 84286 471724 84292 471736
rect 84344 471724 84350 471776
rect 182358 471724 182364 471776
rect 182416 471764 182422 471776
rect 209314 471764 209320 471776
rect 182416 471736 209320 471764
rect 182416 471724 182422 471736
rect 209314 471724 209320 471736
rect 209372 471724 209378 471776
rect 295426 471724 295432 471776
rect 295484 471764 295490 471776
rect 370222 471764 370228 471776
rect 295484 471736 370228 471764
rect 295484 471724 295490 471736
rect 370222 471724 370228 471736
rect 370280 471724 370286 471776
rect 50062 471656 50068 471708
rect 50120 471696 50126 471708
rect 82906 471696 82912 471708
rect 50120 471668 82912 471696
rect 50120 471656 50126 471668
rect 82906 471656 82912 471668
rect 82964 471656 82970 471708
rect 183738 471656 183744 471708
rect 183796 471696 183802 471708
rect 210878 471696 210884 471708
rect 183796 471668 210884 471696
rect 183796 471656 183802 471668
rect 210878 471656 210884 471668
rect 210936 471656 210942 471708
rect 296254 471656 296260 471708
rect 296312 471696 296318 471708
rect 373074 471696 373080 471708
rect 296312 471668 373080 471696
rect 296312 471656 296318 471668
rect 373074 471656 373080 471668
rect 373132 471656 373138 471708
rect 52914 471588 52920 471640
rect 52972 471628 52978 471640
rect 85758 471628 85764 471640
rect 52972 471600 85764 471628
rect 52972 471588 52978 471600
rect 85758 471588 85764 471600
rect 85816 471588 85822 471640
rect 139394 471588 139400 471640
rect 139452 471628 139458 471640
rect 196894 471628 196900 471640
rect 139452 471600 196900 471628
rect 139452 471588 139458 471600
rect 196894 471588 196900 471600
rect 196952 471588 196958 471640
rect 295334 471588 295340 471640
rect 295392 471628 295398 471640
rect 376846 471628 376852 471640
rect 295392 471600 376852 471628
rect 295392 471588 295398 471600
rect 376846 471588 376852 471600
rect 376904 471588 376910 471640
rect 50798 471520 50804 471572
rect 50856 471560 50862 471572
rect 84930 471560 84936 471572
rect 50856 471532 84936 471560
rect 50856 471520 50862 471532
rect 84930 471520 84936 471532
rect 84988 471520 84994 471572
rect 140958 471520 140964 471572
rect 141016 471560 141022 471572
rect 200482 471560 200488 471572
rect 141016 471532 200488 471560
rect 141016 471520 141022 471532
rect 200482 471520 200488 471532
rect 200540 471520 200546 471572
rect 292666 471520 292672 471572
rect 292724 471560 292730 471572
rect 376570 471560 376576 471572
rect 292724 471532 376576 471560
rect 292724 471520 292730 471532
rect 376570 471520 376576 471532
rect 376628 471520 376634 471572
rect 49510 471452 49516 471504
rect 49568 471492 49574 471504
rect 83182 471492 83188 471504
rect 49568 471464 83188 471492
rect 49568 471452 49574 471464
rect 83182 471452 83188 471464
rect 83240 471452 83246 471504
rect 140866 471452 140872 471504
rect 140924 471492 140930 471504
rect 204438 471492 204444 471504
rect 140924 471464 204444 471492
rect 140924 471452 140930 471464
rect 204438 471452 204444 471464
rect 204496 471452 204502 471504
rect 294046 471452 294052 471504
rect 294104 471492 294110 471504
rect 379330 471492 379336 471504
rect 294104 471464 379336 471492
rect 294104 471452 294110 471464
rect 379330 471452 379336 471464
rect 379388 471452 379394 471504
rect 57698 471384 57704 471436
rect 57756 471424 57762 471436
rect 113358 471424 113364 471436
rect 57756 471396 113364 471424
rect 57756 471384 57762 471396
rect 113358 471384 113364 471396
rect 113416 471384 113422 471436
rect 142338 471384 142344 471436
rect 142396 471424 142402 471436
rect 207382 471424 207388 471436
rect 142396 471396 207388 471424
rect 142396 471384 142402 471396
rect 207382 471384 207388 471396
rect 207440 471384 207446 471436
rect 285858 471384 285864 471436
rect 285916 471424 285922 471436
rect 374454 471424 374460 471436
rect 285916 471396 374460 471424
rect 285916 471384 285922 471396
rect 374454 471384 374460 471396
rect 374512 471384 374518 471436
rect 54570 471316 54576 471368
rect 54628 471356 54634 471368
rect 102318 471356 102324 471368
rect 54628 471328 102324 471356
rect 54628 471316 54634 471328
rect 102318 471316 102324 471328
rect 102376 471316 102382 471368
rect 109218 471316 109224 471368
rect 109276 471356 109282 471368
rect 197630 471356 197636 471368
rect 109276 471328 197636 471356
rect 109276 471316 109282 471328
rect 197630 471316 197636 471328
rect 197688 471316 197694 471368
rect 259546 471316 259552 471368
rect 259604 471356 259610 471368
rect 369394 471356 369400 471368
rect 259604 471328 369400 471356
rect 259604 471316 259610 471328
rect 369394 471316 369400 471328
rect 369452 471316 369458 471368
rect 53098 471248 53104 471300
rect 53156 471288 53162 471300
rect 101214 471288 101220 471300
rect 53156 471260 101220 471288
rect 53156 471248 53162 471260
rect 101214 471248 101220 471260
rect 101272 471248 101278 471300
rect 109126 471248 109132 471300
rect 109184 471288 109190 471300
rect 201678 471288 201684 471300
rect 109184 471260 201684 471288
rect 109184 471248 109190 471260
rect 201678 471248 201684 471260
rect 201736 471248 201742 471300
rect 250530 471248 250536 471300
rect 250588 471288 250594 471300
rect 365162 471288 365168 471300
rect 250588 471260 365168 471288
rect 250588 471248 250594 471260
rect 365162 471248 365168 471260
rect 365220 471248 365226 471300
rect 52086 471180 52092 471232
rect 52144 471220 52150 471232
rect 81526 471220 81532 471232
rect 52144 471192 81532 471220
rect 52144 471180 52150 471192
rect 81526 471180 81532 471192
rect 81584 471180 81590 471232
rect 192294 471180 192300 471232
rect 192352 471220 192358 471232
rect 213362 471220 213368 471232
rect 192352 471192 213368 471220
rect 192352 471180 192358 471192
rect 213362 471180 213368 471192
rect 213420 471180 213426 471232
rect 299474 471180 299480 471232
rect 299532 471220 299538 471232
rect 368842 471220 368848 471232
rect 299532 471192 368848 471220
rect 299532 471180 299538 471192
rect 368842 471180 368848 471192
rect 368900 471180 368906 471232
rect 46198 471112 46204 471164
rect 46256 471152 46262 471164
rect 64966 471152 64972 471164
rect 46256 471124 64972 471152
rect 46256 471112 46262 471124
rect 64966 471112 64972 471124
rect 65024 471112 65030 471164
rect 190546 471112 190552 471164
rect 190604 471152 190610 471164
rect 211522 471152 211528 471164
rect 190604 471124 211528 471152
rect 190604 471112 190610 471124
rect 211522 471112 211528 471124
rect 211580 471112 211586 471164
rect 47486 471044 47492 471096
rect 47544 471084 47550 471096
rect 64874 471084 64880 471096
rect 47544 471056 64880 471084
rect 47544 471044 47550 471056
rect 64874 471044 64880 471056
rect 64932 471044 64938 471096
rect 193858 470636 193864 470688
rect 193916 470676 193922 470688
rect 201862 470676 201868 470688
rect 193916 470648 201868 470676
rect 193916 470636 193922 470648
rect 201862 470636 201868 470648
rect 201920 470636 201926 470688
rect 289814 470500 289820 470552
rect 289872 470540 289878 470552
rect 366266 470540 366272 470552
rect 289872 470512 366272 470540
rect 289872 470500 289878 470512
rect 366266 470500 366272 470512
rect 366324 470500 366330 470552
rect 283098 470432 283104 470484
rect 283156 470472 283162 470484
rect 359918 470472 359924 470484
rect 283156 470444 359924 470472
rect 283156 470432 283162 470444
rect 359918 470432 359924 470444
rect 359976 470432 359982 470484
rect 282914 470364 282920 470416
rect 282972 470404 282978 470416
rect 360010 470404 360016 470416
rect 282972 470376 360016 470404
rect 282972 470364 282978 470376
rect 360010 470364 360016 470376
rect 360068 470364 360074 470416
rect 281534 470296 281540 470348
rect 281592 470336 281598 470348
rect 359734 470336 359740 470348
rect 281592 470308 359740 470336
rect 281592 470296 281598 470308
rect 359734 470296 359740 470308
rect 359792 470296 359798 470348
rect 296806 470228 296812 470280
rect 296864 470268 296870 470280
rect 375374 470268 375380 470280
rect 296864 470240 375380 470268
rect 296864 470228 296870 470240
rect 375374 470228 375380 470240
rect 375432 470228 375438 470280
rect 281718 470160 281724 470212
rect 281776 470200 281782 470212
rect 367002 470200 367008 470212
rect 281776 470172 367008 470200
rect 281776 470160 281782 470172
rect 367002 470160 367008 470172
rect 367060 470160 367066 470212
rect 267826 470092 267832 470144
rect 267884 470132 267890 470144
rect 357986 470132 357992 470144
rect 267884 470104 357992 470132
rect 267884 470092 267890 470104
rect 357986 470092 357992 470104
rect 358044 470092 358050 470144
rect 285674 470024 285680 470076
rect 285732 470064 285738 470076
rect 377582 470064 377588 470076
rect 285732 470036 377588 470064
rect 285732 470024 285738 470036
rect 377582 470024 377588 470036
rect 377640 470024 377646 470076
rect 178034 469956 178040 470008
rect 178092 469996 178098 470008
rect 210786 469996 210792 470008
rect 178092 469968 210792 469996
rect 178092 469956 178098 469968
rect 210786 469956 210792 469968
rect 210844 469956 210850 470008
rect 281626 469956 281632 470008
rect 281684 469996 281690 470008
rect 373718 469996 373724 470008
rect 281684 469968 373724 469996
rect 281684 469956 281690 469968
rect 373718 469956 373724 469968
rect 373776 469956 373782 470008
rect 179414 469888 179420 469940
rect 179472 469928 179478 469940
rect 219066 469928 219072 469940
rect 179472 469900 219072 469928
rect 179472 469888 179478 469900
rect 219066 469888 219072 469900
rect 219124 469888 219130 469940
rect 284294 469888 284300 469940
rect 284352 469928 284358 469940
rect 377490 469928 377496 469940
rect 284352 469900 377496 469928
rect 284352 469888 284358 469900
rect 377490 469888 377496 469900
rect 377548 469888 377554 469940
rect 57606 469820 57612 469872
rect 57664 469860 57670 469872
rect 111978 469860 111984 469872
rect 57664 469832 111984 469860
rect 57664 469820 57670 469832
rect 111978 469820 111984 469832
rect 112036 469820 112042 469872
rect 116578 469820 116584 469872
rect 116636 469860 116642 469872
rect 199470 469860 199476 469872
rect 116636 469832 199476 469860
rect 116636 469820 116642 469832
rect 199470 469820 199476 469832
rect 199528 469820 199534 469872
rect 265250 469820 265256 469872
rect 265308 469860 265314 469872
rect 361114 469860 361120 469872
rect 265308 469832 361120 469860
rect 265308 469820 265314 469832
rect 361114 469820 361120 469832
rect 361172 469820 361178 469872
rect 283006 469752 283012 469804
rect 283064 469792 283070 469804
rect 357802 469792 357808 469804
rect 283064 469764 357808 469792
rect 283064 469752 283070 469764
rect 357802 469752 357808 469764
rect 357860 469752 357866 469804
rect 48222 469140 48228 469192
rect 48280 469180 48286 469192
rect 80238 469180 80244 469192
rect 48280 469152 80244 469180
rect 48280 469140 48286 469152
rect 80238 469140 80244 469152
rect 80296 469140 80302 469192
rect 193398 469140 193404 469192
rect 193456 469180 193462 469192
rect 215846 469180 215852 469192
rect 193456 469152 215852 469180
rect 193456 469140 193462 469152
rect 215846 469140 215852 469152
rect 215904 469140 215910 469192
rect 277486 469140 277492 469192
rect 277544 469180 277550 469192
rect 365622 469180 365628 469192
rect 277544 469152 365628 469180
rect 277544 469140 277550 469152
rect 365622 469140 365628 469152
rect 365680 469140 365686 469192
rect 50706 469072 50712 469124
rect 50764 469112 50770 469124
rect 78674 469112 78680 469124
rect 50764 469084 78680 469112
rect 50764 469072 50770 469084
rect 78674 469072 78680 469084
rect 78732 469072 78738 469124
rect 191926 469072 191932 469124
rect 191984 469112 191990 469124
rect 217778 469112 217784 469124
rect 191984 469084 217784 469112
rect 191984 469072 191990 469084
rect 217778 469072 217784 469084
rect 217836 469072 217842 469124
rect 269114 469072 269120 469124
rect 269172 469112 269178 469124
rect 358538 469112 358544 469124
rect 269172 469084 358544 469112
rect 269172 469072 269178 469084
rect 358538 469072 358544 469084
rect 358596 469072 358602 469124
rect 46014 469004 46020 469056
rect 46072 469044 46078 469056
rect 63586 469044 63592 469056
rect 46072 469016 63592 469044
rect 46072 469004 46078 469016
rect 63586 469004 63592 469016
rect 63644 469004 63650 469056
rect 189166 469004 189172 469056
rect 189224 469044 189230 469056
rect 215110 469044 215116 469056
rect 189224 469016 215116 469044
rect 189224 469004 189230 469016
rect 215110 469004 215116 469016
rect 215168 469004 215174 469056
rect 273438 469004 273444 469056
rect 273496 469044 273502 469056
rect 364886 469044 364892 469056
rect 273496 469016 364892 469044
rect 273496 469004 273502 469016
rect 364886 469004 364892 469016
rect 364944 469004 364950 469056
rect 54846 468936 54852 468988
rect 54904 468976 54910 468988
rect 85666 468976 85672 468988
rect 54904 468948 85672 468976
rect 54904 468936 54910 468948
rect 85666 468936 85672 468948
rect 85724 468936 85730 468988
rect 180978 468936 180984 468988
rect 181036 468976 181042 468988
rect 210326 468976 210332 468988
rect 181036 468948 210332 468976
rect 181036 468936 181042 468948
rect 210326 468936 210332 468948
rect 210384 468936 210390 468988
rect 266354 468936 266360 468988
rect 266412 468976 266418 468988
rect 359642 468976 359648 468988
rect 266412 468948 359648 468976
rect 266412 468936 266418 468948
rect 359642 468936 359648 468948
rect 359700 468936 359706 468988
rect 56042 468868 56048 468920
rect 56100 468908 56106 468920
rect 86954 468908 86960 468920
rect 56100 468880 86960 468908
rect 56100 468868 56106 468880
rect 86954 468868 86960 468880
rect 87012 468868 87018 468920
rect 175274 468868 175280 468920
rect 175332 468908 175338 468920
rect 212166 468908 212172 468920
rect 175332 468880 212172 468908
rect 175332 468868 175338 468880
rect 212166 468868 212172 468880
rect 212224 468868 212230 468920
rect 266446 468868 266452 468920
rect 266504 468908 266510 468920
rect 361206 468908 361212 468920
rect 266504 468880 361212 468908
rect 266504 468868 266510 468880
rect 361206 468868 361212 468880
rect 361264 468868 361270 468920
rect 54938 468800 54944 468852
rect 54996 468840 55002 468852
rect 87046 468840 87052 468852
rect 54996 468812 87052 468840
rect 54996 468800 55002 468812
rect 87046 468800 87052 468812
rect 87104 468800 87110 468852
rect 158806 468800 158812 468852
rect 158864 468840 158870 468852
rect 207658 468840 207664 468852
rect 158864 468812 207664 468840
rect 158864 468800 158870 468812
rect 207658 468800 207664 468812
rect 207716 468800 207722 468852
rect 255314 468800 255320 468852
rect 255372 468840 255378 468852
rect 358446 468840 358452 468852
rect 255372 468812 358452 468840
rect 255372 468800 255378 468812
rect 358446 468800 358452 468812
rect 358504 468800 358510 468852
rect 53190 468732 53196 468784
rect 53248 468772 53254 468784
rect 85574 468772 85580 468784
rect 53248 468744 85580 468772
rect 53248 468732 53254 468744
rect 85574 468732 85580 468744
rect 85632 468732 85638 468784
rect 161474 468732 161480 468784
rect 161532 468772 161538 468784
rect 215938 468772 215944 468784
rect 161532 468744 215944 468772
rect 161532 468732 161538 468744
rect 215938 468732 215944 468744
rect 215996 468732 216002 468784
rect 265158 468732 265164 468784
rect 265216 468772 265222 468784
rect 371602 468772 371608 468784
rect 265216 468744 371608 468772
rect 265216 468732 265222 468744
rect 371602 468732 371608 468744
rect 371660 468732 371666 468784
rect 59906 468664 59912 468716
rect 59964 468704 59970 468716
rect 92658 468704 92664 468716
rect 59964 468676 92664 468704
rect 59964 468664 59970 468676
rect 92658 468664 92664 468676
rect 92716 468664 92722 468716
rect 109034 468664 109040 468716
rect 109092 468704 109098 468716
rect 197722 468704 197728 468716
rect 109092 468676 197728 468704
rect 109092 468664 109098 468676
rect 197722 468664 197728 468676
rect 197780 468664 197786 468716
rect 266538 468664 266544 468716
rect 266596 468704 266602 468716
rect 375006 468704 375012 468716
rect 266596 468676 375012 468704
rect 266596 468664 266602 468676
rect 375006 468664 375012 468676
rect 375064 468664 375070 468716
rect 50614 468596 50620 468648
rect 50672 468636 50678 468648
rect 92566 468636 92572 468648
rect 50672 468608 92572 468636
rect 50672 468596 50678 468608
rect 92566 468596 92572 468608
rect 92624 468596 92630 468648
rect 107746 468596 107752 468648
rect 107804 468636 107810 468648
rect 199102 468636 199108 468648
rect 107804 468608 199108 468636
rect 107804 468596 107810 468608
rect 199102 468596 199108 468608
rect 199160 468596 199166 468648
rect 249794 468596 249800 468648
rect 249852 468636 249858 468648
rect 367922 468636 367928 468648
rect 249852 468608 367928 468636
rect 249852 468596 249858 468608
rect 367922 468596 367928 468608
rect 367980 468596 367986 468648
rect 49418 468528 49424 468580
rect 49476 468568 49482 468580
rect 93946 468568 93952 468580
rect 49476 468540 93952 468568
rect 49476 468528 49482 468540
rect 93946 468528 93952 468540
rect 94004 468528 94010 468580
rect 107838 468528 107844 468580
rect 107896 468568 107902 468580
rect 200298 468568 200304 468580
rect 107896 468540 200304 468568
rect 107896 468528 107902 468540
rect 200298 468528 200304 468540
rect 200356 468528 200362 468580
rect 249886 468528 249892 468580
rect 249944 468568 249950 468580
rect 372062 468568 372068 468580
rect 249944 468540 372068 468568
rect 249944 468528 249950 468540
rect 372062 468528 372068 468540
rect 372120 468528 372126 468580
rect 44818 468460 44824 468512
rect 44876 468500 44882 468512
rect 103698 468500 103704 468512
rect 44876 468472 103704 468500
rect 44876 468460 44882 468472
rect 103698 468460 103704 468472
rect 103756 468460 103762 468512
rect 107654 468460 107660 468512
rect 107712 468500 107718 468512
rect 203058 468500 203064 468512
rect 107712 468472 203064 468500
rect 107712 468460 107718 468472
rect 203058 468460 203064 468472
rect 203116 468460 203122 468512
rect 252646 468460 252652 468512
rect 252704 468500 252710 468512
rect 374914 468500 374920 468512
rect 252704 468472 374920 468500
rect 252704 468460 252710 468472
rect 374914 468460 374920 468472
rect 374972 468460 374978 468512
rect 192018 468392 192024 468444
rect 192076 468432 192082 468444
rect 214374 468432 214380 468444
rect 192076 468404 214380 468432
rect 192076 468392 192082 468404
rect 214374 468392 214380 468404
rect 214432 468392 214438 468444
rect 293954 468392 293960 468444
rect 294012 468432 294018 468444
rect 377398 468432 377404 468444
rect 294012 468404 377404 468432
rect 294012 468392 294018 468404
rect 377398 468392 377404 468404
rect 377456 468392 377462 468444
rect 182174 468324 182180 468376
rect 182232 468364 182238 468376
rect 202506 468364 202512 468376
rect 182232 468336 202512 468364
rect 182232 468324 182238 468336
rect 202506 468324 202512 468336
rect 202564 468324 202570 468376
rect 296714 468324 296720 468376
rect 296772 468364 296778 468376
rect 378134 468364 378140 468376
rect 296772 468336 378140 468364
rect 296772 468324 296778 468336
rect 378134 468324 378140 468336
rect 378192 468324 378198 468376
rect 197262 468256 197268 468308
rect 197320 468296 197326 468308
rect 211246 468296 211252 468308
rect 197320 468268 211252 468296
rect 197320 468256 197326 468268
rect 211246 468256 211252 468268
rect 211304 468256 211310 468308
rect 52914 467916 52920 467968
rect 52972 467956 52978 467968
rect 53374 467956 53380 467968
rect 52972 467928 53380 467956
rect 52972 467916 52978 467928
rect 53374 467916 53380 467928
rect 53432 467916 53438 467968
rect 80698 467780 80704 467832
rect 80756 467820 80762 467832
rect 178034 467820 178040 467832
rect 80756 467792 178040 467820
rect 80756 467780 80762 467792
rect 178034 467780 178040 467792
rect 178092 467780 178098 467832
rect 291194 467712 291200 467764
rect 291252 467752 291258 467764
rect 358722 467752 358728 467764
rect 291252 467724 358728 467752
rect 291252 467712 291258 467724
rect 358722 467712 358728 467724
rect 358780 467712 358786 467764
rect 277394 467644 277400 467696
rect 277452 467684 277458 467696
rect 362862 467684 362868 467696
rect 277452 467656 362868 467684
rect 277452 467644 277458 467656
rect 362862 467644 362868 467656
rect 362920 467644 362926 467696
rect 42702 467576 42708 467628
rect 42760 467616 42766 467628
rect 66346 467616 66352 467628
rect 42760 467588 66352 467616
rect 42760 467576 42766 467588
rect 66346 467576 66352 467588
rect 66404 467576 66410 467628
rect 273254 467576 273260 467628
rect 273312 467616 273318 467628
rect 362126 467616 362132 467628
rect 273312 467588 362132 467616
rect 273312 467576 273318 467588
rect 362126 467576 362132 467588
rect 362184 467576 362190 467628
rect 41322 467508 41328 467560
rect 41380 467548 41386 467560
rect 70486 467548 70492 467560
rect 41380 467520 70492 467548
rect 41380 467508 41386 467520
rect 70486 467508 70492 467520
rect 70544 467508 70550 467560
rect 273346 467508 273352 467560
rect 273404 467548 273410 467560
rect 369670 467548 369676 467560
rect 273404 467520 369676 467548
rect 273404 467508 273410 467520
rect 369670 467508 369676 467520
rect 369728 467508 369734 467560
rect 41230 467440 41236 467492
rect 41288 467480 41294 467492
rect 71866 467480 71872 467492
rect 41288 467452 71872 467480
rect 41288 467440 41294 467452
rect 71866 467440 71872 467452
rect 71924 467440 71930 467492
rect 189074 467440 189080 467492
rect 189132 467480 189138 467492
rect 202138 467480 202144 467492
rect 189132 467452 202144 467480
rect 189132 467440 189138 467452
rect 202138 467440 202144 467452
rect 202196 467440 202202 467492
rect 253934 467440 253940 467492
rect 253992 467480 253998 467492
rect 362678 467480 362684 467492
rect 253992 467452 362684 467480
rect 253992 467440 253998 467452
rect 362678 467440 362684 467452
rect 362736 467440 362742 467492
rect 42242 467372 42248 467424
rect 42300 467412 42306 467424
rect 73798 467412 73804 467424
rect 42300 467384 73804 467412
rect 42300 467372 42306 467384
rect 73798 467372 73804 467384
rect 73856 467372 73862 467424
rect 184934 467372 184940 467424
rect 184992 467412 184998 467424
rect 213178 467412 213184 467424
rect 184992 467384 213184 467412
rect 184992 467372 184998 467384
rect 213178 467372 213184 467384
rect 213236 467372 213242 467424
rect 262306 467372 262312 467424
rect 262364 467412 262370 467424
rect 372246 467412 372252 467424
rect 262364 467384 372252 467412
rect 262364 467372 262370 467384
rect 372246 467372 372252 467384
rect 372304 467372 372310 467424
rect 41138 467304 41144 467356
rect 41196 467344 41202 467356
rect 73890 467344 73896 467356
rect 41196 467316 73896 467344
rect 41196 467304 41202 467316
rect 73890 467304 73896 467316
rect 73948 467304 73954 467356
rect 172514 467304 172520 467356
rect 172572 467344 172578 467356
rect 204990 467344 204996 467356
rect 172572 467316 204996 467344
rect 172572 467304 172578 467316
rect 204990 467304 204996 467316
rect 205048 467304 205054 467356
rect 258074 467304 258080 467356
rect 258132 467344 258138 467356
rect 368014 467344 368020 467356
rect 258132 467316 368020 467344
rect 258132 467304 258138 467316
rect 368014 467304 368020 467316
rect 368072 467304 368078 467356
rect 41046 467236 41052 467288
rect 41104 467276 41110 467288
rect 93854 467276 93860 467288
rect 41104 467248 93860 467276
rect 41104 467236 41110 467248
rect 93854 467236 93860 467248
rect 93912 467236 93918 467288
rect 180150 467236 180156 467288
rect 180208 467276 180214 467288
rect 218238 467276 218244 467288
rect 180208 467248 218244 467276
rect 180208 467236 180214 467248
rect 218238 467236 218244 467248
rect 218296 467236 218302 467288
rect 251174 467236 251180 467288
rect 251232 467276 251238 467288
rect 363874 467276 363880 467288
rect 251232 467248 363880 467276
rect 251232 467236 251238 467248
rect 363874 467236 363880 467248
rect 363932 467236 363938 467288
rect 57514 467168 57520 467220
rect 57572 467208 57578 467220
rect 114738 467208 114744 467220
rect 57572 467180 114744 467208
rect 57572 467168 57578 467180
rect 114738 467168 114744 467180
rect 114796 467168 114802 467220
rect 149054 467168 149060 467220
rect 149112 467208 149118 467220
rect 212902 467208 212908 467220
rect 149112 467180 212908 467208
rect 149112 467168 149118 467180
rect 212902 467168 212908 467180
rect 212960 467168 212966 467220
rect 251266 467168 251272 467220
rect 251324 467208 251330 467220
rect 368198 467208 368204 467220
rect 251324 467180 368204 467208
rect 251324 467168 251330 467180
rect 368198 467168 368204 467180
rect 368256 467168 368262 467220
rect 44910 467100 44916 467152
rect 44968 467140 44974 467152
rect 106274 467140 106280 467152
rect 44968 467112 106280 467140
rect 44968 467100 44974 467112
rect 106274 467100 106280 467112
rect 106332 467100 106338 467152
rect 146294 467100 146300 467152
rect 146352 467140 146358 467152
rect 218698 467140 218704 467152
rect 146352 467112 218704 467140
rect 146352 467100 146358 467112
rect 218698 467100 218704 467112
rect 218756 467100 218762 467152
rect 252554 467100 252560 467152
rect 252612 467140 252618 467152
rect 379146 467140 379152 467152
rect 252612 467112 379152 467140
rect 252612 467100 252618 467112
rect 379146 467100 379152 467112
rect 379204 467100 379210 467152
rect 178034 466556 178040 466608
rect 178092 466596 178098 466608
rect 208578 466596 208584 466608
rect 178092 466568 208584 466596
rect 178092 466556 178098 466568
rect 208578 466556 208584 466568
rect 208636 466596 208642 466608
rect 208636 466568 209774 466596
rect 208636 466556 208642 466568
rect 47394 466488 47400 466540
rect 47452 466528 47458 466540
rect 47452 466500 207520 466528
rect 47452 466488 47458 466500
rect 207492 466472 207520 466500
rect 190914 466420 190920 466472
rect 190972 466460 190978 466472
rect 207014 466460 207020 466472
rect 190972 466432 207020 466460
rect 190972 466420 190978 466432
rect 207014 466420 207020 466432
rect 207072 466420 207078 466472
rect 207474 466420 207480 466472
rect 207532 466460 207538 466472
rect 207934 466460 207940 466472
rect 207532 466432 207940 466460
rect 207532 466420 207538 466432
rect 207934 466420 207940 466432
rect 207992 466420 207998 466472
rect 209746 466460 209774 466568
rect 339402 466556 339408 466608
rect 339460 466596 339466 466608
rect 362954 466596 362960 466608
rect 339460 466568 362960 466596
rect 339460 466556 339466 466568
rect 362954 466556 362960 466568
rect 363012 466556 363018 466608
rect 498194 466556 498200 466608
rect 498252 466596 498258 466608
rect 517790 466596 517796 466608
rect 498252 466568 517796 466596
rect 498252 466556 498258 466568
rect 517790 466556 517796 466568
rect 517848 466556 517854 466608
rect 218238 466488 218244 466540
rect 218296 466528 218302 466540
rect 339770 466528 339776 466540
rect 218296 466500 339776 466528
rect 218296 466488 218302 466500
rect 339770 466488 339776 466500
rect 339828 466528 339834 466540
rect 356974 466528 356980 466540
rect 339828 466500 356980 466528
rect 339828 466488 339834 466500
rect 356974 466488 356980 466500
rect 357032 466528 357038 466540
rect 499758 466528 499764 466540
rect 357032 466500 499764 466528
rect 357032 466488 357038 466500
rect 499758 466488 499764 466500
rect 499816 466528 499822 466540
rect 499816 466500 509234 466528
rect 499816 466488 499822 466500
rect 338482 466460 338488 466472
rect 209746 466432 338488 466460
rect 338482 466420 338488 466432
rect 338540 466460 338546 466472
rect 339402 466460 339408 466472
rect 338540 466432 339408 466460
rect 338540 466420 338546 466432
rect 339402 466420 339408 466432
rect 339460 466420 339466 466472
rect 350994 466420 351000 466472
rect 351052 466460 351058 466472
rect 360194 466460 360200 466472
rect 351052 466432 360200 466460
rect 351052 466420 351058 466432
rect 360194 466420 360200 466432
rect 360252 466420 360258 466472
rect 362954 466420 362960 466472
rect 363012 466460 363018 466472
rect 498194 466460 498200 466472
rect 363012 466432 498200 466460
rect 363012 466420 363018 466432
rect 498194 466420 498200 466432
rect 498252 466420 498258 466472
rect 509206 466460 509234 466500
rect 510890 466488 510896 466540
rect 510948 466528 510954 466540
rect 517514 466528 517520 466540
rect 510948 466500 517520 466528
rect 510948 466488 510954 466500
rect 517514 466488 517520 466500
rect 517572 466488 517578 466540
rect 517882 466460 517888 466472
rect 509206 466432 517888 466460
rect 517882 466420 517888 466432
rect 517940 466420 517946 466472
rect 53650 466352 53656 466404
rect 53708 466392 53714 466404
rect 77294 466392 77300 466404
rect 53708 466364 77300 466392
rect 53708 466352 53714 466364
rect 77294 466352 77300 466364
rect 77352 466352 77358 466404
rect 187786 466352 187792 466404
rect 187844 466392 187850 466404
rect 206646 466392 206652 466404
rect 187844 466364 206652 466392
rect 187844 466352 187850 466364
rect 206646 466352 206652 466364
rect 206704 466352 206710 466404
rect 274634 466352 274640 466404
rect 274692 466392 274698 466404
rect 366174 466392 366180 466404
rect 274692 466364 366180 466392
rect 274692 466352 274698 466364
rect 366174 466352 366180 466364
rect 366232 466352 366238 466404
rect 52362 466284 52368 466336
rect 52420 466324 52426 466336
rect 75914 466324 75920 466336
rect 52420 466296 75920 466324
rect 52420 466284 52426 466296
rect 75914 466284 75920 466296
rect 75972 466284 75978 466336
rect 183554 466284 183560 466336
rect 183612 466324 183618 466336
rect 207842 466324 207848 466336
rect 183612 466296 207848 466324
rect 183612 466284 183618 466296
rect 207842 466284 207848 466296
rect 207900 466284 207906 466336
rect 267734 466284 267740 466336
rect 267792 466324 267798 466336
rect 371786 466324 371792 466336
rect 267792 466296 371792 466324
rect 267792 466284 267798 466296
rect 371786 466284 371792 466296
rect 371844 466284 371850 466336
rect 59262 466216 59268 466268
rect 59320 466256 59326 466268
rect 67634 466256 67640 466268
rect 59320 466228 67640 466256
rect 59320 466216 59326 466228
rect 67634 466216 67640 466228
rect 67692 466216 67698 466268
rect 193214 466216 193220 466268
rect 193272 466256 193278 466268
rect 217594 466256 217600 466268
rect 193272 466228 217600 466256
rect 193272 466216 193278 466228
rect 217594 466216 217600 466228
rect 217652 466216 217658 466268
rect 259454 466216 259460 466268
rect 259512 466256 259518 466268
rect 369486 466256 369492 466268
rect 259512 466228 369492 466256
rect 259512 466216 259518 466228
rect 369486 466216 369492 466228
rect 369544 466216 369550 466268
rect 54478 466148 54484 466200
rect 54536 466188 54542 466200
rect 63494 466188 63500 466200
rect 54536 466160 63500 466188
rect 54536 466148 54542 466160
rect 63494 466148 63500 466160
rect 63552 466148 63558 466200
rect 180886 466148 180892 466200
rect 180944 466188 180950 466200
rect 205266 466188 205272 466200
rect 180944 466160 205272 466188
rect 180944 466148 180950 466160
rect 205266 466148 205272 466160
rect 205324 466148 205330 466200
rect 262214 466148 262220 466200
rect 262272 466188 262278 466200
rect 376386 466188 376392 466200
rect 262272 466160 376392 466188
rect 262272 466148 262278 466160
rect 376386 466148 376392 466160
rect 376444 466148 376450 466200
rect 51534 466080 51540 466132
rect 51592 466120 51598 466132
rect 66254 466120 66260 466132
rect 51592 466092 66260 466120
rect 51592 466080 51598 466092
rect 66254 466080 66260 466092
rect 66312 466080 66318 466132
rect 173894 466080 173900 466132
rect 173952 466120 173958 466132
rect 203794 466120 203800 466132
rect 173952 466092 203800 466120
rect 173952 466080 173958 466092
rect 203794 466080 203800 466092
rect 203852 466080 203858 466132
rect 248598 466080 248604 466132
rect 248656 466120 248662 466132
rect 369302 466120 369308 466132
rect 248656 466092 369308 466120
rect 248656 466080 248662 466092
rect 369302 466080 369308 466092
rect 369360 466080 369366 466132
rect 43438 466012 43444 466064
rect 43496 466052 43502 466064
rect 60734 466052 60740 466064
rect 43496 466024 60740 466052
rect 43496 466012 43502 466024
rect 60734 466012 60740 466024
rect 60792 466012 60798 466064
rect 173986 466012 173992 466064
rect 174044 466052 174050 466064
rect 216122 466052 216128 466064
rect 174044 466024 216128 466052
rect 174044 466012 174050 466024
rect 216122 466012 216128 466024
rect 216180 466012 216186 466064
rect 248506 466012 248512 466064
rect 248564 466052 248570 466064
rect 370774 466052 370780 466064
rect 248564 466024 370780 466052
rect 248564 466012 248570 466024
rect 370774 466012 370780 466024
rect 370832 466012 370838 466064
rect 44726 465944 44732 465996
rect 44784 465984 44790 465996
rect 62114 465984 62120 465996
rect 44784 465956 62120 465984
rect 44784 465944 44790 465956
rect 62114 465944 62120 465956
rect 62172 465944 62178 465996
rect 142154 465944 142160 465996
rect 142212 465984 142218 465996
rect 197814 465984 197820 465996
rect 142212 465956 197820 465984
rect 142212 465944 142218 465956
rect 197814 465944 197820 465956
rect 197872 465944 197878 465996
rect 248414 465944 248420 465996
rect 248472 465984 248478 465996
rect 373442 465984 373448 465996
rect 248472 465956 373448 465984
rect 248472 465944 248478 465956
rect 373442 465944 373448 465956
rect 373500 465944 373506 465996
rect 43346 465876 43352 465928
rect 43404 465916 43410 465928
rect 60826 465916 60832 465928
rect 43404 465888 60832 465916
rect 43404 465876 43410 465888
rect 60826 465876 60832 465888
rect 60884 465876 60890 465928
rect 142246 465876 142252 465928
rect 142304 465916 142310 465928
rect 200574 465916 200580 465928
rect 142304 465888 200580 465916
rect 142304 465876 142310 465888
rect 200574 465876 200580 465888
rect 200632 465876 200638 465928
rect 244274 465876 244280 465928
rect 244332 465916 244338 465928
rect 370682 465916 370688 465928
rect 244332 465888 370688 465916
rect 244332 465876 244338 465888
rect 370682 465876 370688 465888
rect 370740 465876 370746 465928
rect 53650 465808 53656 465860
rect 53708 465848 53714 465860
rect 74718 465848 74724 465860
rect 53708 465820 74724 465848
rect 53708 465808 53714 465820
rect 74718 465808 74724 465820
rect 74776 465808 74782 465860
rect 158714 465808 158720 465860
rect 158772 465848 158778 465860
rect 218882 465848 218888 465860
rect 158772 465820 218888 465848
rect 158772 465808 158778 465820
rect 218882 465808 218888 465820
rect 218940 465808 218946 465860
rect 241514 465808 241520 465860
rect 241572 465848 241578 465860
rect 369210 465848 369216 465860
rect 241572 465820 369216 465848
rect 241572 465808 241578 465820
rect 369210 465808 369216 465820
rect 369268 465808 369274 465860
rect 50062 465740 50068 465792
rect 50120 465780 50126 465792
rect 50706 465780 50712 465792
rect 50120 465752 50712 465780
rect 50120 465740 50126 465752
rect 50706 465740 50712 465752
rect 50764 465740 50770 465792
rect 51994 465740 52000 465792
rect 52052 465780 52058 465792
rect 52270 465780 52276 465792
rect 52052 465752 52276 465780
rect 52052 465740 52058 465752
rect 52270 465740 52276 465752
rect 52328 465740 52334 465792
rect 53006 465740 53012 465792
rect 53064 465780 53070 465792
rect 100846 465780 100852 465792
rect 53064 465752 100852 465780
rect 53064 465740 53070 465752
rect 100846 465740 100852 465752
rect 100904 465740 100910 465792
rect 140774 465740 140780 465792
rect 140832 465780 140838 465792
rect 205910 465780 205916 465792
rect 140832 465752 205916 465780
rect 140832 465740 140838 465752
rect 205910 465740 205916 465752
rect 205968 465740 205974 465792
rect 212442 465740 212448 465792
rect 212500 465780 212506 465792
rect 220906 465780 220912 465792
rect 212500 465752 220912 465780
rect 212500 465740 212506 465752
rect 220906 465740 220912 465752
rect 220964 465740 220970 465792
rect 235994 465740 236000 465792
rect 236052 465780 236058 465792
rect 365254 465780 365260 465792
rect 236052 465752 365260 465780
rect 236052 465740 236058 465752
rect 365254 465740 365260 465752
rect 365312 465740 365318 465792
rect 48222 465672 48228 465724
rect 48280 465712 48286 465724
rect 69014 465712 69020 465724
rect 48280 465684 69020 465712
rect 48280 465672 48286 465684
rect 69014 465672 69020 465684
rect 69072 465672 69078 465724
rect 72418 465672 72424 465724
rect 72476 465712 72482 465724
rect 198918 465712 198924 465724
rect 72476 465684 198924 465712
rect 72476 465672 72482 465684
rect 198918 465672 198924 465684
rect 198976 465672 198982 465724
rect 205450 465672 205456 465724
rect 205508 465712 205514 465724
rect 220998 465712 221004 465724
rect 205508 465684 221004 465712
rect 205508 465672 205514 465684
rect 220998 465672 221004 465684
rect 221056 465672 221062 465724
rect 242894 465672 242900 465724
rect 242952 465712 242958 465724
rect 374730 465712 374736 465724
rect 242952 465684 374736 465712
rect 242952 465672 242958 465684
rect 374730 465672 374736 465684
rect 374788 465672 374794 465724
rect 194594 465604 194600 465656
rect 194652 465644 194658 465656
rect 213086 465644 213092 465656
rect 194652 465616 213092 465644
rect 194652 465604 194658 465616
rect 213086 465604 213092 465616
rect 213144 465604 213150 465656
rect 288434 465604 288440 465656
rect 288492 465644 288498 465656
rect 357894 465644 357900 465656
rect 288492 465616 357900 465644
rect 288492 465604 288498 465616
rect 357894 465604 357900 465616
rect 357952 465604 357958 465656
rect 187694 465536 187700 465588
rect 187752 465576 187758 465588
rect 200942 465576 200948 465588
rect 187752 465548 200948 465576
rect 187752 465536 187758 465548
rect 200942 465536 200948 465548
rect 201000 465536 201006 465588
rect 298094 465536 298100 465588
rect 298152 465576 298158 465588
rect 360746 465576 360752 465588
rect 298152 465548 360752 465576
rect 298152 465536 298158 465548
rect 360746 465536 360752 465548
rect 360804 465536 360810 465588
rect 193306 465468 193312 465520
rect 193364 465508 193370 465520
rect 203978 465508 203984 465520
rect 193364 465480 203984 465508
rect 193364 465468 193370 465480
rect 203978 465468 203984 465480
rect 204036 465468 204042 465520
rect 198918 465060 198924 465112
rect 198976 465100 198982 465112
rect 358814 465100 358820 465112
rect 198976 465072 358820 465100
rect 198976 465060 198982 465072
rect 358814 465060 358820 465072
rect 358872 465100 358878 465112
rect 518894 465100 518900 465112
rect 358872 465072 518900 465100
rect 358872 465060 358878 465072
rect 518894 465060 518900 465072
rect 518952 465060 518958 465112
rect 196986 464992 196992 465044
rect 197044 465032 197050 465044
rect 200666 465032 200672 465044
rect 197044 465004 200672 465032
rect 197044 464992 197050 465004
rect 200666 464992 200672 465004
rect 200724 464992 200730 465044
rect 58986 464788 58992 464840
rect 59044 464828 59050 464840
rect 89898 464828 89904 464840
rect 59044 464800 89904 464828
rect 59044 464788 59050 464800
rect 89898 464788 89904 464800
rect 89956 464788 89962 464840
rect 191834 464788 191840 464840
rect 191892 464828 191898 464840
rect 210234 464828 210240 464840
rect 191892 464800 210240 464828
rect 191892 464788 191898 464800
rect 210234 464788 210240 464800
rect 210292 464788 210298 464840
rect 58894 464720 58900 464772
rect 58952 464760 58958 464772
rect 92474 464760 92480 464772
rect 58952 464732 92480 464760
rect 58952 464720 58958 464732
rect 92474 464720 92480 464732
rect 92532 464720 92538 464772
rect 190454 464720 190460 464772
rect 190512 464760 190518 464772
rect 208946 464760 208952 464772
rect 190512 464732 208952 464760
rect 190512 464720 190518 464732
rect 208946 464720 208952 464732
rect 209004 464720 209010 464772
rect 52914 464652 52920 464704
rect 52972 464692 52978 464704
rect 100754 464692 100760 464704
rect 52972 464664 100760 464692
rect 52972 464652 52978 464664
rect 100754 464652 100760 464664
rect 100812 464652 100818 464704
rect 127066 464652 127072 464704
rect 127124 464692 127130 464704
rect 197998 464692 198004 464704
rect 127124 464664 198004 464692
rect 127124 464652 127130 464664
rect 197998 464652 198004 464664
rect 198056 464652 198062 464704
rect 55858 464584 55864 464636
rect 55916 464624 55922 464636
rect 121454 464624 121460 464636
rect 55916 464596 121460 464624
rect 55916 464584 55922 464596
rect 121454 464584 121460 464596
rect 121512 464584 121518 464636
rect 126974 464584 126980 464636
rect 127032 464624 127038 464636
rect 199562 464624 199568 464636
rect 127032 464596 199568 464624
rect 127032 464584 127038 464596
rect 199562 464584 199568 464596
rect 199620 464584 199626 464636
rect 55766 464516 55772 464568
rect 55824 464556 55830 464568
rect 130010 464556 130016 464568
rect 55824 464528 130016 464556
rect 55824 464516 55830 464528
rect 130010 464516 130016 464528
rect 130068 464516 130074 464568
rect 180794 464516 180800 464568
rect 180852 464556 180858 464568
rect 206738 464556 206744 464568
rect 180852 464528 206744 464556
rect 180852 464516 180858 464528
rect 206738 464516 206744 464528
rect 206796 464516 206802 464568
rect 57146 464448 57152 464500
rect 57204 464488 57210 464500
rect 131298 464488 131304 464500
rect 57204 464460 131304 464488
rect 57204 464448 57210 464460
rect 131298 464448 131304 464460
rect 131356 464448 131362 464500
rect 186314 464448 186320 464500
rect 186372 464488 186378 464500
rect 212258 464488 212264 464500
rect 186372 464460 212264 464488
rect 186372 464448 186378 464460
rect 212258 464448 212264 464460
rect 212316 464448 212322 464500
rect 287054 464448 287060 464500
rect 287112 464488 287118 464500
rect 364794 464488 364800 464500
rect 287112 464460 364800 464488
rect 287112 464448 287118 464460
rect 364794 464448 364800 464460
rect 364852 464448 364858 464500
rect 54386 464380 54392 464432
rect 54444 464420 54450 464432
rect 133966 464420 133972 464432
rect 54444 464392 133972 464420
rect 54444 464380 54450 464392
rect 133966 464380 133972 464392
rect 134024 464380 134030 464432
rect 136634 464380 136640 464432
rect 136692 464420 136698 464432
rect 197906 464420 197912 464432
rect 136692 464392 197912 464420
rect 136692 464380 136698 464392
rect 197906 464380 197912 464392
rect 197964 464380 197970 464432
rect 271874 464380 271880 464432
rect 271932 464420 271938 464432
rect 373626 464420 373632 464432
rect 271932 464392 373632 464420
rect 271932 464380 271938 464392
rect 373626 464380 373632 464392
rect 373684 464380 373690 464432
rect 52270 464312 52276 464364
rect 52328 464352 52334 464364
rect 133874 464352 133880 464364
rect 52328 464324 133880 464352
rect 52328 464312 52334 464324
rect 133874 464312 133880 464324
rect 133932 464312 133938 464364
rect 136726 464312 136732 464364
rect 136784 464352 136790 464364
rect 199194 464352 199200 464364
rect 136784 464324 199200 464352
rect 136784 464312 136790 464324
rect 199194 464312 199200 464324
rect 199252 464312 199258 464364
rect 264974 464312 264980 464364
rect 265032 464352 265038 464364
rect 368106 464352 368112 464364
rect 265032 464324 368112 464352
rect 265032 464312 265038 464324
rect 368106 464312 368112 464324
rect 368164 464312 368170 464364
rect 207934 422900 207940 422952
rect 207992 422940 207998 422952
rect 217962 422940 217968 422952
rect 207992 422912 217968 422940
rect 207992 422900 207998 422912
rect 217962 422900 217968 422912
rect 218020 422900 218026 422952
rect 47394 418072 47400 418124
rect 47452 418112 47458 418124
rect 57882 418112 57888 418124
rect 47452 418084 57888 418112
rect 47452 418072 47458 418084
rect 57882 418072 57888 418084
rect 57940 418072 57946 418124
rect 207198 417392 207204 417444
rect 207256 417432 207262 417444
rect 216674 417432 216680 417444
rect 207256 417404 216680 417432
rect 207256 417392 207262 417404
rect 216674 417392 216680 417404
rect 216732 417392 216738 417444
rect 358078 417392 358084 417444
rect 358136 417432 358142 417444
rect 377214 417432 377220 417444
rect 358136 417404 377220 417432
rect 358136 417392 358142 417404
rect 377214 417392 377220 417404
rect 377272 417392 377278 417444
rect 44634 416780 44640 416832
rect 44692 416820 44698 416832
rect 57238 416820 57244 416832
rect 44692 416792 57244 416820
rect 44692 416780 44698 416792
rect 57238 416780 57244 416792
rect 57296 416780 57302 416832
rect 205726 416712 205732 416764
rect 205784 416752 205790 416764
rect 207198 416752 207204 416764
rect 205784 416724 207204 416752
rect 205784 416712 205790 416724
rect 207198 416712 207204 416724
rect 207256 416712 207262 416764
rect 208118 414808 208124 414860
rect 208176 414848 208182 414860
rect 216858 414848 216864 414860
rect 208176 414820 216864 414848
rect 208176 414808 208182 414820
rect 216858 414808 216864 414820
rect 216916 414808 216922 414860
rect 198090 414672 198096 414724
rect 198148 414712 198154 414724
rect 205634 414712 205640 414724
rect 198148 414684 205640 414712
rect 198148 414672 198154 414684
rect 205634 414672 205640 414684
rect 205692 414672 205698 414724
rect 207198 414672 207204 414724
rect 207256 414712 207262 414724
rect 217042 414712 217048 414724
rect 207256 414684 217048 414712
rect 207256 414672 207262 414684
rect 217042 414672 217048 414684
rect 217100 414672 217106 414724
rect 359826 414672 359832 414724
rect 359884 414712 359890 414724
rect 377674 414712 377680 414724
rect 359884 414684 377680 414712
rect 359884 414672 359890 414684
rect 377674 414672 377680 414684
rect 377732 414672 377738 414724
rect 48866 413992 48872 414044
rect 48924 414032 48930 414044
rect 57882 414032 57888 414044
rect 48924 414004 57888 414032
rect 48924 413992 48930 414004
rect 57882 413992 57888 414004
rect 57940 413992 57946 414044
rect 55674 413924 55680 413976
rect 55732 413964 55738 413976
rect 57054 413964 57060 413976
rect 55732 413936 57060 413964
rect 55732 413924 55738 413936
rect 57054 413924 57060 413936
rect 57112 413924 57118 413976
rect 204346 413924 204352 413976
rect 204404 413964 204410 413976
rect 206830 413964 206836 413976
rect 204404 413936 206836 413964
rect 204404 413924 204410 413936
rect 206830 413924 206836 413936
rect 206888 413924 206894 413976
rect 206002 413244 206008 413296
rect 206060 413284 206066 413296
rect 216858 413284 216864 413296
rect 206060 413256 216864 413284
rect 206060 413244 206066 413256
rect 216858 413244 216864 413256
rect 216916 413244 216922 413296
rect 48774 412768 48780 412820
rect 48832 412808 48838 412820
rect 57882 412808 57888 412820
rect 48832 412780 57888 412808
rect 48832 412768 48838 412780
rect 57882 412768 57888 412780
rect 57940 412768 57946 412820
rect 54294 412700 54300 412752
rect 54352 412740 54358 412752
rect 55858 412740 55864 412752
rect 54352 412712 55864 412740
rect 54352 412700 54358 412712
rect 55858 412700 55864 412712
rect 55916 412700 55922 412752
rect 357802 411884 357808 411936
rect 357860 411924 357866 411936
rect 377122 411924 377128 411936
rect 357860 411896 377128 411924
rect 357860 411884 357866 411896
rect 377122 411884 377128 411896
rect 377180 411884 377186 411936
rect 217778 411408 217784 411460
rect 217836 411448 217842 411460
rect 219250 411448 219256 411460
rect 217836 411420 219256 411448
rect 217836 411408 217842 411420
rect 219250 411408 219256 411420
rect 219308 411408 219314 411460
rect 47394 411272 47400 411324
rect 47452 411312 47458 411324
rect 57882 411312 57888 411324
rect 47452 411284 57888 411312
rect 47452 411272 47458 411284
rect 57882 411272 57888 411284
rect 57940 411272 57946 411324
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 14458 411244 14464 411256
rect 3016 411216 14464 411244
rect 3016 411204 3022 411216
rect 14458 411204 14464 411216
rect 14516 411204 14522 411256
rect 51626 410796 51632 410848
rect 51684 410836 51690 410848
rect 55858 410836 55864 410848
rect 51684 410808 55864 410836
rect 51684 410796 51690 410808
rect 55858 410796 55864 410808
rect 55916 410796 55922 410848
rect 206830 410524 206836 410576
rect 206888 410564 206894 410576
rect 216674 410564 216680 410576
rect 206888 410536 216680 410564
rect 206888 410524 206894 410536
rect 216674 410524 216680 410536
rect 216732 410564 216738 410576
rect 216950 410564 216956 410576
rect 216732 410536 216956 410564
rect 216732 410524 216738 410536
rect 216950 410524 216956 410536
rect 217008 410524 217014 410576
rect 360010 410524 360016 410576
rect 360068 410564 360074 410576
rect 377214 410564 377220 410576
rect 360068 410536 377220 410564
rect 360068 410524 360074 410536
rect 377214 410524 377220 410536
rect 377272 410524 377278 410576
rect 377398 410252 377404 410304
rect 377456 410292 377462 410304
rect 379238 410292 379244 410304
rect 377456 410264 379244 410292
rect 377456 410252 377462 410264
rect 379238 410252 379244 410264
rect 379296 410252 379302 410304
rect 51626 409844 51632 409896
rect 51684 409884 51690 409896
rect 56962 409884 56968 409896
rect 51684 409856 56968 409884
rect 51684 409844 51690 409856
rect 56962 409844 56968 409856
rect 57020 409844 57026 409896
rect 359918 409096 359924 409148
rect 359976 409136 359982 409148
rect 377398 409136 377404 409148
rect 359976 409108 377404 409136
rect 359976 409096 359982 409108
rect 377398 409096 377404 409108
rect 377456 409096 377462 409148
rect 52362 408484 52368 408536
rect 52420 408524 52426 408536
rect 57882 408524 57888 408536
rect 52420 408496 57888 408524
rect 52420 408484 52426 408496
rect 57882 408484 57888 408496
rect 57940 408484 57946 408536
rect 216674 407464 216680 407516
rect 216732 407504 216738 407516
rect 217042 407504 217048 407516
rect 216732 407476 217048 407504
rect 216732 407464 216738 407476
rect 217042 407464 217048 407476
rect 217100 407464 217106 407516
rect 216766 398216 216772 398268
rect 216824 398216 216830 398268
rect 216674 398012 216680 398064
rect 216732 398052 216738 398064
rect 216784 398052 216812 398216
rect 216732 398024 216812 398052
rect 216732 398012 216738 398024
rect 198090 397536 198096 397588
rect 198148 397576 198154 397588
rect 199010 397576 199016 397588
rect 198148 397548 199016 397576
rect 198148 397536 198154 397548
rect 199010 397536 199016 397548
rect 199068 397536 199074 397588
rect 198182 396788 198188 396840
rect 198240 396828 198246 396840
rect 199562 396828 199568 396840
rect 198240 396800 199568 396828
rect 198240 396788 198246 396800
rect 199562 396788 199568 396800
rect 199620 396788 199626 396840
rect 520918 396720 520924 396772
rect 520976 396760 520982 396772
rect 580350 396760 580356 396772
rect 520976 396732 580356 396760
rect 520976 396720 520982 396732
rect 580350 396720 580356 396732
rect 580408 396720 580414 396772
rect 216674 392028 216680 392080
rect 216732 392068 216738 392080
rect 217042 392068 217048 392080
rect 216732 392040 217048 392068
rect 216732 392028 216738 392040
rect 217042 392028 217048 392040
rect 217100 392028 217106 392080
rect 43254 391892 43260 391944
rect 43312 391932 43318 391944
rect 57882 391932 57888 391944
rect 43312 391904 57888 391932
rect 43312 391892 43318 391904
rect 57882 391892 57888 391904
rect 57940 391892 57946 391944
rect 209498 391892 209504 391944
rect 209556 391932 209562 391944
rect 216674 391932 216680 391944
rect 209556 391904 216680 391932
rect 209556 391892 209562 391904
rect 216674 391892 216680 391904
rect 216732 391892 216738 391944
rect 359734 391892 359740 391944
rect 359792 391932 359798 391944
rect 376938 391932 376944 391944
rect 359792 391904 376944 391932
rect 359792 391892 359798 391904
rect 376938 391892 376944 391904
rect 376996 391892 377002 391944
rect 207014 390464 207020 390516
rect 207072 390504 207078 390516
rect 216674 390504 216680 390516
rect 207072 390476 216680 390504
rect 207072 390464 207078 390476
rect 216674 390464 216680 390476
rect 216732 390464 216738 390516
rect 360194 390464 360200 390516
rect 360252 390504 360258 390516
rect 376938 390504 376944 390516
rect 360252 390476 376944 390504
rect 360252 390464 360258 390476
rect 376938 390464 376944 390476
rect 376996 390464 377002 390516
rect 57422 390328 57428 390380
rect 57480 390328 57486 390380
rect 57440 390108 57468 390328
rect 57422 390056 57428 390108
rect 57480 390056 57486 390108
rect 44082 389784 44088 389836
rect 44140 389824 44146 389836
rect 57606 389824 57612 389836
rect 44140 389796 57612 389824
rect 44140 389784 44146 389796
rect 57606 389784 57612 389796
rect 57664 389784 57670 389836
rect 206278 389172 206284 389224
rect 206336 389212 206342 389224
rect 207014 389212 207020 389224
rect 206336 389184 207020 389212
rect 206336 389172 206342 389184
rect 207014 389172 207020 389184
rect 207072 389172 207078 389224
rect 358078 389172 358084 389224
rect 358136 389212 358142 389224
rect 360194 389212 360200 389224
rect 358136 389184 360200 389212
rect 358136 389172 358142 389184
rect 360194 389172 360200 389184
rect 360252 389172 360258 389224
rect 46106 389104 46112 389156
rect 46164 389144 46170 389156
rect 57606 389144 57612 389156
rect 46164 389116 57612 389144
rect 46164 389104 46170 389116
rect 57606 389104 57612 389116
rect 57664 389104 57670 389156
rect 203886 389104 203892 389156
rect 203944 389144 203950 389156
rect 216674 389144 216680 389156
rect 203944 389116 216680 389144
rect 203944 389104 203950 389116
rect 216674 389104 216680 389116
rect 216732 389104 216738 389156
rect 359642 389104 359648 389156
rect 359700 389144 359706 389156
rect 376938 389144 376944 389156
rect 359700 389116 376944 389144
rect 359700 389104 359706 389116
rect 376938 389104 376944 389116
rect 376996 389104 377002 389156
rect 56778 388764 56784 388816
rect 56836 388804 56842 388816
rect 59538 388804 59544 388816
rect 56836 388776 59544 388804
rect 56836 388764 56842 388776
rect 59538 388764 59544 388776
rect 59596 388764 59602 388816
rect 57882 388424 57888 388476
rect 57940 388464 57946 388476
rect 58434 388464 58440 388476
rect 57940 388436 58440 388464
rect 57940 388424 57946 388436
rect 58434 388424 58440 388436
rect 58492 388424 58498 388476
rect 57330 388356 57336 388408
rect 57388 388396 57394 388408
rect 57514 388396 57520 388408
rect 57388 388368 57520 388396
rect 57388 388356 57394 388368
rect 57514 388356 57520 388368
rect 57572 388356 57578 388408
rect 216766 388356 216772 388408
rect 216824 388396 216830 388408
rect 217042 388396 217048 388408
rect 216824 388368 217048 388396
rect 216824 388356 216830 388368
rect 217042 388356 217048 388368
rect 217100 388356 217106 388408
rect 57238 387744 57244 387796
rect 57296 387784 57302 387796
rect 58526 387784 58532 387796
rect 57296 387756 58532 387784
rect 57296 387744 57302 387756
rect 58526 387744 58532 387756
rect 58584 387744 58590 387796
rect 372982 382236 372988 382288
rect 373040 382276 373046 382288
rect 376754 382276 376760 382288
rect 373040 382248 376760 382276
rect 373040 382236 373046 382248
rect 376754 382236 376760 382248
rect 376812 382236 376818 382288
rect 57422 381896 57428 381948
rect 57480 381936 57486 381948
rect 59354 381936 59360 381948
rect 57480 381908 59360 381936
rect 57480 381896 57486 381908
rect 59354 381896 59360 381908
rect 59412 381896 59418 381948
rect 55950 380944 55956 380996
rect 56008 380984 56014 380996
rect 59446 380984 59452 380996
rect 56008 380956 59452 380984
rect 56008 380944 56014 380956
rect 59446 380944 59452 380956
rect 59504 380944 59510 380996
rect 197170 380944 197176 380996
rect 197228 380984 197234 380996
rect 198182 380984 198188 380996
rect 197228 380956 198188 380984
rect 197228 380944 197234 380956
rect 198182 380944 198188 380956
rect 198240 380944 198246 380996
rect 57882 380876 57888 380928
rect 57940 380916 57946 380928
rect 60734 380916 60740 380928
rect 57940 380888 60740 380916
rect 57940 380876 57946 380888
rect 60734 380876 60740 380888
rect 60792 380876 60798 380928
rect 196986 380876 196992 380928
rect 197044 380916 197050 380928
rect 197998 380916 198004 380928
rect 197044 380888 198004 380916
rect 197044 380876 197050 380888
rect 197998 380876 198004 380888
rect 198056 380876 198062 380928
rect 198274 380876 198280 380928
rect 198332 380916 198338 380928
rect 199102 380916 199108 380928
rect 198332 380888 199108 380916
rect 198332 380876 198338 380888
rect 199102 380876 199108 380888
rect 199160 380876 199166 380928
rect 217594 380876 217600 380928
rect 217652 380916 217658 380928
rect 276014 380916 276020 380928
rect 217652 380888 276020 380916
rect 217652 380876 217658 380888
rect 276014 380876 276020 380888
rect 276072 380876 276078 380928
rect 376754 380876 376760 380928
rect 376812 380916 376818 380928
rect 421742 380916 421748 380928
rect 376812 380888 421748 380916
rect 376812 380876 376818 380888
rect 421742 380876 421748 380888
rect 421800 380876 421806 380928
rect 54294 380808 54300 380860
rect 54352 380848 54358 380860
rect 56594 380848 56600 380860
rect 54352 380820 56600 380848
rect 54352 380808 54358 380820
rect 56594 380808 56600 380820
rect 56652 380808 56658 380860
rect 216674 380848 216680 380860
rect 60016 380820 216680 380848
rect 48866 380740 48872 380792
rect 48924 380780 48930 380792
rect 60016 380780 60044 380820
rect 216674 380808 216680 380820
rect 216732 380808 216738 380860
rect 216858 380780 216864 380792
rect 48924 380752 60044 380780
rect 60200 380752 216864 380780
rect 48924 380740 48930 380752
rect 48774 380604 48780 380656
rect 48832 380644 48838 380656
rect 60200 380644 60228 380752
rect 216858 380740 216864 380752
rect 216916 380740 216922 380792
rect 364794 380740 364800 380792
rect 364852 380780 364858 380792
rect 379514 380780 379520 380792
rect 364852 380752 379520 380780
rect 364852 380740 364858 380752
rect 379514 380740 379520 380752
rect 379572 380740 379578 380792
rect 216950 380712 216956 380724
rect 48832 380616 60228 380644
rect 64846 380684 216956 380712
rect 48832 380604 48838 380616
rect 51626 380536 51632 380588
rect 51684 380576 51690 380588
rect 64846 380576 64874 380684
rect 216950 380672 216956 380684
rect 217008 380672 217014 380724
rect 373810 380672 373816 380724
rect 373868 380712 373874 380724
rect 378134 380712 378140 380724
rect 373868 380684 378140 380712
rect 373868 380672 373874 380684
rect 378134 380672 378140 380684
rect 378192 380712 378198 380724
rect 434346 380712 434352 380724
rect 378192 380684 434352 380712
rect 378192 380672 378198 380684
rect 434346 380672 434352 380684
rect 434404 380672 434410 380724
rect 155954 380604 155960 380656
rect 156012 380644 156018 380656
rect 204438 380644 204444 380656
rect 156012 380616 204444 380644
rect 156012 380604 156018 380616
rect 204438 380604 204444 380616
rect 204496 380604 204502 380656
rect 360746 380604 360752 380656
rect 360804 380644 360810 380656
rect 376662 380644 376668 380656
rect 360804 380616 376668 380644
rect 360804 380604 360810 380616
rect 376662 380604 376668 380616
rect 376720 380604 376726 380656
rect 377306 380604 377312 380656
rect 377364 380644 377370 380656
rect 425974 380644 425980 380656
rect 377364 380616 425980 380644
rect 377364 380604 377370 380616
rect 425974 380604 425980 380616
rect 426032 380604 426038 380656
rect 51684 380548 64874 380576
rect 51684 380536 51690 380548
rect 158530 380536 158536 380588
rect 158588 380576 158594 380588
rect 205910 380576 205916 380588
rect 158588 380548 205916 380576
rect 158588 380536 158594 380548
rect 205910 380536 205916 380548
rect 205968 380536 205974 380588
rect 207014 380536 207020 380588
rect 207072 380576 207078 380588
rect 213730 380576 213736 380588
rect 207072 380548 213736 380576
rect 207072 380536 207078 380548
rect 213730 380536 213736 380548
rect 213788 380536 213794 380588
rect 373626 380536 373632 380588
rect 373684 380576 373690 380588
rect 433610 380576 433616 380588
rect 373684 380548 433616 380576
rect 373684 380536 373690 380548
rect 433610 380536 433616 380548
rect 433668 380536 433674 380588
rect 58618 380468 58624 380520
rect 58676 380508 58682 380520
rect 105814 380508 105820 380520
rect 58676 380480 105820 380508
rect 58676 380468 58682 380480
rect 105814 380468 105820 380480
rect 105872 380468 105878 380520
rect 138474 380468 138480 380520
rect 138532 380508 138538 380520
rect 200390 380508 200396 380520
rect 138532 380480 200396 380508
rect 138532 380468 138538 380480
rect 200390 380468 200396 380480
rect 200448 380468 200454 380520
rect 202874 380468 202880 380520
rect 202932 380508 202938 380520
rect 213822 380508 213828 380520
rect 202932 380480 213828 380508
rect 202932 380468 202938 380480
rect 213822 380468 213828 380480
rect 213880 380468 213886 380520
rect 359458 380468 359464 380520
rect 359516 380508 359522 380520
rect 421098 380508 421104 380520
rect 359516 380480 421104 380508
rect 359516 380468 359522 380480
rect 421098 380468 421104 380480
rect 421156 380468 421162 380520
rect 59538 380400 59544 380452
rect 59596 380440 59602 380452
rect 118326 380440 118332 380452
rect 59596 380412 118332 380440
rect 59596 380400 59602 380412
rect 118326 380400 118332 380412
rect 118384 380400 118390 380452
rect 135898 380400 135904 380452
rect 135956 380440 135962 380452
rect 200666 380440 200672 380452
rect 135956 380412 200672 380440
rect 135956 380400 135962 380412
rect 200666 380400 200672 380412
rect 200724 380400 200730 380452
rect 202966 380400 202972 380452
rect 203024 380440 203030 380452
rect 274634 380440 274640 380452
rect 203024 380412 274640 380440
rect 203024 380400 203030 380412
rect 274634 380400 274640 380412
rect 274692 380400 274698 380452
rect 370314 380400 370320 380452
rect 370372 380440 370378 380452
rect 436002 380440 436008 380452
rect 370372 380412 436008 380440
rect 370372 380400 370378 380412
rect 436002 380400 436008 380412
rect 436060 380400 436066 380452
rect 52270 380332 52276 380384
rect 52328 380372 52334 380384
rect 113542 380372 113548 380384
rect 52328 380344 113548 380372
rect 52328 380332 52334 380344
rect 113542 380332 113548 380344
rect 113600 380332 113606 380384
rect 123570 380332 123576 380384
rect 123628 380372 123634 380384
rect 204530 380372 204536 380384
rect 123628 380344 204536 380372
rect 123628 380332 123634 380344
rect 204530 380332 204536 380344
rect 204588 380332 204594 380384
rect 208394 380332 208400 380384
rect 208452 380372 208458 380384
rect 218146 380372 218152 380384
rect 208452 380344 218152 380372
rect 208452 380332 208458 380344
rect 218146 380332 218152 380344
rect 218204 380332 218210 380384
rect 367554 380332 367560 380384
rect 367612 380372 367618 380384
rect 438486 380372 438492 380384
rect 367612 380344 438492 380372
rect 367612 380332 367618 380344
rect 438486 380332 438492 380344
rect 438544 380332 438550 380384
rect 48958 380264 48964 380316
rect 49016 380304 49022 380316
rect 110966 380304 110972 380316
rect 49016 380276 110972 380304
rect 49016 380264 49022 380276
rect 110966 380264 110972 380276
rect 111024 380264 111030 380316
rect 148594 380264 148600 380316
rect 148652 380304 148658 380316
rect 196894 380304 196900 380316
rect 148652 380276 196900 380304
rect 148652 380264 148658 380276
rect 196894 380264 196900 380276
rect 196952 380264 196958 380316
rect 201034 380264 201040 380316
rect 201092 380304 201098 380316
rect 295334 380304 295340 380316
rect 201092 380276 295340 380304
rect 201092 380264 201098 380276
rect 295334 380264 295340 380276
rect 295392 380264 295398 380316
rect 369670 380264 369676 380316
rect 369728 380304 369734 380316
rect 440878 380304 440884 380316
rect 369728 380276 440884 380304
rect 369728 380264 369734 380276
rect 440878 380264 440884 380276
rect 440936 380264 440942 380316
rect 58526 380196 58532 380248
rect 58584 380236 58590 380248
rect 120902 380236 120908 380248
rect 58584 380208 120908 380236
rect 58584 380196 58590 380208
rect 120902 380196 120908 380208
rect 120960 380196 120966 380248
rect 133506 380196 133512 380248
rect 133564 380236 133570 380248
rect 199194 380236 199200 380248
rect 133564 380208 199200 380236
rect 133564 380196 133570 380208
rect 199194 380196 199200 380208
rect 199252 380196 199258 380248
rect 200206 380196 200212 380248
rect 200264 380236 200270 380248
rect 301498 380236 301504 380248
rect 200264 380208 301504 380236
rect 200264 380196 200270 380208
rect 301498 380196 301504 380208
rect 301556 380196 301562 380248
rect 364886 380196 364892 380248
rect 364944 380236 364950 380248
rect 443454 380236 443460 380248
rect 364944 380208 443460 380236
rect 364944 380196 364950 380208
rect 443454 380196 443460 380208
rect 443512 380196 443518 380248
rect 54386 380128 54392 380180
rect 54444 380168 54450 380180
rect 115934 380168 115940 380180
rect 54444 380140 115940 380168
rect 54444 380128 54450 380140
rect 115934 380128 115940 380140
rect 115992 380128 115998 380180
rect 128354 380128 128360 380180
rect 128412 380168 128418 380180
rect 197906 380168 197912 380180
rect 128412 380140 197912 380168
rect 128412 380128 128418 380140
rect 197906 380128 197912 380140
rect 197964 380128 197970 380180
rect 201770 380128 201776 380180
rect 201828 380168 201834 380180
rect 311802 380168 311808 380180
rect 201828 380140 311808 380168
rect 201828 380128 201834 380140
rect 311802 380128 311808 380140
rect 311860 380128 311866 380180
rect 365622 380128 365628 380180
rect 365680 380168 365686 380180
rect 465902 380168 465908 380180
rect 365680 380140 465908 380168
rect 365680 380128 365686 380140
rect 465902 380128 465908 380140
rect 465960 380128 465966 380180
rect 160922 380060 160928 380112
rect 160980 380100 160986 380112
rect 207382 380100 207388 380112
rect 160980 380072 207388 380100
rect 160980 380060 160986 380072
rect 207382 380060 207388 380072
rect 207440 380060 207446 380112
rect 166074 379992 166080 380044
rect 166132 380032 166138 380044
rect 200574 380032 200580 380044
rect 166132 380004 200580 380032
rect 166132 379992 166138 380004
rect 200574 379992 200580 380004
rect 200632 379992 200638 380044
rect 213822 379992 213828 380044
rect 213880 380032 213886 380044
rect 235994 380032 236000 380044
rect 213880 380004 236000 380032
rect 213880 379992 213886 380004
rect 235994 379992 236000 380004
rect 236052 379992 236058 380044
rect 366266 379992 366272 380044
rect 366324 380032 366330 380044
rect 366324 380004 373994 380032
rect 366324 379992 366330 380004
rect 55674 379924 55680 379976
rect 55732 379964 55738 379976
rect 59630 379964 59636 379976
rect 55732 379936 59636 379964
rect 55732 379924 55738 379936
rect 59630 379924 59636 379936
rect 59688 379924 59694 379976
rect 163498 379924 163504 379976
rect 163556 379964 163562 379976
rect 197814 379964 197820 379976
rect 163556 379936 197820 379964
rect 163556 379924 163562 379936
rect 197814 379924 197820 379936
rect 197872 379924 197878 379976
rect 215294 379924 215300 379976
rect 215352 379964 215358 379976
rect 216398 379964 216404 379976
rect 215352 379936 216404 379964
rect 215352 379924 215358 379936
rect 216398 379924 216404 379936
rect 216456 379964 216462 379976
rect 237098 379964 237104 379976
rect 216456 379936 237104 379964
rect 216456 379924 216462 379936
rect 237098 379924 237104 379936
rect 237156 379924 237162 379976
rect 239950 379924 239956 379976
rect 240008 379964 240014 379976
rect 259454 379964 259460 379976
rect 240008 379936 259460 379964
rect 240008 379924 240014 379936
rect 259454 379924 259460 379936
rect 259512 379924 259518 379976
rect 212534 379856 212540 379908
rect 212592 379896 212598 379908
rect 217778 379896 217784 379908
rect 212592 379868 217784 379896
rect 212592 379856 212598 379868
rect 217778 379856 217784 379868
rect 217836 379856 217842 379908
rect 218146 379856 218152 379908
rect 218204 379896 218210 379908
rect 218330 379896 218336 379908
rect 218204 379868 218336 379896
rect 218204 379856 218210 379868
rect 218330 379856 218336 379868
rect 218388 379896 218394 379908
rect 244274 379896 244280 379908
rect 218388 379868 244280 379896
rect 218388 379856 218394 379868
rect 244274 379856 244280 379868
rect 244332 379856 244338 379908
rect 213730 379788 213736 379840
rect 213788 379828 213794 379840
rect 243078 379828 243084 379840
rect 213788 379800 243084 379828
rect 213788 379788 213794 379800
rect 243078 379788 243084 379800
rect 243136 379788 243142 379840
rect 215018 379720 215024 379772
rect 215076 379760 215082 379772
rect 215076 379732 219434 379760
rect 215076 379720 215082 379732
rect 207014 379652 207020 379704
rect 207072 379692 207078 379704
rect 208302 379692 208308 379704
rect 207072 379664 208308 379692
rect 207072 379652 207078 379664
rect 208302 379652 208308 379664
rect 208360 379692 208366 379704
rect 209406 379692 209412 379704
rect 208360 379664 209412 379692
rect 208360 379652 208366 379664
rect 209406 379652 209412 379664
rect 209464 379652 209470 379704
rect 212718 379652 212724 379704
rect 212776 379692 212782 379704
rect 219406 379692 219434 379732
rect 220722 379720 220728 379772
rect 220780 379760 220786 379772
rect 254486 379760 254492 379772
rect 220780 379732 254492 379760
rect 220780 379720 220786 379732
rect 254486 379720 254492 379732
rect 254544 379720 254550 379772
rect 373966 379760 373994 380004
rect 379514 379788 379520 379840
rect 379572 379828 379578 379840
rect 379882 379828 379888 379840
rect 379572 379800 379888 379828
rect 379572 379788 379578 379800
rect 379882 379788 379888 379800
rect 379940 379828 379946 379840
rect 408678 379828 408684 379840
rect 379940 379800 408684 379828
rect 379940 379788 379946 379800
rect 408678 379788 408684 379800
rect 408736 379788 408742 379840
rect 381078 379760 381084 379772
rect 373966 379732 381084 379760
rect 381078 379720 381084 379732
rect 381136 379760 381142 379772
rect 413462 379760 413468 379772
rect 381136 379732 413468 379760
rect 381136 379720 381142 379732
rect 413462 379720 413468 379732
rect 413520 379720 413526 379772
rect 256970 379692 256976 379704
rect 212776 379664 217732 379692
rect 219406 379664 256976 379692
rect 212776 379652 212782 379664
rect 204254 379516 204260 379568
rect 204312 379556 204318 379568
rect 215294 379556 215300 379568
rect 204312 379528 215300 379556
rect 204312 379516 204318 379528
rect 215294 379516 215300 379528
rect 215352 379516 215358 379568
rect 216950 379516 216956 379568
rect 217008 379556 217014 379568
rect 217594 379556 217600 379568
rect 217008 379528 217600 379556
rect 217008 379516 217014 379528
rect 217594 379516 217600 379528
rect 217652 379516 217658 379568
rect 217704 379556 217732 379664
rect 256970 379652 256976 379664
rect 257028 379652 257034 379704
rect 371050 379652 371056 379704
rect 371108 379692 371114 379704
rect 376846 379692 376852 379704
rect 371108 379664 376852 379692
rect 371108 379652 371114 379664
rect 376846 379652 376852 379664
rect 376904 379692 376910 379704
rect 377398 379692 377404 379704
rect 376904 379664 377404 379692
rect 376904 379652 376910 379664
rect 377398 379652 377404 379664
rect 377456 379652 377462 379704
rect 379238 379652 379244 379704
rect 379296 379692 379302 379704
rect 380894 379692 380900 379704
rect 379296 379664 380900 379692
rect 379296 379652 379302 379664
rect 380894 379652 380900 379664
rect 380952 379692 380958 379704
rect 425238 379692 425244 379704
rect 380952 379664 425244 379692
rect 380952 379652 380958 379664
rect 425238 379652 425244 379664
rect 425296 379652 425302 379704
rect 217778 379584 217784 379636
rect 217836 379624 217842 379636
rect 219710 379624 219716 379636
rect 217836 379596 219716 379624
rect 217836 379584 217842 379596
rect 219710 379584 219716 379596
rect 219768 379624 219774 379636
rect 220722 379624 220728 379636
rect 219768 379596 220728 379624
rect 219768 379584 219774 379596
rect 220722 379584 220728 379596
rect 220780 379584 220786 379636
rect 255866 379624 255872 379636
rect 220832 379596 255872 379624
rect 220832 379556 220860 379596
rect 255866 379584 255872 379596
rect 255924 379584 255930 379636
rect 376570 379584 376576 379636
rect 376628 379624 376634 379636
rect 422846 379624 422852 379636
rect 376628 379596 422852 379624
rect 376628 379584 376634 379596
rect 422846 379584 422852 379596
rect 422904 379584 422910 379636
rect 217704 379528 220860 379556
rect 221826 379516 221832 379568
rect 221884 379556 221890 379568
rect 265250 379556 265256 379568
rect 221884 379528 265256 379556
rect 221884 379516 221890 379528
rect 265250 379516 265256 379528
rect 265308 379516 265314 379568
rect 376662 379516 376668 379568
rect 376720 379556 376726 379568
rect 436922 379556 436928 379568
rect 376720 379528 436928 379556
rect 376720 379516 376726 379528
rect 436922 379516 436928 379528
rect 436980 379516 436986 379568
rect 86586 379448 86592 379500
rect 86644 379488 86650 379500
rect 208394 379488 208400 379500
rect 86644 379460 208400 379488
rect 86644 379448 86650 379460
rect 208394 379448 208400 379460
rect 208452 379448 208458 379500
rect 220630 379448 220636 379500
rect 220688 379488 220694 379500
rect 220688 379460 274588 379488
rect 220688 379448 220694 379460
rect 47762 379380 47768 379432
rect 47820 379420 47826 379432
rect 88334 379420 88340 379432
rect 47820 379392 88340 379420
rect 47820 379380 47826 379392
rect 88334 379380 88340 379392
rect 88392 379380 88398 379432
rect 92382 379380 92388 379432
rect 92440 379420 92446 379432
rect 212810 379420 212816 379432
rect 92440 379392 212816 379420
rect 92440 379380 92446 379392
rect 212810 379380 212816 379392
rect 212868 379420 212874 379432
rect 213822 379420 213828 379432
rect 212868 379392 213828 379420
rect 212868 379380 212874 379392
rect 213822 379380 213828 379392
rect 213880 379380 213886 379432
rect 215386 379380 215392 379432
rect 215444 379420 215450 379432
rect 219434 379420 219440 379432
rect 215444 379392 219440 379420
rect 215444 379380 215450 379392
rect 219434 379380 219440 379392
rect 219492 379420 219498 379432
rect 273254 379420 273260 379432
rect 219492 379392 273260 379420
rect 219492 379380 219498 379392
rect 273254 379380 273260 379392
rect 273312 379380 273318 379432
rect 274560 379420 274588 379460
rect 274634 379448 274640 379500
rect 274692 379488 274698 379500
rect 323302 379488 323308 379500
rect 274692 379460 323308 379488
rect 274692 379448 274698 379460
rect 323302 379448 323308 379460
rect 323360 379448 323366 379500
rect 368842 379448 368848 379500
rect 368900 379488 368906 379500
rect 439038 379488 439044 379500
rect 368900 379460 439044 379488
rect 368900 379448 368906 379460
rect 439038 379448 439044 379460
rect 439096 379448 439102 379500
rect 275646 379420 275652 379432
rect 274560 379392 275652 379420
rect 275646 379380 275652 379392
rect 275704 379380 275710 379432
rect 295334 379380 295340 379432
rect 295392 379420 295398 379432
rect 310974 379420 310980 379432
rect 295392 379392 310980 379420
rect 295392 379380 295398 379392
rect 310974 379380 310980 379392
rect 311032 379380 311038 379432
rect 311802 379380 311808 379432
rect 311860 379420 311866 379432
rect 315758 379420 315764 379432
rect 311860 379392 315764 379420
rect 311860 379380 311866 379392
rect 315758 379380 315764 379392
rect 315816 379380 315822 379432
rect 377398 379380 377404 379432
rect 377456 379420 377462 379432
rect 427446 379420 427452 379432
rect 377456 379392 427452 379420
rect 377456 379380 377462 379392
rect 427446 379380 427452 379392
rect 427504 379380 427510 379432
rect 88794 379312 88800 379364
rect 88852 379352 88858 379364
rect 209774 379352 209780 379364
rect 88852 379324 209780 379352
rect 88852 379312 88858 379324
rect 209774 379312 209780 379324
rect 209832 379352 209838 379364
rect 211062 379352 211068 379364
rect 209832 379324 211068 379352
rect 209832 379312 209838 379324
rect 211062 379312 211068 379324
rect 211120 379312 211126 379364
rect 220722 379312 220728 379364
rect 220780 379352 220786 379364
rect 274358 379352 274364 379364
rect 220780 379324 274364 379352
rect 220780 379312 220786 379324
rect 274358 379312 274364 379324
rect 274416 379312 274422 379364
rect 301498 379312 301504 379364
rect 301556 379352 301562 379364
rect 313366 379352 313372 379364
rect 301556 379324 313372 379352
rect 301556 379312 301562 379324
rect 313366 379312 313372 379324
rect 313424 379312 313430 379364
rect 375006 379312 375012 379364
rect 375064 379352 375070 379364
rect 408310 379352 408316 379364
rect 375064 379324 408316 379352
rect 375064 379312 375070 379324
rect 408310 379312 408316 379324
rect 408368 379312 408374 379364
rect 55766 379244 55772 379296
rect 55824 379284 55830 379296
rect 90634 379284 90640 379296
rect 55824 379256 90640 379284
rect 55824 379244 55830 379256
rect 90634 379244 90640 379256
rect 90692 379244 90698 379296
rect 90726 379244 90732 379296
rect 90784 379284 90790 379296
rect 209866 379284 209872 379296
rect 90784 379256 209872 379284
rect 90784 379244 90790 379256
rect 209866 379244 209872 379256
rect 209924 379284 209930 379296
rect 219618 379284 219624 379296
rect 209924 379256 219624 379284
rect 209924 379244 209930 379256
rect 219618 379244 219624 379256
rect 219676 379284 219682 379296
rect 220538 379284 220544 379296
rect 219676 379256 220544 379284
rect 219676 379244 219682 379256
rect 220538 379244 220544 379256
rect 220596 379244 220602 379296
rect 91370 379176 91376 379228
rect 91428 379216 91434 379228
rect 91428 379188 209774 379216
rect 91428 379176 91434 379188
rect 59722 379108 59728 379160
rect 59780 379148 59786 379160
rect 93486 379148 93492 379160
rect 59780 379120 93492 379148
rect 59780 379108 59786 379120
rect 93486 379108 93492 379120
rect 93544 379108 93550 379160
rect 93578 379108 93584 379160
rect 93636 379148 93642 379160
rect 195974 379148 195980 379160
rect 93636 379120 195980 379148
rect 93636 379108 93642 379120
rect 195974 379108 195980 379120
rect 196032 379108 196038 379160
rect 47670 379040 47676 379092
rect 47728 379080 47734 379092
rect 108206 379080 108212 379092
rect 47728 379052 108212 379080
rect 47728 379040 47734 379052
rect 108206 379040 108212 379052
rect 108264 379040 108270 379092
rect 112346 379040 112352 379092
rect 112404 379080 112410 379092
rect 205910 379080 205916 379092
rect 112404 379052 205916 379080
rect 112404 379040 112410 379052
rect 205910 379040 205916 379052
rect 205968 379040 205974 379092
rect 209746 379080 209774 379188
rect 213822 379176 213828 379228
rect 213880 379216 213886 379228
rect 220814 379216 220820 379228
rect 213880 379188 220820 379216
rect 213880 379176 213886 379188
rect 220814 379176 220820 379188
rect 220872 379216 220878 379228
rect 221918 379216 221924 379228
rect 220872 379188 221924 379216
rect 220872 379176 220878 379188
rect 221918 379176 221924 379188
rect 221976 379176 221982 379228
rect 211062 379108 211068 379160
rect 211120 379148 211126 379160
rect 219434 379148 219440 379160
rect 211120 379120 219440 379148
rect 211120 379108 211126 379120
rect 219434 379108 219440 379120
rect 219492 379148 219498 379160
rect 220170 379148 220176 379160
rect 219492 379120 220176 379148
rect 219492 379108 219498 379120
rect 220170 379108 220176 379120
rect 220228 379108 220234 379160
rect 220446 379108 220452 379160
rect 220504 379148 220510 379160
rect 220504 379120 229094 379148
rect 220504 379108 220510 379120
rect 211430 379080 211436 379092
rect 209746 379052 211436 379080
rect 211430 379040 211436 379052
rect 211488 379080 211494 379092
rect 221550 379080 221556 379092
rect 211488 379052 221556 379080
rect 211488 379040 211494 379052
rect 221550 379040 221556 379052
rect 221608 379040 221614 379092
rect 53558 378972 53564 379024
rect 53616 379012 53622 379024
rect 101030 379012 101036 379024
rect 53616 378984 101036 379012
rect 53616 378972 53622 378984
rect 101030 378972 101036 378984
rect 101088 378972 101094 379024
rect 195974 378972 195980 379024
rect 196032 379012 196038 379024
rect 197262 379012 197268 379024
rect 196032 378984 197268 379012
rect 196032 378972 196038 378984
rect 197262 378972 197268 378984
rect 197320 379012 197326 379024
rect 220906 379012 220912 379024
rect 197320 378984 220912 379012
rect 197320 378972 197326 378984
rect 220906 378972 220912 378984
rect 220964 379012 220970 379024
rect 222102 379012 222108 379024
rect 220964 378984 222108 379012
rect 220964 378972 220970 378984
rect 222102 378972 222108 378984
rect 222160 378972 222166 379024
rect 57146 378904 57152 378956
rect 57204 378944 57210 378956
rect 103514 378944 103520 378956
rect 57204 378916 103520 378944
rect 57204 378904 57210 378916
rect 103514 378904 103520 378916
rect 103572 378904 103578 378956
rect 205726 378904 205732 378956
rect 205784 378944 205790 378956
rect 206830 378944 206836 378956
rect 205784 378916 206836 378944
rect 205784 378904 205790 378916
rect 206830 378904 206836 378916
rect 206888 378944 206894 378956
rect 219526 378944 219532 378956
rect 206888 378916 219532 378944
rect 206888 378904 206894 378916
rect 219526 378904 219532 378916
rect 219584 378944 219590 378956
rect 220722 378944 220728 378956
rect 219584 378916 220728 378944
rect 219584 378904 219590 378916
rect 220722 378904 220728 378916
rect 220780 378904 220786 378956
rect 229066 378944 229094 379120
rect 371142 378972 371148 379024
rect 371200 379012 371206 379024
rect 381262 379012 381268 379024
rect 371200 378984 381268 379012
rect 371200 378972 371206 378984
rect 381262 378972 381268 378984
rect 381320 378972 381326 379024
rect 247586 378944 247592 378956
rect 229066 378916 247592 378944
rect 247586 378904 247592 378916
rect 247644 378904 247650 378956
rect 357894 378904 357900 378956
rect 357952 378944 357958 378956
rect 379514 378944 379520 378956
rect 357952 378916 379520 378944
rect 357952 378904 357958 378916
rect 379514 378904 379520 378916
rect 379572 378904 379578 378956
rect 50154 378836 50160 378888
rect 50212 378876 50218 378888
rect 98178 378876 98184 378888
rect 50212 378848 98184 378876
rect 50212 378836 50218 378848
rect 98178 378836 98184 378848
rect 98236 378836 98242 378888
rect 111242 378836 111248 378888
rect 111300 378876 111306 378888
rect 199010 378876 199016 378888
rect 111300 378848 199016 378876
rect 111300 378836 111306 378848
rect 199010 378836 199016 378848
rect 199068 378836 199074 378888
rect 219158 378836 219164 378888
rect 219216 378876 219222 378888
rect 245378 378876 245384 378888
rect 219216 378848 245384 378876
rect 219216 378836 219222 378848
rect 245378 378836 245384 378848
rect 245436 378836 245442 378888
rect 373718 378836 373724 378888
rect 373776 378876 373782 378888
rect 396166 378876 396172 378888
rect 373776 378848 396172 378876
rect 373776 378836 373782 378848
rect 396166 378836 396172 378848
rect 396224 378836 396230 378888
rect 108850 378768 108856 378820
rect 108908 378808 108914 378820
rect 208210 378808 208216 378820
rect 108908 378780 208216 378808
rect 108908 378768 108914 378780
rect 208210 378768 208216 378780
rect 208268 378808 208274 378820
rect 268654 378808 268660 378820
rect 208268 378780 268660 378808
rect 208268 378768 208274 378780
rect 268654 378768 268660 378780
rect 268712 378768 268718 378820
rect 359550 378768 359556 378820
rect 359608 378808 359614 378820
rect 375190 378808 375196 378820
rect 359608 378780 375196 378808
rect 359608 378768 359614 378780
rect 375190 378768 375196 378780
rect 375248 378768 375254 378820
rect 379698 378768 379704 378820
rect 379756 378808 379762 378820
rect 379974 378808 379980 378820
rect 379756 378780 379980 378808
rect 379756 378768 379762 378780
rect 379974 378768 379980 378780
rect 380032 378808 380038 378820
rect 405734 378808 405740 378820
rect 380032 378780 405740 378808
rect 380032 378768 380038 378780
rect 405734 378768 405740 378780
rect 405792 378768 405798 378820
rect 213454 378740 213460 378752
rect 200086 378712 213460 378740
rect 49050 378632 49056 378684
rect 49108 378672 49114 378684
rect 96062 378672 96068 378684
rect 49108 378644 96068 378672
rect 49108 378632 49114 378644
rect 96062 378632 96068 378644
rect 96120 378632 96126 378684
rect 115842 378632 115848 378684
rect 115900 378672 115906 378684
rect 200086 378672 200114 378712
rect 213454 378700 213460 378712
rect 213512 378740 213518 378752
rect 219802 378740 219808 378752
rect 213512 378712 219808 378740
rect 213512 378700 213518 378712
rect 219802 378700 219808 378712
rect 219860 378740 219866 378752
rect 220630 378740 220636 378752
rect 219860 378712 220636 378740
rect 219860 378700 219866 378712
rect 220630 378700 220636 378712
rect 220688 378700 220694 378752
rect 115900 378644 200114 378672
rect 115900 378632 115906 378644
rect 220170 378632 220176 378684
rect 220228 378672 220234 378684
rect 248598 378672 248604 378684
rect 220228 378644 248604 378672
rect 220228 378632 220234 378644
rect 248598 378632 248604 378644
rect 248656 378632 248662 378684
rect 46198 378564 46204 378616
rect 46256 378604 46262 378616
rect 46934 378604 46940 378616
rect 46256 378576 46940 378604
rect 46256 378564 46262 378576
rect 46934 378564 46940 378576
rect 46992 378564 46998 378616
rect 85482 378564 85488 378616
rect 85540 378604 85546 378616
rect 213638 378604 213644 378616
rect 85540 378576 213644 378604
rect 85540 378564 85546 378576
rect 213638 378564 213644 378576
rect 213696 378604 213702 378616
rect 219158 378604 219164 378616
rect 213696 378576 219164 378604
rect 213696 378564 213702 378576
rect 219158 378564 219164 378576
rect 219216 378564 219222 378616
rect 221090 378564 221096 378616
rect 221148 378604 221154 378616
rect 221550 378604 221556 378616
rect 221148 378576 221556 378604
rect 221148 378564 221154 378576
rect 221550 378564 221556 378576
rect 221608 378604 221614 378616
rect 251174 378604 251180 378616
rect 221608 378576 251180 378604
rect 221608 378564 221614 378576
rect 251174 378564 251180 378576
rect 251232 378564 251238 378616
rect 47578 378496 47584 378548
rect 47636 378536 47642 378548
rect 49050 378536 49056 378548
rect 47636 378508 49056 378536
rect 47636 378496 47642 378508
rect 49050 378496 49056 378508
rect 49108 378496 49114 378548
rect 114462 378496 114468 378548
rect 114520 378536 114526 378548
rect 205726 378536 205732 378548
rect 114520 378508 205732 378536
rect 114520 378496 114526 378508
rect 205726 378496 205732 378508
rect 205784 378496 205790 378548
rect 220538 378496 220544 378548
rect 220596 378536 220602 378548
rect 250070 378536 250076 378548
rect 220596 378508 250076 378536
rect 220596 378496 220602 378508
rect 250070 378496 250076 378508
rect 250128 378496 250134 378548
rect 374546 378496 374552 378548
rect 374604 378536 374610 378548
rect 375006 378536 375012 378548
rect 374604 378508 375012 378536
rect 374604 378496 374610 378508
rect 375006 378496 375012 378508
rect 375064 378536 375070 378548
rect 396074 378536 396080 378548
rect 375064 378508 396080 378536
rect 375064 378496 375070 378508
rect 396074 378496 396080 378508
rect 396132 378496 396138 378548
rect 199010 378428 199016 378480
rect 199068 378468 199074 378480
rect 209590 378468 209596 378480
rect 199068 378440 209596 378468
rect 199068 378428 199074 378440
rect 209590 378428 209596 378440
rect 209648 378468 209654 378480
rect 271046 378468 271052 378480
rect 209648 378440 271052 378468
rect 209648 378428 209654 378440
rect 271046 378428 271052 378440
rect 271104 378428 271110 378480
rect 381262 378428 381268 378480
rect 381320 378468 381326 378480
rect 412358 378468 412364 378480
rect 381320 378440 412364 378468
rect 381320 378428 381326 378440
rect 412358 378428 412364 378440
rect 412416 378428 412422 378480
rect 208394 378360 208400 378412
rect 208452 378400 208458 378412
rect 211614 378400 211620 378412
rect 208452 378372 211620 378400
rect 208452 378360 208458 378372
rect 211614 378360 211620 378372
rect 211672 378400 211678 378412
rect 245654 378400 245660 378412
rect 211672 378372 245660 378400
rect 211672 378360 211678 378372
rect 245654 378360 245660 378372
rect 245712 378360 245718 378412
rect 379514 378360 379520 378412
rect 379572 378400 379578 378412
rect 379790 378400 379796 378412
rect 379572 378372 379796 378400
rect 379572 378360 379578 378372
rect 379790 378360 379796 378372
rect 379848 378400 379854 378412
rect 411254 378400 411260 378412
rect 379848 378372 411260 378400
rect 379848 378360 379854 378372
rect 411254 378360 411260 378372
rect 411312 378360 411318 378412
rect 113450 378292 113456 378344
rect 113508 378332 113514 378344
rect 215386 378332 215392 378344
rect 113508 378304 215392 378332
rect 113508 378292 113514 378304
rect 215386 378292 215392 378304
rect 215444 378292 215450 378344
rect 221918 378292 221924 378344
rect 221976 378332 221982 378344
rect 252278 378332 252284 378344
rect 221976 378304 252284 378332
rect 221976 378292 221982 378304
rect 252278 378292 252284 378304
rect 252336 378292 252342 378344
rect 342254 378292 342260 378344
rect 342312 378332 342318 378344
rect 343174 378332 343180 378344
rect 342312 378304 343180 378332
rect 342312 378292 342318 378304
rect 343174 378292 343180 378304
rect 343232 378332 343238 378344
rect 359366 378332 359372 378344
rect 343232 378304 359372 378332
rect 343232 378292 343238 378304
rect 359366 378292 359372 378304
rect 359424 378332 359430 378344
rect 359424 378304 364334 378332
rect 359424 378292 359430 378304
rect 49050 378224 49056 378276
rect 49108 378264 49114 378276
rect 81434 378264 81440 378276
rect 49108 378236 81440 378264
rect 49108 378224 49114 378236
rect 81434 378224 81440 378236
rect 81492 378224 81498 378276
rect 205910 378224 205916 378276
rect 205968 378264 205974 378276
rect 206922 378264 206928 378276
rect 205968 378236 206928 378264
rect 205968 378224 205974 378236
rect 206922 378224 206928 378236
rect 206980 378264 206986 378276
rect 211706 378264 211712 378276
rect 206980 378236 211712 378264
rect 206980 378224 206986 378236
rect 211706 378224 211712 378236
rect 211764 378264 211770 378276
rect 271966 378264 271972 378276
rect 211764 378236 271972 378264
rect 211764 378224 211770 378236
rect 271966 378224 271972 378236
rect 272024 378224 272030 378276
rect 276014 378224 276020 378276
rect 276072 378264 276078 378276
rect 277026 378264 277032 378276
rect 276072 378236 277032 378264
rect 276072 378224 276078 378236
rect 277026 378224 277032 378236
rect 277084 378264 277090 378276
rect 356606 378264 356612 378276
rect 277084 378236 356612 378264
rect 277084 378224 277090 378236
rect 356606 378224 356612 378236
rect 356664 378224 356670 378276
rect 364306 378264 364334 378304
rect 375190 378292 375196 378344
rect 375248 378332 375254 378344
rect 407574 378332 407580 378344
rect 375248 378304 407580 378332
rect 375248 378292 375254 378304
rect 407574 378292 407580 378304
rect 407632 378292 407638 378344
rect 439038 378292 439044 378344
rect 439096 378332 439102 378344
rect 516594 378332 516600 378344
rect 439096 378304 516600 378332
rect 439096 378292 439102 378304
rect 516594 378292 516600 378304
rect 516652 378292 516658 378344
rect 503070 378264 503076 378276
rect 364306 378236 503076 378264
rect 503070 378224 503076 378236
rect 503128 378264 503134 378276
rect 517606 378264 517612 378276
rect 503128 378236 517612 378264
rect 503128 378224 503134 378236
rect 517606 378224 517612 378236
rect 517664 378264 517670 378276
rect 580258 378264 580264 378276
rect 517664 378236 580264 378264
rect 517664 378224 517670 378236
rect 580258 378224 580264 378236
rect 580316 378224 580322 378276
rect 46934 378156 46940 378208
rect 46992 378196 46998 378208
rect 80330 378196 80336 378208
rect 46992 378168 80336 378196
rect 46992 378156 46998 378168
rect 80330 378156 80336 378168
rect 80388 378156 80394 378208
rect 87690 378156 87696 378208
rect 87748 378196 87754 378208
rect 219802 378196 219808 378208
rect 87748 378168 219808 378196
rect 87748 378156 87754 378168
rect 219802 378156 219808 378168
rect 219860 378196 219866 378208
rect 220446 378196 220452 378208
rect 219860 378168 220452 378196
rect 219860 378156 219866 378168
rect 220446 378156 220452 378168
rect 220504 378156 220510 378208
rect 222102 378156 222108 378208
rect 222160 378196 222166 378208
rect 253382 378196 253388 378208
rect 222160 378168 253388 378196
rect 222160 378156 222166 378168
rect 253382 378156 253388 378168
rect 253440 378156 253446 378208
rect 273254 378156 273260 378208
rect 273312 378196 273318 378208
rect 303062 378196 303068 378208
rect 273312 378168 303068 378196
rect 273312 378156 273318 378168
rect 303062 378156 303068 378168
rect 303120 378156 303126 378208
rect 343542 378156 343548 378208
rect 343600 378196 343606 378208
rect 503530 378196 503536 378208
rect 343600 378168 503536 378196
rect 343600 378156 343606 378168
rect 503530 378156 503536 378168
rect 503588 378196 503594 378208
rect 517698 378196 517704 378208
rect 503588 378168 517704 378196
rect 503588 378156 503594 378168
rect 517698 378156 517704 378168
rect 517756 378196 517762 378208
rect 580166 378196 580172 378208
rect 517756 378168 580172 378196
rect 517756 378156 517762 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 196710 378088 196716 378140
rect 196768 378128 196774 378140
rect 287606 378128 287612 378140
rect 196768 378100 287612 378128
rect 196768 378088 196774 378100
rect 287606 378088 287612 378100
rect 287664 378088 287670 378140
rect 367002 378088 367008 378140
rect 367060 378128 367066 378140
rect 374546 378128 374552 378140
rect 367060 378100 374552 378128
rect 367060 378088 367066 378100
rect 374546 378088 374552 378100
rect 374604 378088 374610 378140
rect 216766 378020 216772 378072
rect 216824 378060 216830 378072
rect 217318 378060 217324 378072
rect 216824 378032 217324 378060
rect 216824 378020 216830 378032
rect 217318 378020 217324 378032
rect 217376 378020 217382 378072
rect 217502 378020 217508 378072
rect 217560 378060 217566 378072
rect 308398 378060 308404 378072
rect 217560 378032 308404 378060
rect 217560 378020 217566 378032
rect 308398 378020 308404 378032
rect 308456 378020 308462 378072
rect 357250 378020 357256 378072
rect 357308 378060 357314 378072
rect 458358 378060 458364 378072
rect 357308 378032 458364 378060
rect 357308 378020 357314 378032
rect 458358 378020 458364 378032
rect 458416 378020 458422 378072
rect 43346 377952 43352 378004
rect 43404 377992 43410 378004
rect 199654 377992 199660 378004
rect 43404 377964 199660 377992
rect 43404 377952 43410 377964
rect 199654 377952 199660 377964
rect 199712 377952 199718 378004
rect 201586 377952 201592 378004
rect 201644 377992 201650 378004
rect 318334 377992 318340 378004
rect 201644 377964 318340 377992
rect 201644 377952 201650 377964
rect 318334 377952 318340 377964
rect 318392 377952 318398 378004
rect 366174 377952 366180 378004
rect 366232 377992 366238 378004
rect 452746 377992 452752 378004
rect 366232 377964 452752 377992
rect 366232 377952 366238 377964
rect 452746 377952 452752 377964
rect 452804 377952 452810 378004
rect 44726 377884 44732 377936
rect 44784 377924 44790 377936
rect 183462 377924 183468 377936
rect 44784 377896 183468 377924
rect 44784 377884 44790 377896
rect 183462 377884 183468 377896
rect 183520 377884 183526 377936
rect 198826 377884 198832 377936
rect 198884 377924 198890 377936
rect 300854 377924 300860 377936
rect 198884 377896 300860 377924
rect 198884 377884 198890 377896
rect 300854 377884 300860 377896
rect 300912 377884 300918 377936
rect 361298 377884 361304 377936
rect 361356 377924 361362 377936
rect 448146 377924 448152 377936
rect 361356 377896 448152 377924
rect 361356 377884 361362 377896
rect 448146 377884 448152 377896
rect 448204 377884 448210 377936
rect 54478 377816 54484 377868
rect 54536 377856 54542 377868
rect 182266 377856 182272 377868
rect 54536 377828 182272 377856
rect 54536 377816 54542 377828
rect 182266 377816 182272 377828
rect 182324 377816 182330 377868
rect 197538 377816 197544 377868
rect 197596 377856 197602 377868
rect 298094 377856 298100 377868
rect 197596 377828 298100 377856
rect 197596 377816 197602 377828
rect 298094 377816 298100 377828
rect 298152 377816 298158 377868
rect 364242 377816 364248 377868
rect 364300 377856 364306 377868
rect 450998 377856 451004 377868
rect 364300 377828 451004 377856
rect 364300 377816 364306 377828
rect 450998 377816 451004 377828
rect 451056 377816 451062 377868
rect 197446 377748 197452 377800
rect 197504 377788 197510 377800
rect 295886 377788 295892 377800
rect 197504 377760 295892 377788
rect 197504 377748 197510 377760
rect 295886 377748 295892 377760
rect 295944 377748 295950 377800
rect 362126 377748 362132 377800
rect 362184 377788 362190 377800
rect 445846 377788 445852 377800
rect 362184 377760 445852 377788
rect 362184 377748 362190 377760
rect 445846 377748 445852 377760
rect 445904 377748 445910 377800
rect 197354 377680 197360 377732
rect 197412 377720 197418 377732
rect 293310 377720 293316 377732
rect 197412 377692 293316 377720
rect 197412 377680 197418 377692
rect 293310 377680 293316 377692
rect 293368 377680 293374 377732
rect 372430 377680 372436 377732
rect 372488 377720 372494 377732
rect 455506 377720 455512 377732
rect 372488 377692 455512 377720
rect 372488 377680 372494 377692
rect 455506 377680 455512 377692
rect 455564 377680 455570 377732
rect 196802 377612 196808 377664
rect 196860 377652 196866 377664
rect 290918 377652 290924 377664
rect 196860 377624 290924 377652
rect 196860 377612 196866 377624
rect 290918 377612 290924 377624
rect 290976 377612 290982 377664
rect 357066 377612 357072 377664
rect 357124 377652 357130 377664
rect 423398 377652 423404 377664
rect 357124 377624 423404 377652
rect 357124 377612 357130 377624
rect 423398 377612 423404 377624
rect 423456 377612 423462 377664
rect 196618 377544 196624 377596
rect 196676 377584 196682 377596
rect 285950 377584 285956 377596
rect 196676 377556 285956 377584
rect 196676 377544 196682 377556
rect 285950 377544 285956 377556
rect 286008 377544 286014 377596
rect 357986 377544 357992 377596
rect 358044 377584 358050 377596
rect 410610 377584 410616 377596
rect 358044 377556 410616 377584
rect 358044 377544 358050 377556
rect 410610 377544 410616 377556
rect 410668 377544 410674 377596
rect 143626 377476 143632 377528
rect 143684 377516 143690 377528
rect 205818 377516 205824 377528
rect 143684 377488 205824 377516
rect 143684 377476 143690 377488
rect 205818 377476 205824 377488
rect 205876 377476 205882 377528
rect 217410 377476 217416 377528
rect 217468 377516 217474 377528
rect 305730 377516 305736 377528
rect 217468 377488 305736 377516
rect 217468 377476 217474 377488
rect 305730 377476 305736 377488
rect 305788 377476 305794 377528
rect 361482 377476 361488 377528
rect 361540 377516 361546 377528
rect 371142 377516 371148 377528
rect 361540 377488 371148 377516
rect 361540 377476 361546 377488
rect 371142 377476 371148 377488
rect 371200 377476 371206 377528
rect 375098 377476 375104 377528
rect 375156 377516 375162 377528
rect 413094 377516 413100 377528
rect 375156 377488 413100 377516
rect 375156 377476 375162 377488
rect 413094 377476 413100 377488
rect 413152 377476 413158 377528
rect 197078 377408 197084 377460
rect 197136 377448 197142 377460
rect 277854 377448 277860 377460
rect 197136 377420 277860 377448
rect 197136 377408 197142 377420
rect 277854 377408 277860 377420
rect 277912 377408 277918 377460
rect 363506 377408 363512 377460
rect 363564 377448 363570 377460
rect 379974 377448 379980 377460
rect 363564 377420 379980 377448
rect 363564 377408 363570 377420
rect 379974 377408 379980 377420
rect 380032 377448 380038 377460
rect 414566 377448 414572 377460
rect 380032 377420 414572 377448
rect 380032 377408 380038 377420
rect 414566 377408 414572 377420
rect 414624 377408 414630 377460
rect 146018 377340 146024 377392
rect 146076 377380 146082 377392
rect 207290 377380 207296 377392
rect 146076 377352 207296 377380
rect 146076 377340 146082 377352
rect 207290 377340 207296 377352
rect 207348 377340 207354 377392
rect 212350 377340 212356 377392
rect 212408 377380 212414 377392
rect 280798 377380 280804 377392
rect 212408 377352 280804 377380
rect 212408 377340 212414 377352
rect 280798 377340 280804 377352
rect 280856 377340 280862 377392
rect 371142 377340 371148 377392
rect 371200 377380 371206 377392
rect 402974 377380 402980 377392
rect 371200 377352 402980 377380
rect 371200 377340 371206 377352
rect 402974 377340 402980 377352
rect 403032 377340 403038 377392
rect 44634 377272 44640 377324
rect 44692 377312 44698 377324
rect 217318 377312 217324 377324
rect 44692 377284 217324 377312
rect 44692 377272 44698 377284
rect 217318 377272 217324 377284
rect 217376 377272 217382 377324
rect 369026 377272 369032 377324
rect 369084 377312 369090 377324
rect 379238 377312 379244 377324
rect 369084 377284 379244 377312
rect 369084 377272 369090 377284
rect 379238 377272 379244 377284
rect 379296 377312 379302 377324
rect 409966 377312 409972 377324
rect 379296 377284 409972 377312
rect 379296 377272 379302 377284
rect 409966 377272 409972 377284
rect 410024 377272 410030 377324
rect 141050 377204 141056 377256
rect 141108 377244 141114 377256
rect 201862 377244 201868 377256
rect 141108 377216 201868 377244
rect 141108 377204 141114 377216
rect 201862 377204 201868 377216
rect 201920 377204 201926 377256
rect 364150 377204 364156 377256
rect 364208 377244 364214 377256
rect 474734 377244 474740 377256
rect 364208 377216 474740 377244
rect 364208 377204 364214 377216
rect 474734 377204 474740 377216
rect 474792 377204 474798 377256
rect 153562 377136 153568 377188
rect 153620 377176 153626 377188
rect 200482 377176 200488 377188
rect 153620 377148 200488 377176
rect 153620 377136 153626 377148
rect 200482 377136 200488 377148
rect 200540 377136 200546 377188
rect 150986 377068 150992 377120
rect 151044 377108 151050 377120
rect 198182 377108 198188 377120
rect 151044 377080 198188 377108
rect 151044 377068 151050 377080
rect 198182 377068 198188 377080
rect 198240 377068 198246 377120
rect 47394 377000 47400 377052
rect 47452 377040 47458 377052
rect 217686 377040 217692 377052
rect 47452 377012 217692 377040
rect 47452 377000 47458 377012
rect 217686 377000 217692 377012
rect 217744 377000 217750 377052
rect 77202 376660 77208 376712
rect 77260 376700 77266 376712
rect 204254 376700 204260 376712
rect 77260 376672 204260 376700
rect 77260 376660 77266 376672
rect 204254 376660 204260 376672
rect 204312 376660 204318 376712
rect 213086 376660 213092 376712
rect 213144 376700 213150 376712
rect 283006 376700 283012 376712
rect 213144 376672 283012 376700
rect 213144 376660 213150 376672
rect 283006 376660 283012 376672
rect 283064 376660 283070 376712
rect 361390 376660 361396 376712
rect 361448 376700 361454 376712
rect 473446 376700 473452 376712
rect 361448 376672 473452 376700
rect 361448 376660 361454 376672
rect 473446 376660 473452 376672
rect 473504 376660 473510 376712
rect 201494 376592 201500 376644
rect 201552 376632 201558 376644
rect 320910 376632 320916 376644
rect 201552 376604 320916 376632
rect 201552 376592 201558 376604
rect 320910 376592 320916 376604
rect 320968 376592 320974 376644
rect 366910 376592 366916 376644
rect 366968 376632 366974 376644
rect 477586 376632 477592 376644
rect 366968 376604 477592 376632
rect 366968 376592 366974 376604
rect 477586 376592 477592 376604
rect 477644 376592 477650 376644
rect 125962 376524 125968 376576
rect 126020 376564 126026 376576
rect 203150 376564 203156 376576
rect 126020 376536 203156 376564
rect 126020 376524 126026 376536
rect 203150 376524 203156 376536
rect 203208 376524 203214 376576
rect 203978 376524 203984 376576
rect 204036 376564 204042 376576
rect 273438 376564 273444 376576
rect 204036 376536 273444 376564
rect 204036 376524 204042 376536
rect 273438 376524 273444 376536
rect 273496 376524 273502 376576
rect 362862 376524 362868 376576
rect 362920 376564 362926 376576
rect 470870 376564 470876 376576
rect 362920 376536 470876 376564
rect 362920 376524 362926 376536
rect 470870 376524 470876 376536
rect 470928 376524 470934 376576
rect 97718 376456 97724 376508
rect 97776 376496 97782 376508
rect 214466 376496 214472 376508
rect 97776 376468 214472 376496
rect 97776 376456 97782 376468
rect 214466 376456 214472 376468
rect 214524 376496 214530 376508
rect 215018 376496 215024 376508
rect 214524 376468 215024 376496
rect 214524 376456 214530 376468
rect 215018 376456 215024 376468
rect 215076 376456 215082 376508
rect 215846 376456 215852 376508
rect 215904 376496 215910 376508
rect 270954 376496 270960 376508
rect 215904 376468 270960 376496
rect 215904 376456 215910 376468
rect 270954 376456 270960 376468
rect 271012 376456 271018 376508
rect 376478 376456 376484 376508
rect 376536 376496 376542 376508
rect 483382 376496 483388 376508
rect 376536 376468 483388 376496
rect 376536 376456 376542 376468
rect 483382 376456 483388 376468
rect 483440 376456 483446 376508
rect 210234 376388 210240 376440
rect 210292 376428 210298 376440
rect 263594 376428 263600 376440
rect 210292 376400 263600 376428
rect 210292 376388 210298 376400
rect 263594 376388 263600 376400
rect 263652 376388 263658 376440
rect 369578 376388 369584 376440
rect 369636 376428 369642 376440
rect 467926 376428 467932 376440
rect 369636 376400 467932 376428
rect 369636 376388 369642 376400
rect 467926 376388 467932 376400
rect 467984 376388 467990 376440
rect 214374 376320 214380 376372
rect 214432 376360 214438 376372
rect 268102 376360 268108 376372
rect 214432 376332 268108 376360
rect 214432 376320 214438 376332
rect 268102 376320 268108 376332
rect 268160 376320 268166 376372
rect 368290 376320 368296 376372
rect 368348 376360 368354 376372
rect 463510 376360 463516 376372
rect 368348 376332 463516 376360
rect 368348 376320 368354 376332
rect 463510 376320 463516 376332
rect 463568 376320 463574 376372
rect 131022 376252 131028 376304
rect 131080 376292 131086 376304
rect 205634 376292 205640 376304
rect 131080 376264 205640 376292
rect 131080 376252 131086 376264
rect 205634 376252 205640 376264
rect 205692 376252 205698 376304
rect 213362 376252 213368 376304
rect 213420 376292 213426 376304
rect 260926 376292 260932 376304
rect 213420 376264 260932 376292
rect 213420 376252 213426 376264
rect 260926 376252 260932 376264
rect 260984 376252 260990 376304
rect 358538 376252 358544 376304
rect 358596 376292 358602 376304
rect 418246 376292 418252 376304
rect 358596 376264 418252 376292
rect 358596 376252 358602 376264
rect 418246 376252 418252 376264
rect 418304 376252 418310 376304
rect 211522 376184 211528 376236
rect 211580 376224 211586 376236
rect 258350 376224 258356 376236
rect 211580 376196 258356 376224
rect 211580 376184 211586 376196
rect 258350 376184 258356 376196
rect 258408 376184 258414 376236
rect 375282 376184 375288 376236
rect 375340 376224 375346 376236
rect 430666 376224 430672 376236
rect 375340 376196 430672 376224
rect 375340 376184 375346 376196
rect 430666 376184 430672 376196
rect 430724 376184 430730 376236
rect 94682 376116 94688 376168
rect 94740 376156 94746 376168
rect 212534 376156 212540 376168
rect 94740 376128 212540 376156
rect 94740 376116 94746 376128
rect 212534 376116 212540 376128
rect 212592 376116 212598 376168
rect 214006 376116 214012 376168
rect 214064 376156 214070 376168
rect 216306 376156 216312 376168
rect 214064 376128 216312 376156
rect 214064 376116 214070 376128
rect 216306 376116 216312 376128
rect 216364 376116 216370 376168
rect 219250 376116 219256 376168
rect 219308 376156 219314 376168
rect 265342 376156 265348 376168
rect 219308 376128 265348 376156
rect 219308 376116 219314 376128
rect 265342 376116 265348 376128
rect 265400 376116 265406 376168
rect 373166 376116 373172 376168
rect 373224 376156 373230 376168
rect 428182 376156 428188 376168
rect 373224 376128 428188 376156
rect 373224 376116 373230 376128
rect 428182 376116 428188 376128
rect 428240 376116 428246 376168
rect 202138 376048 202144 376100
rect 202196 376088 202202 376100
rect 248230 376088 248236 376100
rect 202196 376060 248236 376088
rect 202196 376048 202202 376060
rect 248230 376048 248236 376060
rect 248288 376048 248294 376100
rect 371786 376048 371792 376100
rect 371844 376088 371850 376100
rect 416038 376088 416044 376100
rect 371844 376060 416044 376088
rect 371844 376048 371850 376060
rect 416038 376048 416044 376060
rect 416096 376048 416102 376100
rect 216214 375980 216220 376032
rect 216272 376020 216278 376032
rect 255958 376020 255964 376032
rect 216272 375992 255964 376020
rect 216272 375980 216278 375992
rect 255958 375980 255964 375992
rect 256016 375980 256022 376032
rect 365530 375980 365536 376032
rect 365588 376020 365594 376032
rect 374546 376020 374552 376032
rect 365588 375992 374552 376020
rect 365588 375980 365594 375992
rect 374546 375980 374552 375992
rect 374604 376020 374610 376032
rect 415394 376020 415400 376032
rect 374604 375992 415400 376020
rect 374604 375980 374610 375992
rect 415394 375980 415400 375992
rect 415452 375980 415458 376032
rect 208946 375912 208952 375964
rect 209004 375952 209010 375964
rect 253566 375952 253572 375964
rect 209004 375924 253572 375952
rect 209004 375912 209010 375924
rect 253566 375912 253572 375924
rect 253624 375912 253630 375964
rect 374454 375912 374460 375964
rect 374512 375952 374518 375964
rect 377306 375952 377312 375964
rect 374512 375924 377312 375952
rect 374512 375912 374518 375924
rect 377306 375912 377312 375924
rect 377364 375952 377370 375964
rect 403618 375952 403624 375964
rect 377364 375924 403624 375952
rect 377364 375912 377370 375924
rect 403618 375912 403624 375924
rect 403676 375912 403682 375964
rect 99466 375844 99472 375896
rect 99524 375884 99530 375896
rect 214006 375884 214012 375896
rect 99524 375856 214012 375884
rect 99524 375844 99530 375856
rect 214006 375844 214012 375856
rect 214064 375844 214070 375896
rect 215110 375844 215116 375896
rect 215168 375884 215174 375896
rect 250622 375884 250628 375896
rect 215168 375856 250628 375884
rect 215168 375844 215174 375856
rect 250622 375844 250628 375856
rect 250680 375844 250686 375896
rect 239950 375816 239956 375828
rect 219406 375788 239956 375816
rect 104066 375708 104072 375760
rect 104124 375748 104130 375760
rect 216582 375748 216588 375760
rect 104124 375720 216588 375748
rect 104124 375708 104130 375720
rect 216582 375708 216588 375720
rect 216640 375748 216646 375760
rect 217226 375748 217232 375760
rect 216640 375720 217232 375748
rect 216640 375708 216646 375720
rect 217226 375708 217232 375720
rect 217284 375708 217290 375760
rect 100754 375640 100760 375692
rect 100812 375680 100818 375692
rect 216490 375680 216496 375692
rect 100812 375652 216496 375680
rect 100812 375640 100818 375652
rect 216490 375640 216496 375652
rect 216548 375640 216554 375692
rect 216306 375572 216312 375624
rect 216364 375612 216370 375624
rect 219406 375612 219434 375788
rect 239950 375776 239956 375788
rect 240008 375776 240014 375828
rect 216364 375584 219434 375612
rect 216364 375572 216370 375584
rect 357066 375408 357072 375420
rect 280080 375380 357072 375408
rect 101950 375300 101956 375352
rect 102008 375340 102014 375352
rect 213914 375340 213920 375352
rect 102008 375312 213920 375340
rect 102008 375300 102014 375312
rect 213914 375300 213920 375312
rect 213972 375300 213978 375352
rect 218054 375300 218060 375352
rect 218112 375340 218118 375352
rect 218238 375340 218244 375352
rect 218112 375312 218244 375340
rect 218112 375300 218118 375312
rect 218238 375300 218244 375312
rect 218296 375340 218302 375352
rect 219342 375340 219348 375352
rect 218296 375312 219348 375340
rect 218296 375300 218302 375312
rect 219342 375300 219348 375312
rect 219400 375340 219406 375352
rect 266354 375340 266360 375352
rect 219400 375312 266360 375340
rect 219400 375300 219406 375312
rect 266354 375300 266360 375312
rect 266412 375300 266418 375352
rect 215110 375232 215116 375284
rect 215168 375272 215174 375284
rect 215478 375272 215484 375284
rect 215168 375244 215484 375272
rect 215168 375232 215174 375244
rect 215478 375232 215484 375244
rect 215536 375272 215542 375284
rect 262766 375272 262772 375284
rect 215536 375244 262772 375272
rect 215536 375232 215542 375244
rect 262766 375232 262772 375244
rect 262824 375232 262830 375284
rect 107562 375164 107568 375216
rect 107620 375204 107626 375216
rect 207014 375204 207020 375216
rect 107620 375176 207020 375204
rect 107620 375164 107626 375176
rect 207014 375164 207020 375176
rect 207072 375164 207078 375216
rect 208302 375164 208308 375216
rect 208360 375204 208366 375216
rect 279142 375204 279148 375216
rect 208360 375176 279148 375204
rect 208360 375164 208366 375176
rect 279142 375164 279148 375176
rect 279200 375204 279206 375216
rect 280080 375204 280108 375380
rect 357066 375368 357072 375380
rect 357124 375368 357130 375420
rect 374362 375368 374368 375420
rect 374420 375408 374426 375420
rect 375466 375408 375472 375420
rect 374420 375380 375472 375408
rect 374420 375368 374426 375380
rect 375466 375368 375472 375380
rect 375524 375368 375530 375420
rect 368934 375300 368940 375352
rect 368992 375340 368998 375352
rect 369578 375340 369584 375352
rect 368992 375312 369584 375340
rect 368992 375300 368998 375312
rect 369578 375300 369584 375312
rect 369636 375300 369642 375352
rect 428274 375340 428280 375352
rect 369826 375312 428280 375340
rect 369596 375272 369624 375300
rect 369826 375272 369854 375312
rect 428274 375300 428280 375312
rect 428332 375300 428338 375352
rect 369596 375244 369854 375272
rect 373074 375232 373080 375284
rect 373132 375272 373138 375284
rect 431126 375272 431132 375284
rect 373132 375244 431132 375272
rect 373132 375232 373138 375244
rect 431126 375232 431132 375244
rect 431184 375232 431190 375284
rect 279200 375176 280108 375204
rect 279200 375164 279206 375176
rect 367646 375164 367652 375216
rect 367704 375204 367710 375216
rect 370038 375204 370044 375216
rect 367704 375176 370044 375204
rect 367704 375164 367710 375176
rect 370038 375164 370044 375176
rect 370096 375164 370102 375216
rect 375466 375164 375472 375216
rect 375524 375204 375530 375216
rect 432230 375204 432236 375216
rect 375524 375176 432236 375204
rect 375524 375164 375530 375176
rect 432230 375164 432236 375176
rect 432288 375164 432294 375216
rect 213914 375096 213920 375148
rect 213972 375136 213978 375148
rect 217502 375136 217508 375148
rect 213972 375108 217508 375136
rect 213972 375096 213978 375108
rect 217502 375096 217508 375108
rect 217560 375136 217566 375148
rect 261662 375136 261668 375148
rect 217560 375108 261668 375136
rect 217560 375096 217566 375108
rect 261662 375096 261668 375108
rect 261720 375096 261726 375148
rect 379330 375096 379336 375148
rect 379388 375136 379394 375148
rect 423950 375136 423956 375148
rect 379388 375108 423956 375136
rect 379388 375096 379394 375108
rect 423950 375096 423956 375108
rect 424008 375096 424014 375148
rect 106458 375028 106464 375080
rect 106516 375068 106522 375080
rect 218054 375068 218060 375080
rect 106516 375040 218060 375068
rect 106516 375028 106522 375040
rect 218054 375028 218060 375040
rect 218112 375028 218118 375080
rect 375558 375028 375564 375080
rect 375616 375068 375622 375080
rect 376570 375068 376576 375080
rect 375616 375040 376576 375068
rect 375616 375028 375622 375040
rect 376570 375028 376576 375040
rect 376628 375068 376634 375080
rect 405366 375068 405372 375080
rect 376628 375040 405372 375068
rect 376628 375028 376634 375040
rect 405366 375028 405372 375040
rect 405424 375028 405430 375080
rect 368382 374960 368388 375012
rect 368440 375000 368446 375012
rect 375742 375000 375748 375012
rect 368440 374972 375748 375000
rect 368440 374960 368446 374972
rect 375742 374960 375748 374972
rect 375800 375000 375806 375012
rect 416958 375000 416964 375012
rect 375800 374972 416964 375000
rect 375800 374960 375806 374972
rect 416958 374960 416964 374972
rect 417016 374960 417022 375012
rect 362770 374892 362776 374944
rect 362828 374932 362834 374944
rect 377122 374932 377128 374944
rect 362828 374904 377128 374932
rect 362828 374892 362834 374904
rect 377122 374892 377128 374904
rect 377180 374932 377186 374944
rect 418154 374932 418160 374944
rect 377180 374904 418160 374932
rect 377180 374892 377186 374904
rect 418154 374892 418160 374904
rect 418212 374892 418218 374944
rect 358722 374824 358728 374876
rect 358780 374864 358786 374876
rect 376478 374864 376484 374876
rect 358780 374836 376484 374864
rect 358780 374824 358786 374836
rect 376478 374824 376484 374836
rect 376536 374864 376542 374876
rect 418338 374864 418344 374876
rect 376536 374836 418344 374864
rect 376536 374824 376542 374836
rect 418338 374824 418344 374836
rect 418396 374824 418402 374876
rect 207014 374756 207020 374808
rect 207072 374796 207078 374808
rect 208118 374796 208124 374808
rect 207072 374768 208124 374796
rect 207072 374756 207078 374768
rect 208118 374756 208124 374768
rect 208176 374796 208182 374808
rect 217870 374796 217876 374808
rect 208176 374768 217876 374796
rect 208176 374756 208182 374768
rect 217870 374756 217876 374768
rect 217928 374796 217934 374808
rect 217928 374768 219434 374796
rect 217928 374756 217934 374768
rect 102962 374688 102968 374740
rect 103020 374728 103026 374740
rect 215110 374728 215116 374740
rect 103020 374700 215116 374728
rect 103020 374688 103026 374700
rect 215110 374688 215116 374700
rect 215168 374688 215174 374740
rect 219406 374728 219434 374768
rect 357158 374756 357164 374808
rect 357216 374796 357222 374808
rect 375558 374796 375564 374808
rect 357216 374768 375564 374796
rect 357216 374756 357222 374768
rect 375558 374756 375564 374768
rect 375616 374756 375622 374808
rect 378134 374796 378140 374808
rect 376496 374768 378140 374796
rect 267550 374728 267556 374740
rect 219406 374700 267556 374728
rect 267550 374688 267556 374700
rect 267608 374688 267614 374740
rect 371694 374688 371700 374740
rect 371752 374728 371758 374740
rect 376496 374728 376524 374768
rect 378134 374756 378140 374768
rect 378192 374796 378198 374808
rect 426434 374796 426440 374808
rect 378192 374768 426440 374796
rect 378192 374756 378198 374768
rect 426434 374756 426440 374768
rect 426492 374756 426498 374808
rect 429378 374728 429384 374740
rect 371752 374700 376524 374728
rect 376680 374700 429384 374728
rect 371752 374688 371758 374700
rect 183462 374620 183468 374672
rect 183520 374660 183526 374672
rect 197354 374660 197360 374672
rect 183520 374632 197360 374660
rect 183520 374620 183526 374632
rect 197354 374620 197360 374632
rect 197412 374660 197418 374672
rect 342254 374660 342260 374672
rect 197412 374632 342260 374660
rect 197412 374620 197418 374632
rect 342254 374620 342260 374632
rect 342312 374620 342318 374672
rect 370222 374620 370228 374672
rect 370280 374660 370286 374672
rect 372430 374660 372436 374672
rect 370280 374632 372436 374660
rect 370280 374620 370286 374632
rect 372430 374620 372436 374632
rect 372488 374620 372494 374672
rect 372448 374592 372476 374620
rect 376680 374592 376708 374700
rect 429378 374688 429384 374700
rect 429436 374688 429442 374740
rect 437750 374660 437756 374672
rect 372448 374564 376708 374592
rect 379486 374632 437756 374660
rect 370038 374484 370044 374536
rect 370096 374524 370102 374536
rect 370406 374524 370412 374536
rect 370096 374496 370412 374524
rect 370096 374484 370102 374496
rect 370406 374484 370412 374496
rect 370464 374524 370470 374536
rect 379486 374524 379514 374632
rect 437750 374620 437756 374632
rect 437808 374620 437814 374672
rect 370464 374496 379514 374524
rect 370464 374484 370470 374496
rect 199378 371832 199384 371884
rect 199436 371872 199442 371884
rect 199930 371872 199936 371884
rect 199436 371844 199936 371872
rect 199436 371832 199442 371844
rect 199930 371832 199936 371844
rect 199988 371872 199994 371884
rect 359182 371872 359188 371884
rect 199988 371844 359188 371872
rect 199988 371832 199994 371844
rect 359182 371832 359188 371844
rect 359240 371832 359246 371884
rect 359182 371220 359188 371272
rect 359240 371260 359246 371272
rect 359458 371260 359464 371272
rect 359240 371232 359464 371260
rect 359240 371220 359246 371232
rect 359458 371220 359464 371232
rect 359516 371220 359522 371272
rect 199470 370472 199476 370524
rect 199528 370512 199534 370524
rect 359090 370512 359096 370524
rect 199528 370484 359096 370512
rect 199528 370472 199534 370484
rect 359090 370472 359096 370484
rect 359148 370472 359154 370524
rect 359826 370472 359832 370524
rect 359884 370512 359890 370524
rect 518986 370512 518992 370524
rect 359884 370484 518992 370512
rect 359884 370472 359890 370484
rect 518986 370472 518992 370484
rect 519044 370472 519050 370524
rect 199654 369112 199660 369164
rect 199712 369152 199718 369164
rect 199838 369152 199844 369164
rect 199712 369124 199844 369152
rect 199712 369112 199718 369124
rect 199838 369112 199844 369124
rect 199896 369152 199902 369164
rect 359090 369152 359096 369164
rect 199896 369124 359096 369152
rect 199896 369112 199902 369124
rect 359090 369112 359096 369124
rect 359148 369152 359154 369164
rect 359826 369152 359832 369164
rect 359148 369124 359832 369152
rect 359148 369112 359154 369124
rect 359826 369112 359832 369124
rect 359884 369112 359890 369164
rect 199562 366324 199568 366376
rect 199620 366364 199626 366376
rect 358998 366364 359004 366376
rect 199620 366336 359004 366364
rect 199620 366324 199626 366336
rect 358998 366324 359004 366336
rect 359056 366364 359062 366376
rect 519262 366364 519268 366376
rect 359056 366336 519268 366364
rect 359056 366324 359062 366336
rect 519262 366324 519268 366336
rect 519320 366364 519326 366376
rect 519630 366364 519636 366376
rect 519320 366336 519636 366364
rect 519320 366324 519326 366336
rect 519630 366324 519636 366336
rect 519688 366324 519694 366376
rect 359182 364964 359188 365016
rect 359240 365004 359246 365016
rect 359550 365004 359556 365016
rect 359240 364976 359556 365004
rect 359240 364964 359246 364976
rect 359550 364964 359556 364976
rect 359608 365004 359614 365016
rect 518894 365004 518900 365016
rect 359608 364976 518900 365004
rect 359608 364964 359614 364976
rect 518894 364964 518900 364976
rect 518952 365004 518958 365016
rect 519078 365004 519084 365016
rect 518952 364976 519084 365004
rect 518952 364964 518958 364976
rect 519078 364964 519084 364976
rect 519136 364964 519142 365016
rect 359458 363604 359464 363656
rect 359516 363644 359522 363656
rect 519170 363644 519176 363656
rect 359516 363616 519176 363644
rect 359516 363604 359522 363616
rect 519170 363604 519176 363616
rect 519228 363604 519234 363656
rect 199746 362176 199752 362228
rect 199804 362216 199810 362228
rect 358906 362216 358912 362228
rect 199804 362188 358912 362216
rect 199804 362176 199810 362188
rect 358906 362176 358912 362188
rect 358964 362216 358970 362228
rect 359182 362216 359188 362228
rect 358964 362188 359188 362216
rect 358964 362176 358970 362188
rect 359182 362176 359188 362188
rect 359240 362216 359246 362228
rect 519446 362216 519452 362228
rect 359240 362188 519452 362216
rect 359240 362176 359246 362188
rect 519446 362176 519452 362188
rect 519504 362176 519510 362228
rect 202598 360204 202604 360256
rect 202656 360244 202662 360256
rect 206278 360244 206284 360256
rect 202656 360216 206284 360244
rect 202656 360204 202662 360216
rect 206278 360204 206284 360216
rect 206336 360204 206342 360256
rect 500770 359660 500776 359712
rect 500828 359700 500834 359712
rect 518066 359700 518072 359712
rect 500828 359672 518072 359700
rect 500828 359660 500834 359672
rect 518066 359660 518072 359672
rect 518124 359660 518130 359712
rect 197446 359524 197452 359576
rect 197504 359564 197510 359576
rect 208578 359564 208584 359576
rect 197504 359536 208584 359564
rect 197504 359524 197510 359536
rect 208578 359524 208584 359536
rect 208636 359524 208642 359576
rect 339862 359524 339868 359576
rect 339920 359564 339926 359576
rect 356974 359564 356980 359576
rect 339920 359536 356980 359564
rect 339920 359524 339926 359536
rect 356974 359524 356980 359536
rect 357032 359564 357038 359576
rect 357158 359564 357164 359576
rect 357032 359536 357164 359564
rect 357032 359524 357038 359536
rect 357158 359524 357164 359536
rect 357216 359524 357222 359576
rect 498930 359524 498936 359576
rect 498988 359564 498994 359576
rect 517974 359564 517980 359576
rect 498988 359536 517980 359564
rect 498988 359524 498994 359536
rect 517974 359524 517980 359536
rect 518032 359524 518038 359576
rect 190914 359456 190920 359508
rect 190972 359496 190978 359508
rect 201494 359496 201500 359508
rect 190972 359468 201500 359496
rect 190972 359456 190978 359468
rect 201494 359456 201500 359468
rect 201552 359496 201558 359508
rect 202598 359496 202604 359508
rect 201552 359468 202604 359496
rect 201552 359456 201558 359468
rect 202598 359456 202604 359468
rect 202656 359456 202662 359508
rect 351730 359456 351736 359508
rect 351788 359496 351794 359508
rect 358078 359496 358084 359508
rect 351788 359468 358084 359496
rect 351788 359456 351794 359468
rect 358078 359456 358084 359468
rect 358136 359456 358142 359508
rect 360194 359252 360200 359304
rect 360252 359292 360258 359304
rect 362954 359292 362960 359304
rect 360252 359264 362960 359292
rect 360252 359252 360258 359264
rect 362954 359252 362960 359264
rect 363012 359252 363018 359304
rect 179690 358844 179696 358896
rect 179748 358884 179754 358896
rect 179748 358856 197584 358884
rect 179748 358844 179754 358856
rect 178586 358776 178592 358828
rect 178644 358816 178650 358828
rect 197446 358816 197452 358828
rect 178644 358788 197452 358816
rect 178644 358776 178650 358788
rect 197446 358776 197452 358788
rect 197504 358776 197510 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 18598 358748 18604 358760
rect 3384 358720 18604 358748
rect 3384 358708 3390 358720
rect 18598 358708 18604 358720
rect 18656 358708 18662 358760
rect 55950 358708 55956 358760
rect 56008 358748 56014 358760
rect 59446 358748 59452 358760
rect 56008 358720 59452 358748
rect 56008 358708 56014 358720
rect 59446 358708 59452 358720
rect 59504 358708 59510 358760
rect 197556 358748 197584 358856
rect 342254 358844 342260 358896
rect 342312 358884 342318 358896
rect 343542 358884 343548 358896
rect 342312 358856 343548 358884
rect 342312 358844 342318 358856
rect 343542 358844 343548 358856
rect 343600 358884 343606 358896
rect 358538 358884 358544 358896
rect 343600 358856 358544 358884
rect 343600 358844 343606 358856
rect 358538 358844 358544 358856
rect 358596 358844 358602 358896
rect 338482 358776 338488 358828
rect 338540 358816 338546 358828
rect 360194 358816 360200 358828
rect 338540 358788 360200 358816
rect 338540 358776 338546 358788
rect 360194 358776 360200 358788
rect 360252 358776 360258 358828
rect 510890 358776 510896 358828
rect 510948 358816 510954 358828
rect 517514 358816 517520 358828
rect 510948 358788 517520 358816
rect 510948 358776 510954 358788
rect 517514 358776 517520 358788
rect 517572 358776 517578 358828
rect 198090 358748 198096 358760
rect 197556 358720 198096 358748
rect 198090 358708 198096 358720
rect 198148 358748 198154 358760
rect 203886 358748 203892 358760
rect 198148 358720 203892 358748
rect 198148 358708 198154 358720
rect 203886 358708 203892 358720
rect 203944 358708 203950 358760
rect 218514 358708 218520 358760
rect 218572 358748 218578 358760
rect 221366 358748 221372 358760
rect 218572 358720 221372 358748
rect 218572 358708 218578 358720
rect 221366 358708 221372 358720
rect 221424 358708 221430 358760
rect 379422 358708 379428 358760
rect 379480 358748 379486 358760
rect 380986 358748 380992 358760
rect 379480 358720 380992 358748
rect 379480 358708 379486 358720
rect 380986 358708 380992 358720
rect 381044 358708 381050 358760
rect 219250 358640 219256 358692
rect 219308 358680 219314 358692
rect 220906 358680 220912 358692
rect 219308 358652 220912 358680
rect 219308 358640 219314 358652
rect 220906 358640 220912 358652
rect 220964 358640 220970 358692
rect 375282 358640 375288 358692
rect 375340 358680 375346 358692
rect 381078 358680 381084 358692
rect 375340 358652 381084 358680
rect 375340 358640 375346 358652
rect 381078 358640 381084 358652
rect 381136 358640 381142 358692
rect 217042 358572 217048 358624
rect 217100 358612 217106 358624
rect 220814 358612 220820 358624
rect 217100 358584 220820 358612
rect 217100 358572 217106 358584
rect 220814 358572 220820 358584
rect 220872 358572 220878 358624
rect 214374 358504 214380 358556
rect 214432 358544 214438 358556
rect 220998 358544 221004 358556
rect 214432 358516 221004 358544
rect 214432 358504 214438 358516
rect 220998 358504 221004 358516
rect 221056 358504 221062 358556
rect 219158 358232 219164 358284
rect 219216 358272 219222 358284
rect 221090 358272 221096 358284
rect 219216 358244 221096 358272
rect 219216 358232 219222 358244
rect 221090 358232 221096 358244
rect 221148 358232 221154 358284
rect 215662 358096 215668 358148
rect 215720 358136 215726 358148
rect 221182 358136 221188 358148
rect 215720 358108 221188 358136
rect 215720 358096 215726 358108
rect 221182 358096 221188 358108
rect 221240 358096 221246 358148
rect 182818 358028 182824 358080
rect 182876 358068 182882 358080
rect 201586 358068 201592 358080
rect 182876 358040 201592 358068
rect 182876 358028 182882 358040
rect 201586 358028 201592 358040
rect 201644 358068 201650 358080
rect 342254 358068 342260 358080
rect 201644 358040 342260 358068
rect 201644 358028 201650 358040
rect 342254 358028 342260 358040
rect 342312 358028 342318 358080
rect 377030 357960 377036 358012
rect 377088 358000 377094 358012
rect 381262 358000 381268 358012
rect 377088 357972 381268 358000
rect 377088 357960 377094 357972
rect 381262 357960 381268 357972
rect 381320 357960 381326 358012
rect 57146 357824 57152 357876
rect 57204 357864 57210 357876
rect 59354 357864 59360 357876
rect 57204 357836 59360 357864
rect 57204 357824 57210 357836
rect 59354 357824 59360 357836
rect 59412 357824 59418 357876
rect 378686 357824 378692 357876
rect 378744 357864 378750 357876
rect 380894 357864 380900 357876
rect 378744 357836 380900 357864
rect 378744 357824 378750 357836
rect 380894 357824 380900 357836
rect 380952 357824 380958 357876
rect 215846 357484 215852 357536
rect 215904 357524 215910 357536
rect 221274 357524 221280 357536
rect 215904 357496 221280 357524
rect 215904 357484 215910 357496
rect 221274 357484 221280 357496
rect 221332 357484 221338 357536
rect 375834 357484 375840 357536
rect 375892 357524 375898 357536
rect 381170 357524 381176 357536
rect 375892 357496 381176 357524
rect 375892 357484 375898 357496
rect 381170 357484 381176 357496
rect 381228 357484 381234 357536
rect 58618 357348 58624 357400
rect 58676 357388 58682 357400
rect 60734 357388 60740 357400
rect 58676 357360 60740 357388
rect 58676 357348 58682 357360
rect 60734 357348 60740 357360
rect 60792 357348 60798 357400
rect 55122 303900 55128 303952
rect 55180 303940 55186 303952
rect 56594 303940 56600 303952
rect 55180 303912 56600 303940
rect 55180 303900 55186 303912
rect 56594 303900 56600 303912
rect 56652 303900 56658 303952
rect 46290 303560 46296 303612
rect 46348 303600 46354 303612
rect 57330 303600 57336 303612
rect 46348 303572 57336 303600
rect 46348 303560 46354 303572
rect 57330 303560 57336 303572
rect 57388 303600 57394 303612
rect 57606 303600 57612 303612
rect 57388 303572 57612 303600
rect 57388 303560 57394 303572
rect 57606 303560 57612 303572
rect 57664 303560 57670 303612
rect 46382 300772 46388 300824
rect 46440 300812 46446 300824
rect 56962 300812 56968 300824
rect 46440 300784 56968 300812
rect 46440 300772 46446 300784
rect 56962 300772 56968 300784
rect 57020 300812 57026 300824
rect 57422 300812 57428 300824
rect 57020 300784 57428 300812
rect 57020 300772 57026 300784
rect 57422 300772 57428 300784
rect 57480 300772 57486 300824
rect 520182 288396 520188 288448
rect 520240 288436 520246 288448
rect 580258 288436 580264 288448
rect 520240 288408 580264 288436
rect 520240 288396 520246 288408
rect 580258 288396 580264 288408
rect 580316 288396 580322 288448
rect 518986 287036 518992 287088
rect 519044 287076 519050 287088
rect 519446 287076 519452 287088
rect 519044 287048 519452 287076
rect 519044 287036 519050 287048
rect 519446 287036 519452 287048
rect 519504 287076 519510 287088
rect 580350 287076 580356 287088
rect 519504 287048 580356 287076
rect 519504 287036 519510 287048
rect 580350 287036 580356 287048
rect 580408 287036 580414 287088
rect 200942 284248 200948 284300
rect 201000 284288 201006 284300
rect 216674 284288 216680 284300
rect 201000 284260 216680 284288
rect 201000 284248 201006 284260
rect 216674 284248 216680 284260
rect 216732 284248 216738 284300
rect 361206 284248 361212 284300
rect 361264 284288 361270 284300
rect 376938 284288 376944 284300
rect 361264 284260 376944 284288
rect 361264 284248 361270 284260
rect 376938 284248 376944 284260
rect 376996 284248 377002 284300
rect 201494 282820 201500 282872
rect 201552 282860 201558 282872
rect 216674 282860 216680 282872
rect 201552 282832 216680 282860
rect 201552 282820 201558 282832
rect 216674 282820 216680 282832
rect 216732 282820 216738 282872
rect 368198 282820 368204 282872
rect 368256 282860 368262 282872
rect 376754 282860 376760 282872
rect 368256 282832 376760 282860
rect 368256 282820 368262 282832
rect 376754 282820 376760 282832
rect 376812 282820 376818 282872
rect 203794 282752 203800 282804
rect 203852 282792 203858 282804
rect 216766 282792 216772 282804
rect 203852 282764 216772 282792
rect 203852 282752 203858 282764
rect 216766 282752 216772 282764
rect 216824 282752 216830 282804
rect 55122 282208 55128 282260
rect 55180 282248 55186 282260
rect 58710 282248 58716 282260
rect 55180 282220 58716 282248
rect 55180 282208 55186 282220
rect 58710 282208 58716 282220
rect 58768 282208 58774 282260
rect 51626 282140 51632 282192
rect 51684 282180 51690 282192
rect 58526 282180 58532 282192
rect 51684 282152 58532 282180
rect 51684 282140 51690 282152
rect 58526 282140 58532 282152
rect 58584 282140 58590 282192
rect 358078 282140 358084 282192
rect 358136 282180 358142 282192
rect 376938 282180 376944 282192
rect 358136 282152 376944 282180
rect 358136 282140 358142 282152
rect 376938 282140 376944 282152
rect 376996 282140 377002 282192
rect 44082 281460 44088 281512
rect 44140 281500 44146 281512
rect 57238 281500 57244 281512
rect 44140 281472 57244 281500
rect 44140 281460 44146 281472
rect 57238 281460 57244 281472
rect 57296 281500 57302 281512
rect 57514 281500 57520 281512
rect 57296 281472 57520 281500
rect 57296 281460 57302 281472
rect 57514 281460 57520 281472
rect 57572 281460 57578 281512
rect 374454 274728 374460 274780
rect 374512 274768 374518 274780
rect 375006 274768 375012 274780
rect 374512 274740 375012 274768
rect 374512 274728 374518 274740
rect 375006 274728 375012 274740
rect 375064 274728 375070 274780
rect 212902 274660 212908 274712
rect 212960 274700 212966 274712
rect 215386 274700 215392 274712
rect 212960 274672 215392 274700
rect 212960 274660 212966 274672
rect 215386 274660 215392 274672
rect 215444 274660 215450 274712
rect 219342 273572 219348 273624
rect 219400 273612 219406 273624
rect 219894 273612 219900 273624
rect 219400 273584 219900 273612
rect 219400 273572 219406 273584
rect 219894 273572 219900 273584
rect 219952 273612 219958 273624
rect 266354 273612 266360 273624
rect 219952 273584 266360 273612
rect 219952 273572 219958 273584
rect 266354 273572 266360 273584
rect 266412 273572 266418 273624
rect 55858 273504 55864 273556
rect 55916 273544 55922 273556
rect 110966 273544 110972 273556
rect 55916 273516 110972 273544
rect 55916 273504 55922 273516
rect 110966 273504 110972 273516
rect 111024 273504 111030 273556
rect 200850 273504 200856 273556
rect 200908 273544 200914 273556
rect 250714 273544 250720 273556
rect 200908 273516 250720 273544
rect 200908 273504 200914 273516
rect 250714 273504 250720 273516
rect 250772 273504 250778 273556
rect 44818 273436 44824 273488
rect 44876 273476 44882 273488
rect 133414 273476 133420 273488
rect 44876 273448 133420 273476
rect 44876 273436 44882 273448
rect 133414 273436 133420 273448
rect 133472 273436 133478 273488
rect 215386 273436 215392 273488
rect 215444 273476 215450 273488
rect 273346 273476 273352 273488
rect 215444 273448 273352 273476
rect 215444 273436 215450 273448
rect 273346 273436 273352 273448
rect 273404 273436 273410 273488
rect 370314 273436 370320 273488
rect 370372 273476 370378 273488
rect 379330 273476 379336 273488
rect 370372 273448 379336 273476
rect 370372 273436 370378 273448
rect 379330 273436 379336 273448
rect 379388 273436 379394 273488
rect 45186 273368 45192 273420
rect 45244 273408 45250 273420
rect 135898 273408 135904 273420
rect 45244 273380 135904 273408
rect 45244 273368 45250 273380
rect 135898 273368 135904 273380
rect 135956 273368 135962 273420
rect 213454 273368 213460 273420
rect 213512 273408 213518 273420
rect 215018 273408 215024 273420
rect 213512 273380 215024 273408
rect 213512 273368 213518 273380
rect 215018 273368 215024 273380
rect 215076 273408 215082 273420
rect 275738 273408 275744 273420
rect 215076 273380 275744 273408
rect 215076 273368 215082 273380
rect 275738 273368 275744 273380
rect 275796 273368 275802 273420
rect 369026 273368 369032 273420
rect 369084 273408 369090 273420
rect 378134 273408 378140 273420
rect 369084 273380 378140 273408
rect 369084 273368 369090 273380
rect 378134 273368 378140 273380
rect 378192 273408 378198 273420
rect 378594 273408 378600 273420
rect 378192 273380 378600 273408
rect 378192 273368 378198 273380
rect 378594 273368 378600 273380
rect 378652 273368 378658 273420
rect 45094 273300 45100 273352
rect 45152 273340 45158 273352
rect 138474 273340 138480 273352
rect 45152 273312 138480 273340
rect 45152 273300 45158 273312
rect 138474 273300 138480 273312
rect 138532 273300 138538 273352
rect 215754 273300 215760 273352
rect 215812 273340 215818 273352
rect 278038 273340 278044 273352
rect 215812 273312 278044 273340
rect 215812 273300 215818 273312
rect 278038 273300 278044 273312
rect 278096 273300 278102 273352
rect 362678 273300 362684 273352
rect 362736 273340 362742 273352
rect 421098 273340 421104 273352
rect 362736 273312 421104 273340
rect 362736 273300 362742 273312
rect 421098 273300 421104 273312
rect 421156 273300 421162 273352
rect 45002 273232 45008 273284
rect 45060 273272 45066 273284
rect 140866 273272 140872 273284
rect 45060 273244 140872 273272
rect 45060 273232 45066 273244
rect 140866 273232 140872 273244
rect 140924 273232 140930 273284
rect 205266 273232 205272 273284
rect 205324 273272 205330 273284
rect 283466 273272 283472 273284
rect 205324 273244 283472 273272
rect 205324 273232 205330 273244
rect 283466 273232 283472 273244
rect 283524 273232 283530 273284
rect 369394 273232 369400 273284
rect 369452 273272 369458 273284
rect 450998 273272 451004 273284
rect 369452 273244 451004 273272
rect 369452 273232 369458 273244
rect 450998 273232 451004 273244
rect 451056 273232 451062 273284
rect 371142 273164 371148 273216
rect 371200 273204 371206 273216
rect 375190 273204 375196 273216
rect 371200 273176 375196 273204
rect 371200 273164 371206 273176
rect 375190 273164 375196 273176
rect 375248 273164 375254 273216
rect 379330 273164 379336 273216
rect 379388 273204 379394 273216
rect 423766 273204 423772 273216
rect 379388 273176 423772 273204
rect 379388 273164 379394 273176
rect 423766 273164 423772 273176
rect 423824 273164 423830 273216
rect 53834 273096 53840 273148
rect 53892 273136 53898 273148
rect 100754 273136 100760 273148
rect 53892 273108 100760 273136
rect 53892 273096 53898 273108
rect 100754 273096 100760 273108
rect 100812 273096 100818 273148
rect 378594 273096 378600 273148
rect 378652 273136 378658 273148
rect 426434 273136 426440 273148
rect 378652 273108 426440 273136
rect 378652 273096 378658 273108
rect 426434 273096 426440 273108
rect 426492 273096 426498 273148
rect 365438 273028 365444 273080
rect 365496 273068 365502 273080
rect 423398 273068 423404 273080
rect 365496 273040 423404 273068
rect 365496 273028 365502 273040
rect 423398 273028 423404 273040
rect 423456 273028 423462 273080
rect 60826 273000 60832 273012
rect 45526 272972 60832 273000
rect 42518 272824 42524 272876
rect 42576 272864 42582 272876
rect 45526 272864 45554 272972
rect 60826 272960 60832 272972
rect 60884 272960 60890 273012
rect 210326 272960 210332 273012
rect 210384 273000 210390 273012
rect 288158 273000 288164 273012
rect 210384 272972 288164 273000
rect 210384 272960 210390 272972
rect 288158 272960 288164 272972
rect 288216 272960 288222 273012
rect 372338 272960 372344 273012
rect 372396 273000 372402 273012
rect 373166 273000 373172 273012
rect 372396 272972 373172 273000
rect 372396 272960 372402 272972
rect 373166 272960 373172 272972
rect 373224 273000 373230 273012
rect 431126 273000 431132 273012
rect 373224 272972 431132 273000
rect 373224 272960 373230 272972
rect 431126 272960 431132 272972
rect 431184 272960 431190 273012
rect 58618 272892 58624 272944
rect 58676 272932 58682 272944
rect 61102 272932 61108 272944
rect 58676 272904 61108 272932
rect 58676 272892 58682 272904
rect 61102 272892 61108 272904
rect 61160 272932 61166 272944
rect 61470 272932 61476 272944
rect 61160 272904 61476 272932
rect 61160 272892 61166 272904
rect 61470 272892 61476 272904
rect 61528 272892 61534 272944
rect 206738 272892 206744 272944
rect 206796 272932 206802 272944
rect 285950 272932 285956 272944
rect 206796 272904 285956 272932
rect 206796 272892 206802 272904
rect 285950 272892 285956 272904
rect 286008 272892 286014 272944
rect 358446 272892 358452 272944
rect 358504 272932 358510 272944
rect 425974 272932 425980 272944
rect 358504 272904 425980 272932
rect 358504 272892 358510 272904
rect 425974 272892 425980 272904
rect 426032 272892 426038 272944
rect 42576 272836 45554 272864
rect 42576 272824 42582 272836
rect 59630 272824 59636 272876
rect 59688 272864 59694 272876
rect 60734 272864 60740 272876
rect 59688 272836 60740 272864
rect 59688 272824 59694 272836
rect 60734 272824 60740 272836
rect 60792 272864 60798 272876
rect 61746 272864 61752 272876
rect 60792 272836 61752 272864
rect 60792 272824 60798 272836
rect 61746 272824 61752 272836
rect 61804 272824 61810 272876
rect 209314 272824 209320 272876
rect 209372 272864 209378 272876
rect 290918 272864 290924 272876
rect 209372 272836 290924 272864
rect 209372 272824 209378 272836
rect 290918 272824 290924 272836
rect 290976 272824 290982 272876
rect 356882 272824 356888 272876
rect 356940 272864 356946 272876
rect 428182 272864 428188 272876
rect 356940 272836 428188 272864
rect 356940 272824 356946 272836
rect 428182 272824 428188 272836
rect 428240 272824 428246 272876
rect 50430 272756 50436 272808
rect 50488 272796 50494 272808
rect 90726 272796 90732 272808
rect 50488 272768 90732 272796
rect 50488 272756 50494 272768
rect 90726 272756 90732 272768
rect 90784 272756 90790 272808
rect 210878 272756 210884 272808
rect 210936 272796 210942 272808
rect 300854 272796 300860 272808
rect 210936 272768 300860 272796
rect 210936 272756 210942 272768
rect 300854 272756 300860 272768
rect 300912 272756 300918 272808
rect 370958 272756 370964 272808
rect 371016 272796 371022 272808
rect 468478 272796 468484 272808
rect 371016 272768 468484 272796
rect 371016 272756 371022 272768
rect 468478 272756 468484 272768
rect 468536 272756 468542 272808
rect 47854 272688 47860 272740
rect 47912 272728 47918 272740
rect 93670 272728 93676 272740
rect 47912 272700 93676 272728
rect 47912 272688 47918 272700
rect 93670 272688 93676 272700
rect 93728 272688 93734 272740
rect 202506 272688 202512 272740
rect 202564 272728 202570 272740
rect 293310 272728 293316 272740
rect 202564 272700 293316 272728
rect 202564 272688 202570 272700
rect 293310 272688 293316 272700
rect 293368 272688 293374 272740
rect 376294 272688 376300 272740
rect 376352 272728 376358 272740
rect 473446 272728 473452 272740
rect 376352 272700 473452 272728
rect 376352 272688 376358 272700
rect 473446 272688 473452 272700
rect 473504 272688 473510 272740
rect 49234 272620 49240 272672
rect 49292 272660 49298 272672
rect 95878 272660 95884 272672
rect 49292 272632 95884 272660
rect 49292 272620 49298 272632
rect 95878 272620 95884 272632
rect 95936 272620 95942 272672
rect 205174 272620 205180 272672
rect 205232 272660 205238 272672
rect 298462 272660 298468 272672
rect 205232 272632 298468 272660
rect 205232 272620 205238 272632
rect 298462 272620 298468 272632
rect 298520 272620 298526 272672
rect 364058 272620 364064 272672
rect 364116 272660 364122 272672
rect 470870 272660 470876 272672
rect 364116 272632 470876 272660
rect 364116 272620 364122 272632
rect 470870 272620 470876 272632
rect 470928 272620 470934 272672
rect 51902 272552 51908 272604
rect 51960 272592 51966 272604
rect 98454 272592 98460 272604
rect 51960 272564 98460 272592
rect 51960 272552 51966 272564
rect 98454 272552 98460 272564
rect 98512 272552 98518 272604
rect 207842 272552 207848 272604
rect 207900 272592 207906 272604
rect 305822 272592 305828 272604
rect 207900 272564 305828 272592
rect 207900 272552 207906 272564
rect 305822 272552 305828 272564
rect 305880 272552 305886 272604
rect 366818 272552 366824 272604
rect 366876 272592 366882 272604
rect 475838 272592 475844 272604
rect 366876 272564 475844 272592
rect 366876 272552 366882 272564
rect 475838 272552 475844 272564
rect 475896 272552 475902 272604
rect 45278 272484 45284 272536
rect 45336 272524 45342 272536
rect 143534 272524 143540 272536
rect 45336 272496 143540 272524
rect 45336 272484 45342 272496
rect 143534 272484 143540 272496
rect 143592 272484 143598 272536
rect 208210 272484 208216 272536
rect 208268 272524 208274 272536
rect 210878 272524 210884 272536
rect 208268 272496 210884 272524
rect 208268 272484 208274 272496
rect 210878 272484 210884 272496
rect 210936 272484 210942 272536
rect 212258 272484 212264 272536
rect 212316 272524 212322 272536
rect 320910 272524 320916 272536
rect 212316 272496 320916 272524
rect 212316 272484 212322 272496
rect 320910 272484 320916 272496
rect 320968 272484 320974 272536
rect 368106 272484 368112 272536
rect 368164 272524 368170 272536
rect 478414 272524 478420 272536
rect 368164 272496 478420 272524
rect 368164 272484 368170 272496
rect 478414 272484 478420 272496
rect 478472 272484 478478 272536
rect 46658 272416 46664 272468
rect 46716 272456 46722 272468
rect 47486 272456 47492 272468
rect 46716 272428 47492 272456
rect 46716 272416 46722 272428
rect 47486 272416 47492 272428
rect 47544 272456 47550 272468
rect 47544 272428 55214 272456
rect 47544 272416 47550 272428
rect 46566 272348 46572 272400
rect 46624 272388 46630 272400
rect 47670 272388 47676 272400
rect 46624 272360 47676 272388
rect 46624 272348 46630 272360
rect 47670 272348 47676 272360
rect 47728 272348 47734 272400
rect 55186 272388 55214 272428
rect 58526 272416 58532 272468
rect 58584 272456 58590 272468
rect 59722 272456 59728 272468
rect 58584 272428 59728 272456
rect 58584 272416 58590 272428
rect 59722 272416 59728 272428
rect 59780 272456 59786 272468
rect 99374 272456 99380 272468
rect 59780 272428 99380 272456
rect 59780 272416 59786 272428
rect 99374 272416 99380 272428
rect 99432 272416 99438 272468
rect 374546 272416 374552 272468
rect 374604 272456 374610 272468
rect 396718 272456 396724 272468
rect 374604 272428 396724 272456
rect 374604 272416 374610 272428
rect 396718 272416 396724 272428
rect 396776 272416 396782 272468
rect 76006 272388 76012 272400
rect 55186 272360 76012 272388
rect 76006 272348 76012 272360
rect 76064 272348 76070 272400
rect 65334 272280 65340 272332
rect 65392 272320 65398 272332
rect 95970 272320 95976 272332
rect 65392 272292 95976 272320
rect 65392 272280 65398 272292
rect 95970 272280 95976 272292
rect 96028 272280 96034 272332
rect 67358 272212 67364 272264
rect 67416 272252 67422 272264
rect 96982 272252 96988 272264
rect 67416 272224 96988 272252
rect 67416 272212 67422 272224
rect 96982 272212 96988 272224
rect 97040 272212 97046 272264
rect 46750 272144 46756 272196
rect 46808 272184 46814 272196
rect 46934 272184 46940 272196
rect 46808 272156 46940 272184
rect 46808 272144 46814 272156
rect 46934 272144 46940 272156
rect 46992 272144 46998 272196
rect 60826 272144 60832 272196
rect 60884 272184 60890 272196
rect 94222 272184 94228 272196
rect 60884 272156 94228 272184
rect 60884 272144 60890 272156
rect 94222 272144 94228 272156
rect 94280 272144 94286 272196
rect 53926 272076 53932 272128
rect 53984 272116 53990 272128
rect 86954 272116 86960 272128
rect 53984 272088 86960 272116
rect 53984 272076 53990 272088
rect 86954 272076 86960 272088
rect 87012 272076 87018 272128
rect 49326 272008 49332 272060
rect 49384 272048 49390 272060
rect 82814 272048 82820 272060
rect 49384 272020 82820 272048
rect 49384 272008 49390 272020
rect 82814 272008 82820 272020
rect 82872 272008 82878 272060
rect 83458 272008 83464 272060
rect 83516 272048 83522 272060
rect 97994 272048 98000 272060
rect 83516 272020 98000 272048
rect 83516 272008 83522 272020
rect 97994 272008 98000 272020
rect 98052 272008 98058 272060
rect 47670 271940 47676 271992
rect 47728 271980 47734 271992
rect 75914 271980 75920 271992
rect 47728 271952 75920 271980
rect 47728 271940 47734 271952
rect 75914 271940 75920 271952
rect 75972 271940 75978 271992
rect 213730 271940 213736 271992
rect 213788 271980 213794 271992
rect 216214 271980 216220 271992
rect 213788 271952 216220 271980
rect 213788 271940 213794 271952
rect 216214 271940 216220 271952
rect 216272 271980 216278 271992
rect 235994 271980 236000 271992
rect 216272 271952 236000 271980
rect 216272 271940 216278 271952
rect 235994 271940 236000 271952
rect 236052 271940 236058 271992
rect 421558 271940 421564 271992
rect 421616 271980 421622 271992
rect 437934 271980 437940 271992
rect 421616 271952 437940 271980
rect 421616 271940 421622 271952
rect 437934 271940 437940 271952
rect 437992 271940 437998 271992
rect 98638 271872 98644 271924
rect 98696 271912 98702 271924
rect 100754 271912 100760 271924
rect 98696 271884 100760 271912
rect 98696 271872 98702 271884
rect 100754 271872 100760 271884
rect 100812 271872 100818 271924
rect 114462 271872 114468 271924
rect 114520 271912 114526 271924
rect 127618 271912 127624 271924
rect 114520 271884 127624 271912
rect 114520 271872 114526 271884
rect 127618 271872 127624 271884
rect 127676 271872 127682 271924
rect 210878 271872 210884 271924
rect 210936 271912 210942 271924
rect 268194 271912 268200 271924
rect 210936 271884 268200 271912
rect 210936 271872 210942 271884
rect 268194 271872 268200 271884
rect 268252 271872 268258 271924
rect 356974 271872 356980 271924
rect 357032 271912 357038 271924
rect 359366 271912 359372 271924
rect 357032 271884 359372 271912
rect 357032 271872 357038 271884
rect 359366 271872 359372 271884
rect 359424 271872 359430 271924
rect 360286 271912 360292 271924
rect 359476 271884 360292 271912
rect 43530 271804 43536 271856
rect 43588 271844 43594 271856
rect 129734 271844 129740 271856
rect 43588 271816 129740 271844
rect 43588 271804 43594 271816
rect 129734 271804 129740 271816
rect 129792 271804 129798 271856
rect 151354 271804 151360 271856
rect 151412 271844 151418 271856
rect 197998 271844 198004 271856
rect 151412 271816 198004 271844
rect 151412 271804 151418 271816
rect 197998 271804 198004 271816
rect 198056 271804 198062 271856
rect 213178 271804 213184 271856
rect 213236 271844 213242 271856
rect 313274 271844 313280 271856
rect 213236 271816 313280 271844
rect 213236 271804 213242 271816
rect 313274 271804 313280 271816
rect 313332 271804 313338 271856
rect 343542 271804 343548 271856
rect 343600 271844 343606 271856
rect 358538 271844 358544 271856
rect 343600 271816 358544 271844
rect 343600 271804 343606 271816
rect 358538 271804 358544 271816
rect 358596 271844 358602 271856
rect 359476 271844 359504 271884
rect 360286 271872 360292 271884
rect 360344 271872 360350 271924
rect 374454 271872 374460 271924
rect 374512 271912 374518 271924
rect 375190 271912 375196 271924
rect 374512 271884 375196 271912
rect 374512 271872 374518 271884
rect 375190 271872 375196 271884
rect 375248 271912 375254 271924
rect 402974 271912 402980 271924
rect 375248 271884 402980 271912
rect 375248 271872 375254 271884
rect 402974 271872 402980 271884
rect 403032 271872 403038 271924
rect 358596 271816 359504 271844
rect 358596 271804 358602 271816
rect 366726 271804 366732 271856
rect 366784 271844 366790 271856
rect 455782 271844 455788 271856
rect 366784 271816 455788 271844
rect 366784 271804 366790 271816
rect 455782 271804 455788 271816
rect 455840 271804 455846 271856
rect 42334 271736 42340 271788
rect 42392 271776 42398 271788
rect 123202 271776 123208 271788
rect 42392 271748 123208 271776
rect 42392 271736 42398 271748
rect 123202 271736 123208 271748
rect 123260 271736 123266 271788
rect 157242 271736 157248 271788
rect 157300 271776 157306 271788
rect 203058 271776 203064 271788
rect 157300 271748 203064 271776
rect 157300 271736 157306 271748
rect 203058 271736 203064 271748
rect 203116 271736 203122 271788
rect 212074 271736 212080 271788
rect 212132 271776 212138 271788
rect 307754 271776 307760 271788
rect 212132 271748 307760 271776
rect 212132 271736 212138 271748
rect 307754 271736 307760 271748
rect 307812 271736 307818 271788
rect 373534 271736 373540 271788
rect 373592 271776 373598 271788
rect 458174 271776 458180 271788
rect 373592 271748 458180 271776
rect 373592 271736 373598 271748
rect 458174 271736 458180 271748
rect 458232 271736 458238 271788
rect 42426 271668 42432 271720
rect 42484 271708 42490 271720
rect 53834 271708 53840 271720
rect 42484 271680 53840 271708
rect 42484 271668 42490 271680
rect 53834 271668 53840 271680
rect 53892 271708 53898 271720
rect 54386 271708 54392 271720
rect 53892 271680 54392 271708
rect 53892 271668 53898 271680
rect 54386 271668 54392 271680
rect 54444 271668 54450 271720
rect 57146 271668 57152 271720
rect 57204 271708 57210 271720
rect 128354 271708 128360 271720
rect 57204 271680 128360 271708
rect 57204 271668 57210 271680
rect 128354 271668 128360 271680
rect 128412 271668 128418 271720
rect 154482 271668 154488 271720
rect 154540 271708 154546 271720
rect 200298 271708 200304 271720
rect 154540 271680 200304 271708
rect 154540 271668 154546 271680
rect 200298 271668 200304 271680
rect 200356 271668 200362 271720
rect 200758 271668 200764 271720
rect 200816 271708 200822 271720
rect 268010 271708 268016 271720
rect 200816 271680 268016 271708
rect 200816 271668 200822 271680
rect 268010 271668 268016 271680
rect 268068 271668 268074 271720
rect 369486 271668 369492 271720
rect 369544 271708 369550 271720
rect 452654 271708 452660 271720
rect 369544 271680 452660 271708
rect 369544 271668 369550 271680
rect 452654 271668 452660 271680
rect 452712 271668 452718 271720
rect 46474 271600 46480 271652
rect 46532 271640 46538 271652
rect 53926 271640 53932 271652
rect 46532 271612 53932 271640
rect 46532 271600 46538 271612
rect 53926 271600 53932 271612
rect 53984 271600 53990 271652
rect 55950 271600 55956 271652
rect 56008 271640 56014 271652
rect 125594 271640 125600 271652
rect 56008 271612 125600 271640
rect 56008 271600 56014 271612
rect 125594 271600 125600 271612
rect 125652 271600 125658 271652
rect 158622 271600 158628 271652
rect 158680 271640 158686 271652
rect 201678 271640 201684 271652
rect 158680 271612 201684 271640
rect 158680 271600 158686 271612
rect 201678 271600 201684 271612
rect 201736 271600 201742 271652
rect 214834 271600 214840 271652
rect 214892 271640 214898 271652
rect 280154 271640 280160 271652
rect 214892 271612 280160 271640
rect 214892 271600 214898 271612
rect 280154 271600 280160 271612
rect 280212 271600 280218 271652
rect 365346 271600 365352 271652
rect 365404 271640 365410 271652
rect 445754 271640 445760 271652
rect 365404 271612 445760 271640
rect 365404 271600 365410 271612
rect 445754 271600 445760 271612
rect 445812 271600 445818 271652
rect 54570 271532 54576 271584
rect 54628 271572 54634 271584
rect 120074 271572 120080 271584
rect 54628 271544 120080 271572
rect 54628 271532 54634 271544
rect 120074 271532 120080 271544
rect 120132 271532 120138 271584
rect 161290 271532 161296 271584
rect 161348 271572 161354 271584
rect 197630 271572 197636 271584
rect 161348 271544 197636 271572
rect 161348 271532 161354 271544
rect 197630 271532 197636 271544
rect 197688 271532 197694 271584
rect 214926 271532 214932 271584
rect 214984 271572 214990 271584
rect 276014 271572 276020 271584
rect 214984 271544 276020 271572
rect 214984 271532 214990 271544
rect 276014 271532 276020 271544
rect 276072 271532 276078 271584
rect 372154 271532 372160 271584
rect 372212 271572 372218 271584
rect 447134 271572 447140 271584
rect 372212 271544 447140 271572
rect 372212 271532 372218 271544
rect 447134 271532 447140 271544
rect 447192 271532 447198 271584
rect 52914 271464 52920 271516
rect 52972 271504 52978 271516
rect 117314 271504 117320 271516
rect 52972 271476 117320 271504
rect 52972 271464 52978 271476
rect 117314 271464 117320 271476
rect 117372 271464 117378 271516
rect 164142 271464 164148 271516
rect 164200 271504 164206 271516
rect 197722 271504 197728 271516
rect 164200 271476 197728 271504
rect 164200 271464 164206 271476
rect 197722 271464 197728 271476
rect 197780 271464 197786 271516
rect 205082 271464 205088 271516
rect 205140 271504 205146 271516
rect 264974 271504 264980 271516
rect 205140 271476 264980 271504
rect 205140 271464 205146 271476
rect 264974 271464 264980 271476
rect 265032 271464 265038 271516
rect 363966 271464 363972 271516
rect 364024 271504 364030 271516
rect 437474 271504 437480 271516
rect 364024 271476 437480 271504
rect 364024 271464 364030 271476
rect 437474 271464 437480 271476
rect 437532 271464 437538 271516
rect 48130 271396 48136 271448
rect 48188 271436 48194 271448
rect 51902 271436 51908 271448
rect 48188 271408 51908 271436
rect 48188 271396 48194 271408
rect 51902 271396 51908 271408
rect 51960 271396 51966 271448
rect 53098 271396 53104 271448
rect 53156 271436 53162 271448
rect 115934 271436 115940 271448
rect 53156 271408 115940 271436
rect 53156 271396 53162 271408
rect 115934 271396 115940 271408
rect 115992 271396 115998 271448
rect 210786 271396 210792 271448
rect 210844 271436 210850 271448
rect 270494 271436 270500 271448
rect 210844 271408 270500 271436
rect 210844 271396 210850 271408
rect 270494 271396 270500 271408
rect 270552 271396 270558 271448
rect 361022 271396 361028 271448
rect 361080 271436 361086 271448
rect 433334 271436 433340 271448
rect 361080 271408 433340 271436
rect 361080 271396 361086 271408
rect 433334 271396 433340 271408
rect 433392 271396 433398 271448
rect 48038 271328 48044 271380
rect 48096 271368 48102 271380
rect 52454 271368 52460 271380
rect 48096 271340 52460 271368
rect 48096 271328 48102 271340
rect 52454 271328 52460 271340
rect 52512 271328 52518 271380
rect 53006 271328 53012 271380
rect 53064 271368 53070 271380
rect 113542 271368 113548 271380
rect 53064 271340 113548 271368
rect 53064 271328 53070 271340
rect 113542 271328 113548 271340
rect 113600 271328 113606 271380
rect 219066 271328 219072 271380
rect 219124 271368 219130 271380
rect 277670 271368 277676 271380
rect 219124 271340 277676 271368
rect 219124 271328 219130 271340
rect 277670 271328 277676 271340
rect 277728 271328 277734 271380
rect 368014 271328 368020 271380
rect 368072 271368 368078 271380
rect 440234 271368 440240 271380
rect 368072 271340 440240 271368
rect 368072 271328 368078 271340
rect 440234 271328 440240 271340
rect 440292 271328 440298 271380
rect 503622 271328 503628 271380
rect 503680 271368 503686 271380
rect 517606 271368 517612 271380
rect 503680 271340 517612 271368
rect 503680 271328 503686 271340
rect 517606 271328 517612 271340
rect 517664 271328 517670 271380
rect 51810 271260 51816 271312
rect 51868 271300 51874 271312
rect 104894 271300 104900 271312
rect 51868 271272 104900 271300
rect 51868 271260 51874 271272
rect 104894 271260 104900 271272
rect 104952 271260 104958 271312
rect 183462 271260 183468 271312
rect 183520 271300 183526 271312
rect 197354 271300 197360 271312
rect 183520 271272 197360 271300
rect 183520 271260 183526 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 209222 271260 209228 271312
rect 209280 271300 209286 271312
rect 263594 271300 263600 271312
rect 209280 271272 263600 271300
rect 209280 271260 209286 271272
rect 263594 271260 263600 271272
rect 263652 271260 263658 271312
rect 362586 271260 362592 271312
rect 362644 271300 362650 271312
rect 434714 271300 434720 271312
rect 362644 271272 434720 271300
rect 362644 271260 362650 271272
rect 434714 271260 434720 271272
rect 434772 271260 434778 271312
rect 51718 271192 51724 271244
rect 51776 271232 51782 271244
rect 103514 271232 103520 271244
rect 51776 271204 103520 271232
rect 51776 271192 51782 271204
rect 103514 271192 103520 271204
rect 103572 271192 103578 271244
rect 206554 271192 206560 271244
rect 206612 271232 206618 271244
rect 260834 271232 260840 271244
rect 206612 271204 260840 271232
rect 206612 271192 206618 271204
rect 260834 271192 260840 271204
rect 260892 271192 260898 271244
rect 343542 271192 343548 271244
rect 343600 271232 343606 271244
rect 356974 271232 356980 271244
rect 343600 271204 356980 271232
rect 343600 271192 343606 271204
rect 356974 271192 356980 271204
rect 357032 271192 357038 271244
rect 370866 271192 370872 271244
rect 370924 271232 370930 271244
rect 442994 271232 443000 271244
rect 370924 271204 443000 271232
rect 370924 271192 370930 271204
rect 442994 271192 443000 271204
rect 443052 271192 443058 271244
rect 503622 271192 503628 271244
rect 503680 271232 503686 271244
rect 517698 271232 517704 271244
rect 503680 271204 517704 271232
rect 503680 271192 503686 271204
rect 517698 271192 517704 271204
rect 517756 271192 517762 271244
rect 50246 271124 50252 271176
rect 50304 271164 50310 271176
rect 100754 271164 100760 271176
rect 50304 271136 100760 271164
rect 50304 271124 50310 271136
rect 100754 271124 100760 271136
rect 100812 271124 100818 271176
rect 183462 271124 183468 271176
rect 183520 271164 183526 271176
rect 201586 271164 201592 271176
rect 183520 271136 201592 271164
rect 183520 271124 183526 271136
rect 201586 271124 201592 271136
rect 201644 271124 201650 271176
rect 202414 271124 202420 271176
rect 202472 271164 202478 271176
rect 252554 271164 252560 271176
rect 202472 271136 252560 271164
rect 202472 271124 202478 271136
rect 252554 271124 252560 271136
rect 252612 271124 252618 271176
rect 277118 271124 277124 271176
rect 277176 271164 277182 271176
rect 356606 271164 356612 271176
rect 277176 271136 356612 271164
rect 277176 271124 277182 271136
rect 356606 271124 356612 271136
rect 356664 271164 356670 271176
rect 356882 271164 356888 271176
rect 356664 271136 356888 271164
rect 356664 271124 356670 271136
rect 356882 271124 356888 271136
rect 356940 271124 356946 271176
rect 374914 271124 374920 271176
rect 374972 271164 374978 271176
rect 413094 271164 413100 271176
rect 374972 271136 413100 271164
rect 374972 271124 374978 271136
rect 413094 271124 413100 271136
rect 413152 271124 413158 271176
rect 440142 271124 440148 271176
rect 440200 271164 440206 271176
rect 516594 271164 516600 271176
rect 440200 271136 516600 271164
rect 440200 271124 440206 271136
rect 516594 271124 516600 271136
rect 516652 271124 516658 271176
rect 54662 271056 54668 271108
rect 54720 271096 54726 271108
rect 88334 271096 88340 271108
rect 54720 271068 88340 271096
rect 54720 271056 54726 271068
rect 88334 271056 88340 271068
rect 88392 271056 88398 271108
rect 212166 271056 212172 271108
rect 212224 271096 212230 271108
rect 258258 271096 258264 271108
rect 212224 271068 258264 271096
rect 212224 271056 212230 271068
rect 258258 271056 258264 271068
rect 258316 271056 258322 271108
rect 379054 271056 379060 271108
rect 379112 271096 379118 271108
rect 416038 271096 416044 271108
rect 379112 271068 416044 271096
rect 379112 271056 379118 271068
rect 416038 271056 416044 271068
rect 416096 271056 416102 271108
rect 46106 270988 46112 271040
rect 46164 271028 46170 271040
rect 77294 271028 77300 271040
rect 46164 271000 77300 271028
rect 46164 270988 46170 271000
rect 77294 270988 77300 271000
rect 77352 270988 77358 271040
rect 210694 270988 210700 271040
rect 210752 271028 210758 271040
rect 255314 271028 255320 271040
rect 210752 271000 255320 271028
rect 210752 270988 210758 271000
rect 255314 270988 255320 271000
rect 255372 270988 255378 271040
rect 374822 270988 374828 271040
rect 374880 271028 374886 271040
rect 409874 271028 409880 271040
rect 374880 271000 409880 271028
rect 374880 270988 374886 271000
rect 409874 270988 409880 271000
rect 409932 270988 409938 271040
rect 47762 270920 47768 270972
rect 47820 270960 47826 270972
rect 78674 270960 78680 270972
rect 47820 270932 78680 270960
rect 47820 270920 47826 270932
rect 78674 270920 78680 270932
rect 78732 270920 78738 270972
rect 216122 270920 216128 270972
rect 216180 270960 216186 270972
rect 247034 270960 247040 270972
rect 216180 270932 247040 270960
rect 216180 270920 216186 270932
rect 247034 270920 247040 270932
rect 247092 270920 247098 270972
rect 379146 270920 379152 270972
rect 379204 270960 379210 270972
rect 407114 270960 407120 270972
rect 379204 270932 407120 270960
rect 379204 270920 379210 270932
rect 407114 270920 407120 270932
rect 407172 270920 407178 270972
rect 50338 270444 50344 270496
rect 50396 270484 50402 270496
rect 51810 270484 51816 270496
rect 50396 270456 51816 270484
rect 50396 270444 50402 270456
rect 51810 270444 51816 270456
rect 51868 270444 51874 270496
rect 59814 270444 59820 270496
rect 59872 270484 59878 270496
rect 107654 270484 107660 270496
rect 59872 270456 107660 270484
rect 59872 270444 59878 270456
rect 107654 270444 107660 270456
rect 107712 270444 107718 270496
rect 115842 270444 115848 270496
rect 115900 270484 115906 270496
rect 196986 270484 196992 270496
rect 115900 270456 196992 270484
rect 115900 270444 115906 270456
rect 196986 270444 196992 270456
rect 197044 270444 197050 270496
rect 211706 270444 211712 270496
rect 211764 270484 211770 270496
rect 212166 270484 212172 270496
rect 211764 270456 212172 270484
rect 211764 270444 211770 270456
rect 212166 270444 212172 270456
rect 212224 270444 212230 270496
rect 215110 270444 215116 270496
rect 215168 270484 215174 270496
rect 216398 270484 216404 270496
rect 215168 270456 216404 270484
rect 215168 270444 215174 270456
rect 216398 270444 216404 270456
rect 216456 270444 216462 270496
rect 219802 270444 219808 270496
rect 219860 270484 219866 270496
rect 220630 270484 220636 270496
rect 219860 270456 220636 270484
rect 219860 270444 219866 270456
rect 220630 270444 220636 270456
rect 220688 270484 220694 270496
rect 247034 270484 247040 270496
rect 220688 270456 247040 270484
rect 220688 270444 220694 270456
rect 247034 270444 247040 270456
rect 247092 270444 247098 270496
rect 280062 270444 280068 270496
rect 280120 270484 280126 270496
rect 356606 270484 356612 270496
rect 280120 270456 356612 270484
rect 280120 270444 280126 270456
rect 356606 270444 356612 270456
rect 356664 270484 356670 270496
rect 357066 270484 357072 270496
rect 356664 270456 357072 270484
rect 356664 270444 356670 270456
rect 357066 270444 357072 270456
rect 357124 270444 357130 270496
rect 369762 270444 369768 270496
rect 369820 270484 369826 270496
rect 371694 270484 371700 270496
rect 369820 270456 371700 270484
rect 369820 270444 369826 270456
rect 371694 270444 371700 270456
rect 371752 270444 371758 270496
rect 377030 270444 377036 270496
rect 377088 270484 377094 270496
rect 378042 270484 378048 270496
rect 377088 270456 378048 270484
rect 377088 270444 377094 270456
rect 378042 270444 378048 270456
rect 378100 270484 378106 270496
rect 411254 270484 411260 270496
rect 378100 270456 411260 270484
rect 378100 270444 378106 270456
rect 411254 270444 411260 270456
rect 411312 270444 411318 270496
rect 81434 270376 81440 270428
rect 81492 270416 81498 270428
rect 109034 270416 109040 270428
rect 81492 270388 109040 270416
rect 81492 270376 81498 270388
rect 109034 270376 109040 270388
rect 109092 270376 109098 270428
rect 117222 270376 117228 270428
rect 117280 270416 117286 270428
rect 197170 270416 197176 270428
rect 117280 270388 197176 270416
rect 117280 270376 117286 270388
rect 197170 270376 197176 270388
rect 197228 270376 197234 270428
rect 211614 270376 211620 270428
rect 211672 270416 211678 270428
rect 213086 270416 213092 270428
rect 211672 270388 213092 270416
rect 211672 270376 211678 270388
rect 213086 270376 213092 270388
rect 213144 270376 213150 270428
rect 213638 270376 213644 270428
rect 213696 270416 213702 270428
rect 215662 270416 215668 270428
rect 213696 270388 215668 270416
rect 213696 270376 213702 270388
rect 215662 270376 215668 270388
rect 215720 270376 215726 270428
rect 216674 270376 216680 270428
rect 216732 270416 216738 270428
rect 217226 270416 217232 270428
rect 216732 270388 217232 270416
rect 216732 270376 216738 270388
rect 217226 270376 217232 270388
rect 217284 270416 217290 270428
rect 263594 270416 263600 270428
rect 217284 270388 263600 270416
rect 217284 270376 217290 270388
rect 263594 270376 263600 270388
rect 263652 270376 263658 270428
rect 369670 270376 369676 270428
rect 369728 270416 369734 270428
rect 401686 270416 401692 270428
rect 369728 270388 401692 270416
rect 369728 270376 369734 270388
rect 401686 270376 401692 270388
rect 401744 270376 401750 270428
rect 63494 270308 63500 270360
rect 63552 270348 63558 270360
rect 92474 270348 92480 270360
rect 63552 270320 92480 270348
rect 63552 270308 63558 270320
rect 92474 270308 92480 270320
rect 92532 270308 92538 270360
rect 219158 270308 219164 270360
rect 219216 270348 219222 270360
rect 251174 270348 251180 270360
rect 219216 270320 251180 270348
rect 219216 270308 219222 270320
rect 251174 270308 251180 270320
rect 251232 270308 251238 270360
rect 376294 270308 376300 270360
rect 376352 270348 376358 270360
rect 377122 270348 377128 270360
rect 376352 270320 377128 270348
rect 376352 270308 376358 270320
rect 377122 270308 377128 270320
rect 377180 270308 377186 270360
rect 411346 270348 411352 270360
rect 379808 270320 411352 270348
rect 379808 270292 379836 270320
rect 411346 270308 411352 270320
rect 411404 270308 411410 270360
rect 53926 270240 53932 270292
rect 53984 270280 53990 270292
rect 84194 270280 84200 270292
rect 53984 270252 84200 270280
rect 53984 270240 53990 270252
rect 84194 270240 84200 270252
rect 84252 270240 84258 270292
rect 220722 270240 220728 270292
rect 220780 270280 220786 270292
rect 249794 270280 249800 270292
rect 220780 270252 249800 270280
rect 220780 270240 220786 270252
rect 249794 270240 249800 270252
rect 249852 270240 249858 270292
rect 375098 270240 375104 270292
rect 375156 270280 375162 270292
rect 377490 270280 377496 270292
rect 375156 270252 377496 270280
rect 375156 270240 375162 270252
rect 377490 270240 377496 270252
rect 377548 270240 377554 270292
rect 378594 270240 378600 270292
rect 378652 270280 378658 270292
rect 379790 270280 379796 270292
rect 378652 270252 379796 270280
rect 378652 270240 378658 270252
rect 379790 270240 379796 270252
rect 379848 270240 379854 270292
rect 379882 270240 379888 270292
rect 379940 270280 379946 270292
rect 408494 270280 408500 270292
rect 379940 270252 408500 270280
rect 379940 270240 379946 270252
rect 408494 270240 408500 270252
rect 408552 270240 408558 270292
rect 53834 270172 53840 270224
rect 53892 270212 53898 270224
rect 85574 270212 85580 270224
rect 53892 270184 85580 270212
rect 53892 270172 53898 270184
rect 85574 270172 85580 270184
rect 85632 270172 85638 270224
rect 219342 270172 219348 270224
rect 219400 270212 219406 270224
rect 248506 270212 248512 270224
rect 219400 270184 248512 270212
rect 219400 270172 219406 270184
rect 248506 270172 248512 270184
rect 248564 270172 248570 270224
rect 370958 270172 370964 270224
rect 371016 270212 371022 270224
rect 373626 270212 373632 270224
rect 371016 270184 373632 270212
rect 371016 270172 371022 270184
rect 373626 270172 373632 270184
rect 373684 270212 373690 270224
rect 400214 270212 400220 270224
rect 373684 270184 400220 270212
rect 373684 270172 373690 270184
rect 400214 270172 400220 270184
rect 400272 270172 400278 270224
rect 80054 270104 80060 270156
rect 80112 270144 80118 270156
rect 111794 270144 111800 270156
rect 80112 270116 111800 270144
rect 80112 270104 80118 270116
rect 111794 270104 111800 270116
rect 111852 270104 111858 270156
rect 216766 270104 216772 270156
rect 216824 270144 216830 270156
rect 219618 270144 219624 270156
rect 216824 270116 219624 270144
rect 216824 270104 216830 270116
rect 219618 270104 219624 270116
rect 219676 270144 219682 270156
rect 220722 270144 220728 270156
rect 219676 270116 220728 270144
rect 219676 270104 219682 270116
rect 220722 270104 220728 270116
rect 220780 270104 220786 270156
rect 224218 270104 224224 270156
rect 224276 270144 224282 270156
rect 245654 270144 245660 270156
rect 224276 270116 245660 270144
rect 224276 270104 224282 270116
rect 245654 270104 245660 270116
rect 245712 270104 245718 270156
rect 375650 270104 375656 270156
rect 375708 270144 375714 270156
rect 379698 270144 379704 270156
rect 375708 270116 379704 270144
rect 375708 270104 375714 270116
rect 379698 270104 379704 270116
rect 379756 270144 379762 270156
rect 405734 270144 405740 270156
rect 379756 270116 405740 270144
rect 379756 270104 379762 270116
rect 405734 270104 405740 270116
rect 405792 270104 405798 270156
rect 51810 270036 51816 270088
rect 51868 270076 51874 270088
rect 84654 270076 84660 270088
rect 51868 270048 84660 270076
rect 51868 270036 51874 270048
rect 84654 270036 84660 270048
rect 84712 270036 84718 270088
rect 217042 270036 217048 270088
rect 217100 270076 217106 270088
rect 219066 270076 219072 270088
rect 217100 270048 219072 270076
rect 217100 270036 217106 270048
rect 219066 270036 219072 270048
rect 219124 270076 219130 270088
rect 251266 270076 251272 270088
rect 219124 270048 251272 270076
rect 219124 270036 219130 270048
rect 251266 270036 251272 270048
rect 251324 270036 251330 270088
rect 371694 270036 371700 270088
rect 371752 270076 371758 270088
rect 397454 270076 397460 270088
rect 371752 270048 397460 270076
rect 371752 270036 371758 270048
rect 397454 270036 397460 270048
rect 397512 270036 397518 270088
rect 55950 269968 55956 270020
rect 56008 270008 56014 270020
rect 88334 270008 88340 270020
rect 56008 269980 88340 270008
rect 56008 269968 56014 269980
rect 88334 269968 88340 269980
rect 88392 269968 88398 270020
rect 219250 269968 219256 270020
rect 219308 270008 219314 270020
rect 252554 270008 252560 270020
rect 219308 269980 252560 270008
rect 219308 269968 219314 269980
rect 252554 269968 252560 269980
rect 252612 269968 252618 270020
rect 372522 269968 372528 270020
rect 372580 270008 372586 270020
rect 373902 270008 373908 270020
rect 372580 269980 373908 270008
rect 372580 269968 372586 269980
rect 373902 269968 373908 269980
rect 373960 270008 373966 270020
rect 398834 270008 398840 270020
rect 373960 269980 398840 270008
rect 373960 269968 373966 269980
rect 398834 269968 398840 269980
rect 398892 269968 398898 270020
rect 57974 269900 57980 269952
rect 58032 269940 58038 269952
rect 91094 269940 91100 269952
rect 58032 269912 91100 269940
rect 58032 269900 58038 269912
rect 91094 269900 91100 269912
rect 91152 269900 91158 269952
rect 215662 269900 215668 269952
rect 215720 269940 215726 269952
rect 224126 269940 224132 269952
rect 215720 269912 224132 269940
rect 215720 269900 215726 269912
rect 224126 269900 224132 269912
rect 224184 269900 224190 269952
rect 224402 269900 224408 269952
rect 224460 269940 224466 269952
rect 265158 269940 265164 269952
rect 224460 269912 265164 269940
rect 224460 269900 224466 269912
rect 265158 269900 265164 269912
rect 265216 269900 265222 269952
rect 377490 269900 377496 269952
rect 377548 269940 377554 269952
rect 407114 269940 407120 269952
rect 377548 269912 407120 269940
rect 377548 269900 377554 269912
rect 407114 269900 407120 269912
rect 407172 269900 407178 269952
rect 57054 269832 57060 269884
rect 57112 269872 57118 269884
rect 89714 269872 89720 269884
rect 57112 269844 89720 269872
rect 57112 269832 57118 269844
rect 89714 269832 89720 269844
rect 89772 269832 89778 269884
rect 213086 269832 213092 269884
rect 213144 269872 213150 269884
rect 224218 269872 224224 269884
rect 213144 269844 224224 269872
rect 213144 269832 213150 269844
rect 224218 269832 224224 269844
rect 224276 269832 224282 269884
rect 224310 269832 224316 269884
rect 224368 269872 224374 269884
rect 262214 269872 262220 269884
rect 224368 269844 262220 269872
rect 224368 269832 224374 269844
rect 262214 269832 262220 269844
rect 262272 269832 262278 269884
rect 374362 269832 374368 269884
rect 374420 269872 374426 269884
rect 379882 269872 379888 269884
rect 374420 269844 379888 269872
rect 374420 269832 374426 269844
rect 379882 269832 379888 269844
rect 379940 269832 379946 269884
rect 389266 269832 389272 269884
rect 389324 269872 389330 269884
rect 420914 269872 420920 269884
rect 389324 269844 420920 269872
rect 389324 269832 389330 269844
rect 420914 269832 420920 269844
rect 420972 269832 420978 269884
rect 46658 269764 46664 269816
rect 46716 269804 46722 269816
rect 59814 269804 59820 269816
rect 46716 269776 59820 269804
rect 46716 269764 46722 269776
rect 59814 269764 59820 269776
rect 59872 269764 59878 269816
rect 77846 269764 77852 269816
rect 77904 269804 77910 269816
rect 113174 269804 113180 269816
rect 77904 269776 113180 269804
rect 77904 269764 77910 269776
rect 113174 269764 113180 269776
rect 113232 269764 113238 269816
rect 217870 269764 217876 269816
rect 217928 269804 217934 269816
rect 218606 269804 218612 269816
rect 217928 269776 218612 269804
rect 217928 269764 217934 269776
rect 218606 269764 218612 269776
rect 218664 269804 218670 269816
rect 266354 269804 266360 269816
rect 218664 269776 266360 269804
rect 218664 269764 218670 269776
rect 266354 269764 266360 269776
rect 266412 269764 266418 269816
rect 371786 269764 371792 269816
rect 371844 269804 371850 269816
rect 379146 269804 379152 269816
rect 371844 269776 379152 269804
rect 371844 269764 371850 269776
rect 379146 269764 379152 269776
rect 379204 269764 379210 269816
rect 379606 269764 379612 269816
rect 379664 269804 379670 269816
rect 412910 269804 412916 269816
rect 379664 269776 412916 269804
rect 379664 269764 379670 269776
rect 412910 269764 412916 269776
rect 412968 269764 412974 269816
rect 209406 269696 209412 269748
rect 209464 269736 209470 269748
rect 210786 269736 210792 269748
rect 209464 269708 210792 269736
rect 209464 269696 209470 269708
rect 210786 269696 210792 269708
rect 210844 269736 210850 269748
rect 239122 269736 239128 269748
rect 210844 269708 239128 269736
rect 210844 269696 210850 269708
rect 239122 269696 239128 269708
rect 239180 269696 239186 269748
rect 373718 269696 373724 269748
rect 373776 269736 373782 269748
rect 376202 269736 376208 269748
rect 373776 269708 376208 269736
rect 373776 269696 373782 269708
rect 376202 269696 376208 269708
rect 376260 269736 376266 269748
rect 396074 269736 396080 269748
rect 376260 269708 396080 269736
rect 376260 269696 376266 269708
rect 396074 269696 396080 269708
rect 396132 269696 396138 269748
rect 224126 269628 224132 269680
rect 224184 269668 224190 269680
rect 244274 269668 244280 269680
rect 224184 269640 244280 269668
rect 224184 269628 224190 269640
rect 244274 269628 244280 269640
rect 244332 269628 244338 269680
rect 377122 269628 377128 269680
rect 377180 269668 377186 269680
rect 391934 269668 391940 269680
rect 377180 269640 391940 269668
rect 377180 269628 377186 269640
rect 391934 269628 391940 269640
rect 391992 269628 391998 269680
rect 212166 269560 212172 269612
rect 212224 269600 212230 269612
rect 271874 269600 271880 269612
rect 212224 269572 271880 269600
rect 212224 269560 212230 269572
rect 271874 269560 271880 269572
rect 271932 269560 271938 269612
rect 216398 269492 216404 269544
rect 216456 269532 216462 269544
rect 224310 269532 224316 269544
rect 216456 269504 224316 269532
rect 216456 269492 216462 269504
rect 224310 269492 224316 269504
rect 224368 269492 224374 269544
rect 217962 269424 217968 269476
rect 218020 269464 218026 269476
rect 220630 269464 220636 269476
rect 218020 269436 220636 269464
rect 218020 269424 218026 269436
rect 220630 269424 220636 269436
rect 220688 269424 220694 269476
rect 219250 269288 219256 269340
rect 219308 269328 219314 269340
rect 219802 269328 219808 269340
rect 219308 269300 219808 269328
rect 219308 269288 219314 269300
rect 219802 269288 219808 269300
rect 219860 269288 219866 269340
rect 54754 269220 54760 269272
rect 54812 269260 54818 269272
rect 55950 269260 55956 269272
rect 54812 269232 55956 269260
rect 54812 269220 54818 269232
rect 55950 269220 55956 269232
rect 56008 269220 56014 269272
rect 218514 269220 218520 269272
rect 218572 269260 218578 269272
rect 219618 269260 219624 269272
rect 218572 269232 219624 269260
rect 218572 269220 218578 269232
rect 219618 269220 219624 269232
rect 219676 269260 219682 269272
rect 224402 269260 224408 269272
rect 219676 269232 224408 269260
rect 219676 269220 219682 269232
rect 224402 269220 224408 269232
rect 224460 269220 224466 269272
rect 379146 269152 379152 269204
rect 379204 269192 379210 269204
rect 389174 269192 389180 269204
rect 379204 269164 389180 269192
rect 379204 269152 379210 269164
rect 389174 269152 389180 269164
rect 389232 269152 389238 269204
rect 376478 269084 376484 269136
rect 376536 269124 376542 269136
rect 390554 269124 390560 269136
rect 376536 269096 390560 269124
rect 376536 269084 376542 269096
rect 390554 269084 390560 269096
rect 390612 269084 390618 269136
rect 47946 269016 47952 269068
rect 48004 269056 48010 269068
rect 53834 269056 53840 269068
rect 48004 269028 53840 269056
rect 48004 269016 48010 269028
rect 53834 269016 53840 269028
rect 53892 269056 53898 269068
rect 54570 269056 54576 269068
rect 53892 269028 54576 269056
rect 53892 269016 53898 269028
rect 54570 269016 54576 269028
rect 54628 269016 54634 269068
rect 214466 269016 214472 269068
rect 214524 269056 214530 269068
rect 216030 269056 216036 269068
rect 214524 269028 216036 269056
rect 214524 269016 214530 269028
rect 216030 269016 216036 269028
rect 216088 269016 216094 269068
rect 219710 269016 219716 269068
rect 219768 269056 219774 269068
rect 253934 269056 253940 269068
rect 219768 269028 253940 269056
rect 219768 269016 219774 269028
rect 253934 269016 253940 269028
rect 253992 269016 253998 269068
rect 376570 269016 376576 269068
rect 376628 269056 376634 269068
rect 379054 269056 379060 269068
rect 376628 269028 379060 269056
rect 376628 269016 376634 269028
rect 379054 269016 379060 269028
rect 379112 269016 379118 269068
rect 383562 269016 383568 269068
rect 383620 269056 383626 269068
rect 436186 269056 436192 269068
rect 383620 269028 436192 269056
rect 383620 269016 383626 269028
rect 436186 269016 436192 269028
rect 436244 269016 436250 269068
rect 45370 268948 45376 269000
rect 45428 268988 45434 269000
rect 144914 268988 144920 269000
rect 45428 268960 144920 268988
rect 45428 268948 45434 268960
rect 144914 268948 144920 268960
rect 144972 268948 144978 269000
rect 213546 268948 213552 269000
rect 213604 268988 213610 269000
rect 242894 268988 242900 269000
rect 213604 268960 242900 268988
rect 213604 268948 213610 268960
rect 242894 268948 242900 268960
rect 242952 268948 242958 269000
rect 372246 268948 372252 269000
rect 372304 268988 372310 269000
rect 373810 268988 373816 269000
rect 372304 268960 373816 268988
rect 372304 268948 372310 268960
rect 373810 268948 373816 268960
rect 373868 268988 373874 269000
rect 433334 268988 433340 269000
rect 373868 268960 433340 268988
rect 373868 268948 373874 268960
rect 433334 268948 433340 268960
rect 433392 268948 433398 269000
rect 42242 268880 42248 268932
rect 42300 268920 42306 268932
rect 107746 268920 107752 268932
rect 42300 268892 107752 268920
rect 42300 268880 42306 268892
rect 107746 268880 107752 268892
rect 107804 268880 107810 268932
rect 213270 268880 213276 268932
rect 213328 268920 213334 268932
rect 215846 268920 215852 268932
rect 213328 268892 215852 268920
rect 213328 268880 213334 268892
rect 215846 268880 215852 268892
rect 215904 268880 215910 268932
rect 231854 268880 231860 268932
rect 231912 268920 231918 268932
rect 259454 268920 259460 268932
rect 231912 268892 259460 268920
rect 231912 268880 231918 268892
rect 259454 268880 259460 268892
rect 259512 268880 259518 268932
rect 375926 268880 375932 268932
rect 375984 268920 375990 268932
rect 376754 268920 376760 268932
rect 375984 268892 376760 268920
rect 375984 268880 375990 268892
rect 376754 268880 376760 268892
rect 376812 268920 376818 268932
rect 383378 268920 383384 268932
rect 376812 268892 383384 268920
rect 376812 268880 376818 268892
rect 383378 268880 383384 268892
rect 383436 268880 383442 268932
rect 383470 268880 383476 268932
rect 383528 268920 383534 268932
rect 416774 268920 416780 268932
rect 383528 268892 416780 268920
rect 383528 268880 383534 268892
rect 416774 268880 416780 268892
rect 416832 268880 416838 268932
rect 49142 268812 49148 268864
rect 49200 268852 49206 268864
rect 110414 268852 110420 268864
rect 49200 268824 110420 268852
rect 49200 268812 49206 268824
rect 110414 268812 110420 268824
rect 110472 268812 110478 268864
rect 216490 268812 216496 268864
rect 216548 268852 216554 268864
rect 230474 268852 230480 268864
rect 216548 268824 230480 268852
rect 216548 268812 216554 268824
rect 230474 268812 230480 268824
rect 230532 268852 230538 268864
rect 259546 268852 259552 268864
rect 230532 268824 259552 268852
rect 230532 268812 230538 268824
rect 259546 268812 259552 268824
rect 259604 268812 259610 268864
rect 379974 268812 379980 268864
rect 380032 268852 380038 268864
rect 414014 268852 414020 268864
rect 380032 268824 414020 268852
rect 380032 268812 380038 268824
rect 414014 268812 414020 268824
rect 414072 268812 414078 268864
rect 43898 268744 43904 268796
rect 43956 268784 43962 268796
rect 57974 268784 57980 268796
rect 43956 268756 57980 268784
rect 43956 268744 43962 268756
rect 57974 268744 57980 268756
rect 58032 268744 58038 268796
rect 229186 268744 229192 268796
rect 229244 268784 229250 268796
rect 260834 268784 260840 268796
rect 229244 268756 260840 268784
rect 229244 268744 229250 268756
rect 260834 268744 260840 268756
rect 260892 268744 260898 268796
rect 379238 268744 379244 268796
rect 379296 268784 379302 268796
rect 409874 268784 409880 268796
rect 379296 268756 409880 268784
rect 379296 268744 379302 268756
rect 409874 268744 409880 268756
rect 409932 268744 409938 268796
rect 43806 268676 43812 268728
rect 43864 268716 43870 268728
rect 57054 268716 57060 268728
rect 43864 268688 57060 268716
rect 43864 268676 43870 268688
rect 57054 268676 57060 268688
rect 57112 268676 57118 268728
rect 215846 268676 215852 268728
rect 215904 268716 215910 268728
rect 255314 268716 255320 268728
rect 215904 268688 255320 268716
rect 215904 268676 215910 268688
rect 255314 268676 255320 268688
rect 255372 268676 255378 268728
rect 389174 268676 389180 268728
rect 389232 268716 389238 268728
rect 419534 268716 419540 268728
rect 389232 268688 419540 268716
rect 389232 268676 389238 268688
rect 419534 268676 419540 268688
rect 419592 268676 419598 268728
rect 46842 268608 46848 268660
rect 46900 268648 46906 268660
rect 53926 268648 53932 268660
rect 46900 268620 53932 268648
rect 46900 268608 46906 268620
rect 53926 268608 53932 268620
rect 53984 268648 53990 268660
rect 54478 268648 54484 268660
rect 53984 268620 54484 268648
rect 53984 268608 53990 268620
rect 54478 268608 54484 268620
rect 54536 268608 54542 268660
rect 207934 268608 207940 268660
rect 207992 268648 207998 268660
rect 218514 268648 218520 268660
rect 207992 268620 218520 268648
rect 207992 268608 207998 268620
rect 218514 268608 218520 268620
rect 218572 268648 218578 268660
rect 258074 268648 258080 268660
rect 218572 268620 258080 268648
rect 218572 268608 218578 268620
rect 258074 268608 258080 268620
rect 258132 268608 258138 268660
rect 374914 268608 374920 268660
rect 374972 268648 374978 268660
rect 375742 268648 375748 268660
rect 374972 268620 375748 268648
rect 374972 268608 374978 268620
rect 375742 268608 375748 268620
rect 375800 268648 375806 268660
rect 383470 268648 383476 268660
rect 375800 268620 383476 268648
rect 375800 268608 375806 268620
rect 383470 268608 383476 268620
rect 383528 268608 383534 268660
rect 390554 268608 390560 268660
rect 390612 268648 390618 268660
rect 418246 268648 418252 268660
rect 390612 268620 418252 268648
rect 390612 268608 390618 268620
rect 418246 268608 418252 268620
rect 418304 268608 418310 268660
rect 50430 268540 50436 268592
rect 50488 268580 50494 268592
rect 63494 268580 63500 268592
rect 50488 268552 63500 268580
rect 50488 268540 50494 268552
rect 63494 268540 63500 268552
rect 63552 268540 63558 268592
rect 216030 268540 216036 268592
rect 216088 268580 216094 268592
rect 256694 268580 256700 268592
rect 216088 268552 256700 268580
rect 216088 268540 216094 268552
rect 256694 268540 256700 268552
rect 256752 268540 256758 268592
rect 377306 268540 377312 268592
rect 377364 268580 377370 268592
rect 403526 268580 403532 268592
rect 377364 268552 403532 268580
rect 377364 268540 377370 268552
rect 403526 268540 403532 268552
rect 403584 268540 403590 268592
rect 43714 268472 43720 268524
rect 43772 268512 43778 268524
rect 46474 268512 46480 268524
rect 43772 268484 46480 268512
rect 43772 268472 43778 268484
rect 46474 268472 46480 268484
rect 46532 268512 46538 268524
rect 80054 268512 80060 268524
rect 46532 268484 80060 268512
rect 46532 268472 46538 268484
rect 80054 268472 80060 268484
rect 80112 268472 80118 268524
rect 209498 268472 209504 268524
rect 209556 268512 209562 268524
rect 213454 268512 213460 268524
rect 209556 268484 213460 268512
rect 209556 268472 209562 268484
rect 213454 268472 213460 268484
rect 213512 268512 213518 268524
rect 269114 268512 269120 268524
rect 213512 268484 269120 268512
rect 213512 268472 213518 268484
rect 269114 268472 269120 268484
rect 269172 268472 269178 268524
rect 391934 268472 391940 268524
rect 391992 268512 391998 268524
rect 418154 268512 418160 268524
rect 391992 268484 418160 268512
rect 391992 268472 391998 268484
rect 418154 268472 418160 268484
rect 418212 268472 418218 268524
rect 43622 268404 43628 268456
rect 43680 268444 43686 268456
rect 47854 268444 47860 268456
rect 43680 268416 47860 268444
rect 43680 268404 43686 268416
rect 47854 268404 47860 268416
rect 47912 268444 47918 268456
rect 81434 268444 81440 268456
rect 47912 268416 81440 268444
rect 47912 268404 47918 268416
rect 81434 268404 81440 268416
rect 81492 268404 81498 268456
rect 209590 268404 209596 268456
rect 209648 268444 209654 268456
rect 213362 268444 213368 268456
rect 209648 268416 213368 268444
rect 209648 268404 209654 268416
rect 213362 268404 213368 268416
rect 213420 268444 213426 268456
rect 270494 268444 270500 268456
rect 213420 268416 270500 268444
rect 213420 268404 213426 268416
rect 270494 268404 270500 268416
rect 270552 268404 270558 268456
rect 45462 268336 45468 268388
rect 45520 268376 45526 268388
rect 50430 268376 50436 268388
rect 45520 268348 50436 268376
rect 45520 268336 45526 268348
rect 50430 268336 50436 268348
rect 50488 268336 50494 268388
rect 53098 268336 53104 268388
rect 53156 268376 53162 268388
rect 106366 268376 106372 268388
rect 53156 268348 106372 268376
rect 53156 268336 53162 268348
rect 106366 268336 106372 268348
rect 106424 268336 106430 268388
rect 206830 268336 206836 268388
rect 206888 268376 206894 268388
rect 212074 268376 212080 268388
rect 206888 268348 212080 268376
rect 206888 268336 206894 268348
rect 212074 268336 212080 268348
rect 212132 268376 212138 268388
rect 273162 268376 273168 268388
rect 212132 268348 273168 268376
rect 212132 268336 212138 268348
rect 273162 268336 273168 268348
rect 273220 268336 273226 268388
rect 379054 268336 379060 268388
rect 379112 268376 379118 268388
rect 404354 268376 404360 268388
rect 379112 268348 404360 268376
rect 379112 268336 379118 268348
rect 404354 268336 404360 268348
rect 404412 268336 404418 268388
rect 44910 268268 44916 268320
rect 44968 268308 44974 268320
rect 147674 268308 147680 268320
rect 44968 268280 147680 268308
rect 44968 268268 44974 268280
rect 147674 268268 147680 268280
rect 147732 268268 147738 268320
rect 216306 268268 216312 268320
rect 216364 268308 216370 268320
rect 231854 268308 231860 268320
rect 216364 268280 231860 268308
rect 216364 268268 216370 268280
rect 231854 268268 231860 268280
rect 231912 268268 231918 268320
rect 215110 268200 215116 268252
rect 215168 268240 215174 268252
rect 218330 268240 218336 268252
rect 215168 268212 218336 268240
rect 215168 268200 215174 268212
rect 218330 268200 218336 268212
rect 218388 268240 218394 268252
rect 244366 268240 244372 268252
rect 218388 268212 244372 268240
rect 218388 268200 218394 268212
rect 244366 268200 244372 268212
rect 244424 268200 244430 268252
rect 375558 268200 375564 268252
rect 375616 268240 375622 268252
rect 377306 268240 377312 268252
rect 375616 268212 377312 268240
rect 375616 268200 375622 268212
rect 377306 268200 377312 268212
rect 377364 268200 377370 268252
rect 357158 253960 357164 253972
rect 356440 253932 357164 253960
rect 191742 253852 191748 253904
rect 191800 253892 191806 253904
rect 201402 253892 201408 253904
rect 191800 253864 201408 253892
rect 191800 253852 191806 253864
rect 201402 253852 201408 253864
rect 201460 253892 201466 253904
rect 202874 253892 202880 253904
rect 201460 253864 202880 253892
rect 201460 253852 201466 253864
rect 202874 253852 202880 253864
rect 202932 253852 202938 253904
rect 340782 253852 340788 253904
rect 340840 253892 340846 253904
rect 356440 253892 356468 253932
rect 357158 253920 357164 253932
rect 357216 253960 357222 253972
rect 357526 253960 357532 253972
rect 357216 253932 357532 253960
rect 357216 253920 357222 253932
rect 357526 253920 357532 253932
rect 357584 253920 357590 253972
rect 340840 253864 356468 253892
rect 340840 253852 340846 253864
rect 500862 253308 500868 253360
rect 500920 253348 500926 253360
rect 517790 253348 517796 253360
rect 500920 253320 517796 253348
rect 500920 253308 500926 253320
rect 517790 253308 517796 253320
rect 517848 253308 517854 253360
rect 180518 253240 180524 253292
rect 180576 253280 180582 253292
rect 197630 253280 197636 253292
rect 180576 253252 197636 253280
rect 180576 253240 180582 253252
rect 197630 253240 197636 253252
rect 197688 253280 197694 253292
rect 198090 253280 198096 253292
rect 197688 253252 198096 253280
rect 197688 253240 197694 253252
rect 198090 253240 198096 253252
rect 198148 253240 198154 253292
rect 339402 253240 339408 253292
rect 339460 253280 339466 253292
rect 360194 253280 360200 253292
rect 339460 253252 360200 253280
rect 339460 253240 339466 253252
rect 360194 253240 360200 253252
rect 360252 253240 360258 253292
rect 499206 253240 499212 253292
rect 499264 253280 499270 253292
rect 517698 253280 517704 253292
rect 499264 253252 517704 253280
rect 499264 253240 499270 253252
rect 517698 253240 517704 253252
rect 517756 253280 517762 253292
rect 517974 253280 517980 253292
rect 517756 253252 517980 253280
rect 517756 253240 517762 253252
rect 517974 253240 517980 253252
rect 518032 253240 518038 253292
rect 179322 253172 179328 253224
rect 179380 253212 179386 253224
rect 197538 253212 197544 253224
rect 179380 253184 197544 253212
rect 179380 253172 179386 253184
rect 197538 253172 197544 253184
rect 197596 253172 197602 253224
rect 351822 253172 351828 253224
rect 351880 253212 351886 253224
rect 358078 253212 358084 253224
rect 351880 253184 358084 253212
rect 351880 253172 351886 253184
rect 358078 253172 358084 253184
rect 358136 253172 358142 253224
rect 517790 253172 517796 253224
rect 517848 253212 517854 253224
rect 518066 253212 518072 253224
rect 517848 253184 518072 253212
rect 517848 253172 517854 253184
rect 518066 253172 518072 253184
rect 518124 253172 518130 253224
rect 510890 252560 510896 252612
rect 510948 252600 510954 252612
rect 517514 252600 517520 252612
rect 510948 252572 517520 252600
rect 510948 252560 510954 252572
rect 517514 252560 517520 252572
rect 517572 252560 517578 252612
rect 58710 252492 58716 252544
rect 58768 252532 58774 252544
rect 60826 252532 60832 252544
rect 58768 252504 60832 252532
rect 58768 252492 58774 252504
rect 60826 252492 60832 252504
rect 60884 252492 60890 252544
rect 374822 252492 374828 252544
rect 374880 252532 374886 252544
rect 375282 252532 375288 252544
rect 374880 252504 375288 252532
rect 374880 252492 374886 252504
rect 375282 252492 375288 252504
rect 375340 252532 375346 252544
rect 436094 252532 436100 252544
rect 375340 252504 436100 252532
rect 375340 252492 375346 252504
rect 436094 252492 436100 252504
rect 436152 252492 436158 252544
rect 373626 252424 373632 252476
rect 373684 252464 373690 252476
rect 375834 252464 375840 252476
rect 373684 252436 375840 252464
rect 373684 252424 373690 252436
rect 375834 252424 375840 252436
rect 375892 252464 375898 252476
rect 434714 252464 434720 252476
rect 375892 252436 434720 252464
rect 375892 252424 375898 252436
rect 434714 252424 434720 252436
rect 434772 252424 434778 252476
rect 372154 252356 372160 252408
rect 372212 252396 372218 252408
rect 372430 252396 372436 252408
rect 372212 252368 372436 252396
rect 372212 252356 372218 252368
rect 372430 252356 372436 252368
rect 372488 252396 372494 252408
rect 429194 252396 429200 252408
rect 372488 252368 429200 252396
rect 372488 252356 372494 252368
rect 429194 252356 429200 252368
rect 429252 252356 429258 252408
rect 55858 252152 55864 252204
rect 55916 252192 55922 252204
rect 60734 252192 60740 252204
rect 55916 252164 60740 252192
rect 55916 252152 55922 252164
rect 60734 252152 60740 252164
rect 60792 252152 60798 252204
rect 75822 252016 75828 252068
rect 75880 252056 75886 252068
rect 98638 252056 98644 252068
rect 75880 252028 98644 252056
rect 75880 252016 75886 252028
rect 98638 252016 98644 252028
rect 98696 252016 98702 252068
rect 377122 252016 377128 252068
rect 377180 252056 377186 252068
rect 389174 252056 389180 252068
rect 377180 252028 389180 252056
rect 377180 252016 377186 252028
rect 389174 252016 389180 252028
rect 389232 252016 389238 252068
rect 52914 251948 52920 252000
rect 52972 251988 52978 252000
rect 83458 251988 83464 252000
rect 52972 251960 83464 251988
rect 52972 251948 52978 251960
rect 83458 251948 83464 251960
rect 83516 251948 83522 252000
rect 371050 251948 371056 252000
rect 371108 251988 371114 252000
rect 379698 251988 379704 252000
rect 371108 251960 379704 251988
rect 371108 251948 371114 251960
rect 379698 251948 379704 251960
rect 379756 251988 379762 252000
rect 425698 251988 425704 252000
rect 379756 251960 425704 251988
rect 379756 251948 379762 251960
rect 425698 251948 425704 251960
rect 425756 251948 425762 252000
rect 58618 251880 58624 251932
rect 58676 251920 58682 251932
rect 106274 251920 106280 251932
rect 58676 251892 106280 251920
rect 58676 251880 58682 251892
rect 106274 251880 106280 251892
rect 106332 251880 106338 251932
rect 214466 251880 214472 251932
rect 214524 251920 214530 251932
rect 229094 251920 229100 251932
rect 214524 251892 229100 251920
rect 214524 251880 214530 251892
rect 229094 251880 229100 251892
rect 229152 251880 229158 251932
rect 370406 251880 370412 251932
rect 370464 251920 370470 251932
rect 373534 251920 373540 251932
rect 370464 251892 373540 251920
rect 370464 251880 370470 251892
rect 373534 251880 373540 251892
rect 373592 251920 373598 251932
rect 421558 251920 421564 251932
rect 373592 251892 421564 251920
rect 373592 251880 373598 251892
rect 421558 251880 421564 251892
rect 421616 251880 421622 251932
rect 57606 251812 57612 251864
rect 57664 251852 57670 251864
rect 104894 251852 104900 251864
rect 57664 251824 104900 251852
rect 57664 251812 57670 251824
rect 104894 251812 104900 251824
rect 104952 251812 104958 251864
rect 214834 251812 214840 251864
rect 214892 251852 214898 251864
rect 230474 251852 230480 251864
rect 214892 251824 230480 251852
rect 214892 251812 214898 251824
rect 230474 251812 230480 251824
rect 230532 251812 230538 251864
rect 369578 251812 369584 251864
rect 369636 251852 369642 251864
rect 372430 251852 372436 251864
rect 369636 251824 372436 251852
rect 369636 251812 369642 251824
rect 372430 251812 372436 251824
rect 372488 251852 372494 251864
rect 427078 251852 427084 251864
rect 372488 251824 427084 251852
rect 372488 251812 372494 251824
rect 427078 251812 427084 251824
rect 427136 251812 427142 251864
rect 50522 251132 50528 251184
rect 50580 251172 50586 251184
rect 75822 251172 75828 251184
rect 50580 251144 75828 251172
rect 50580 251132 50586 251144
rect 75822 251132 75828 251144
rect 75880 251132 75886 251184
rect 43990 251064 43996 251116
rect 44048 251104 44054 251116
rect 56870 251104 56876 251116
rect 44048 251076 56876 251104
rect 44048 251064 44054 251076
rect 56870 251064 56876 251076
rect 56928 251104 56934 251116
rect 57606 251104 57612 251116
rect 56928 251076 57612 251104
rect 56928 251064 56934 251076
rect 57606 251064 57612 251076
rect 57664 251064 57670 251116
rect 42610 250996 42616 251048
rect 42668 251036 42674 251048
rect 52914 251036 52920 251048
rect 42668 251008 52920 251036
rect 42668 250996 42674 251008
rect 52914 250996 52920 251008
rect 52972 250996 52978 251048
rect 519446 183540 519452 183592
rect 519504 183580 519510 183592
rect 520182 183580 520188 183592
rect 519504 183552 520188 183580
rect 519504 183540 519510 183552
rect 520182 183540 520188 183552
rect 520240 183580 520246 183592
rect 580258 183580 580264 183592
rect 520240 183552 580264 183580
rect 520240 183540 520246 183552
rect 580258 183540 580264 183552
rect 580316 183540 580322 183592
rect 520090 183472 520096 183524
rect 520148 183512 520154 183524
rect 580350 183512 580356 183524
rect 520148 183484 580356 183512
rect 520148 183472 520154 183484
rect 580350 183472 580356 183484
rect 580408 183472 580414 183524
rect 204990 177964 204996 178016
rect 205048 178004 205054 178016
rect 217042 178004 217048 178016
rect 205048 177976 217048 178004
rect 205048 177964 205054 177976
rect 217042 177964 217048 177976
rect 217100 177964 217106 178016
rect 363874 177964 363880 178016
rect 363932 178004 363938 178016
rect 377030 178004 377036 178016
rect 363932 177976 377036 178004
rect 363932 177964 363938 177976
rect 377030 177964 377036 177976
rect 377088 177964 377094 178016
rect 216766 176808 216772 176860
rect 216824 176848 216830 176860
rect 217042 176848 217048 176860
rect 216824 176820 217048 176848
rect 216824 176808 216830 176820
rect 217042 176808 217048 176820
rect 217100 176808 217106 176860
rect 202874 176604 202880 176656
rect 202932 176644 202938 176656
rect 216674 176644 216680 176656
rect 202932 176616 216680 176644
rect 202932 176604 202938 176616
rect 216674 176604 216680 176616
rect 216732 176604 216738 176656
rect 202138 176128 202144 176180
rect 202196 176168 202202 176180
rect 202874 176168 202880 176180
rect 202196 176140 202880 176168
rect 202196 176128 202202 176140
rect 202874 176128 202880 176140
rect 202932 176128 202938 176180
rect 358078 175924 358084 175976
rect 358136 175964 358142 175976
rect 376938 175964 376944 175976
rect 358136 175936 376944 175964
rect 358136 175924 358142 175936
rect 376938 175924 376944 175936
rect 376996 175924 377002 175976
rect 207658 175176 207664 175228
rect 207716 175216 207722 175228
rect 217134 175216 217140 175228
rect 207716 175188 217140 175216
rect 207716 175176 207722 175188
rect 217134 175176 217140 175188
rect 217192 175176 217198 175228
rect 365254 175176 365260 175228
rect 365312 175216 365318 175228
rect 377398 175216 377404 175228
rect 365312 175188 377404 175216
rect 365312 175176 365318 175188
rect 377398 175176 377404 175188
rect 377456 175176 377462 175228
rect 216766 175108 216772 175160
rect 216824 175148 216830 175160
rect 217042 175148 217048 175160
rect 216824 175120 217048 175148
rect 216824 175108 216830 175120
rect 217042 175108 217048 175120
rect 217100 175108 217106 175160
rect 51994 166948 52000 167000
rect 52052 166988 52058 167000
rect 101030 166988 101036 167000
rect 52052 166960 101036 166988
rect 52052 166948 52058 166960
rect 101030 166948 101036 166960
rect 101088 166948 101094 167000
rect 197446 166948 197452 167000
rect 197504 166988 197510 167000
rect 201494 166988 201500 167000
rect 197504 166960 201500 166988
rect 197504 166948 197510 166960
rect 201494 166948 201500 166960
rect 201552 166948 201558 167000
rect 362494 166948 362500 167000
rect 362552 166988 362558 167000
rect 423398 166988 423404 167000
rect 362552 166960 423404 166988
rect 362552 166948 362558 166960
rect 423398 166948 423404 166960
rect 423456 166948 423462 167000
rect 50890 166880 50896 166932
rect 50948 166920 50954 166932
rect 103514 166920 103520 166932
rect 50948 166892 103520 166920
rect 50948 166880 50954 166892
rect 103514 166880 103520 166892
rect 103572 166880 103578 166932
rect 358262 166880 358268 166932
rect 358320 166920 358326 166932
rect 418430 166920 418436 166932
rect 358320 166892 418436 166920
rect 358320 166880 358326 166892
rect 418430 166880 418436 166892
rect 418488 166880 418494 166932
rect 50798 166812 50804 166864
rect 50856 166852 50862 166864
rect 108298 166852 108304 166864
rect 50856 166824 108304 166852
rect 50856 166812 50862 166824
rect 108298 166812 108304 166824
rect 108356 166812 108362 166864
rect 214742 166812 214748 166864
rect 214800 166852 214806 166864
rect 260926 166852 260932 166864
rect 214800 166824 260932 166852
rect 214800 166812 214806 166824
rect 260926 166812 260932 166824
rect 260984 166812 260990 166864
rect 358354 166812 358360 166864
rect 358412 166852 358418 166864
rect 421006 166852 421012 166864
rect 358412 166824 421012 166852
rect 358412 166812 358418 166824
rect 421006 166812 421012 166824
rect 421064 166812 421070 166864
rect 58986 166744 58992 166796
rect 59044 166784 59050 166796
rect 140866 166784 140872 166796
rect 59044 166756 140872 166784
rect 59044 166744 59050 166756
rect 140866 166744 140872 166756
rect 140924 166744 140930 166796
rect 203518 166744 203524 166796
rect 203576 166784 203582 166796
rect 265894 166784 265900 166796
rect 203576 166756 265900 166784
rect 203576 166744 203582 166756
rect 265894 166744 265900 166756
rect 265952 166744 265958 166796
rect 356790 166744 356796 166796
rect 356848 166784 356854 166796
rect 445846 166784 445852 166796
rect 356848 166756 445852 166784
rect 356848 166744 356854 166756
rect 445846 166744 445852 166756
rect 445904 166744 445910 166796
rect 56226 166676 56232 166728
rect 56284 166716 56290 166728
rect 138474 166716 138480 166728
rect 56284 166688 138480 166716
rect 56284 166676 56290 166688
rect 138474 166676 138480 166688
rect 138532 166676 138538 166728
rect 203702 166676 203708 166728
rect 203760 166716 203766 166728
rect 270862 166716 270868 166728
rect 203760 166688 270868 166716
rect 203760 166676 203766 166688
rect 270862 166676 270868 166688
rect 270920 166676 270926 166728
rect 369302 166676 369308 166728
rect 369360 166716 369366 166728
rect 470962 166716 470968 166728
rect 369360 166688 470968 166716
rect 369360 166676 369366 166688
rect 470962 166676 470968 166688
rect 471020 166676 471026 166728
rect 59998 166608 60004 166660
rect 60056 166648 60062 166660
rect 145926 166648 145932 166660
rect 60056 166620 145932 166648
rect 60056 166608 60062 166620
rect 145926 166608 145932 166620
rect 145984 166608 145990 166660
rect 204898 166608 204904 166660
rect 204956 166648 204962 166660
rect 285950 166648 285956 166660
rect 204956 166620 285956 166648
rect 204956 166608 204962 166620
rect 285950 166608 285956 166620
rect 286008 166608 286014 166660
rect 373442 166608 373448 166660
rect 373500 166648 373506 166660
rect 475838 166648 475844 166660
rect 373500 166620 475844 166648
rect 373500 166608 373506 166620
rect 475838 166608 475844 166620
rect 475896 166608 475902 166660
rect 59170 166540 59176 166592
rect 59228 166580 59234 166592
rect 148502 166580 148508 166592
rect 59228 166552 148508 166580
rect 59228 166540 59234 166552
rect 148502 166540 148508 166552
rect 148560 166540 148566 166592
rect 210602 166540 210608 166592
rect 210660 166580 210666 166592
rect 295886 166580 295892 166592
rect 210660 166552 295892 166580
rect 210660 166540 210666 166552
rect 295886 166540 295892 166552
rect 295944 166540 295950 166592
rect 370774 166540 370780 166592
rect 370832 166580 370838 166592
rect 473446 166580 473452 166592
rect 370832 166552 473452 166580
rect 370832 166540 370838 166552
rect 473446 166540 473452 166552
rect 473504 166540 473510 166592
rect 59906 166472 59912 166524
rect 59964 166512 59970 166524
rect 150894 166512 150900 166524
rect 59964 166484 150900 166512
rect 59964 166472 59970 166484
rect 150894 166472 150900 166484
rect 150952 166472 150958 166524
rect 206462 166472 206468 166524
rect 206520 166512 206526 166524
rect 293402 166512 293408 166524
rect 206520 166484 293408 166512
rect 206520 166472 206526 166484
rect 293402 166472 293408 166484
rect 293460 166472 293466 166524
rect 372062 166472 372068 166524
rect 372120 166512 372126 166524
rect 480898 166512 480904 166524
rect 372120 166484 480904 166512
rect 372120 166472 372126 166484
rect 480898 166472 480904 166484
rect 480956 166472 480962 166524
rect 58894 166404 58900 166456
rect 58952 166444 58958 166456
rect 153286 166444 153292 166456
rect 58952 166416 153292 166444
rect 58952 166404 58958 166416
rect 153286 166404 153292 166416
rect 153344 166404 153350 166456
rect 203610 166404 203616 166456
rect 203668 166444 203674 166456
rect 291010 166444 291016 166456
rect 203668 166416 291016 166444
rect 203668 166404 203674 166416
rect 291010 166404 291016 166416
rect 291068 166404 291074 166456
rect 367922 166404 367928 166456
rect 367980 166444 367986 166456
rect 478414 166444 478420 166456
rect 367980 166416 478420 166444
rect 367980 166404 367986 166416
rect 478414 166404 478420 166416
rect 478472 166404 478478 166456
rect 41046 166336 41052 166388
rect 41104 166376 41110 166388
rect 163314 166376 163320 166388
rect 41104 166348 163320 166376
rect 41104 166336 41110 166348
rect 163314 166336 163320 166348
rect 163372 166336 163378 166388
rect 209130 166336 209136 166388
rect 209188 166376 209194 166388
rect 298462 166376 298468 166388
rect 209188 166348 298468 166376
rect 209188 166336 209194 166348
rect 298462 166336 298468 166348
rect 298520 166336 298526 166388
rect 365162 166336 365168 166388
rect 365220 166376 365226 166388
rect 483382 166376 483388 166388
rect 365220 166348 483388 166376
rect 365220 166336 365226 166348
rect 483382 166336 483388 166348
rect 483440 166336 483446 166388
rect 41138 166268 41144 166320
rect 41196 166308 41202 166320
rect 165890 166308 165896 166320
rect 41196 166280 165896 166308
rect 41196 166268 41202 166280
rect 165890 166268 165896 166280
rect 165948 166268 165954 166320
rect 202322 166268 202328 166320
rect 202380 166308 202386 166320
rect 305914 166308 305920 166320
rect 202380 166280 305920 166308
rect 202380 166268 202386 166280
rect 305914 166268 305920 166280
rect 305972 166268 305978 166320
rect 366634 166268 366640 166320
rect 366692 166308 366698 166320
rect 485958 166308 485964 166320
rect 366692 166280 485964 166308
rect 366692 166268 366698 166280
rect 485958 166268 485964 166280
rect 486016 166268 486022 166320
rect 49510 166200 49516 166252
rect 49568 166240 49574 166252
rect 98454 166240 98460 166252
rect 49568 166212 98460 166240
rect 49568 166200 49574 166212
rect 98454 166200 98460 166212
rect 98512 166200 98518 166252
rect 374638 166200 374644 166252
rect 374696 166240 374702 166252
rect 430942 166240 430948 166252
rect 374696 166212 430948 166240
rect 374696 166200 374702 166212
rect 430942 166200 430948 166212
rect 431000 166200 431006 166252
rect 50706 166132 50712 166184
rect 50764 166172 50770 166184
rect 96062 166172 96068 166184
rect 50764 166144 96068 166172
rect 50764 166132 50770 166144
rect 96062 166132 96068 166144
rect 96120 166132 96126 166184
rect 373350 166132 373356 166184
rect 373408 166172 373414 166184
rect 428182 166172 428188 166184
rect 373408 166144 428188 166172
rect 373408 166132 373414 166144
rect 428182 166132 428188 166144
rect 428240 166132 428246 166184
rect 357618 165588 357624 165640
rect 357676 165628 357682 165640
rect 360286 165628 360292 165640
rect 357676 165600 360292 165628
rect 357676 165588 357682 165600
rect 360286 165588 360292 165600
rect 360344 165588 360350 165640
rect 373626 165588 373632 165640
rect 373684 165628 373690 165640
rect 373810 165628 373816 165640
rect 373684 165600 373816 165628
rect 373684 165588 373690 165600
rect 373810 165588 373816 165600
rect 373868 165628 373874 165640
rect 433334 165628 433340 165640
rect 373868 165600 433340 165628
rect 373868 165588 373874 165600
rect 433334 165588 433340 165600
rect 433392 165588 433398 165640
rect 50522 165520 50528 165572
rect 50580 165560 50586 165572
rect 51626 165560 51632 165572
rect 50580 165532 51632 165560
rect 50580 165520 50586 165532
rect 51626 165520 51632 165532
rect 51684 165520 51690 165572
rect 54202 165520 54208 165572
rect 54260 165560 54266 165572
rect 132494 165560 132500 165572
rect 54260 165532 132500 165560
rect 54260 165520 54266 165532
rect 132494 165520 132500 165532
rect 132552 165520 132558 165572
rect 209038 165520 209044 165572
rect 209096 165560 209102 165572
rect 325878 165560 325884 165572
rect 209096 165532 325884 165560
rect 209096 165520 209102 165532
rect 325878 165520 325884 165532
rect 325936 165520 325942 165572
rect 343266 165520 343272 165572
rect 343324 165560 343330 165572
rect 356974 165560 356980 165572
rect 343324 165532 356980 165560
rect 343324 165520 343330 165532
rect 356974 165520 356980 165532
rect 357032 165560 357038 165572
rect 357434 165560 357440 165572
rect 357032 165532 357440 165560
rect 357032 165520 357038 165532
rect 357434 165520 357440 165532
rect 357492 165520 357498 165572
rect 362402 165520 362408 165572
rect 362460 165560 362466 165572
rect 458358 165560 458364 165572
rect 362460 165532 458364 165560
rect 362460 165520 362466 165532
rect 458358 165520 458364 165532
rect 458416 165520 458422 165572
rect 55030 165452 55036 165504
rect 55088 165492 55094 165504
rect 128354 165492 128360 165504
rect 55088 165464 128360 165492
rect 55088 165452 55094 165464
rect 128354 165452 128360 165464
rect 128412 165452 128418 165504
rect 214650 165452 214656 165504
rect 214708 165492 214714 165504
rect 308398 165492 308404 165504
rect 214708 165464 308404 165492
rect 214708 165452 214714 165464
rect 308398 165452 308404 165464
rect 308456 165452 308462 165504
rect 360930 165452 360936 165504
rect 360988 165492 360994 165504
rect 447318 165492 447324 165504
rect 360988 165464 447324 165492
rect 360988 165452 360994 165464
rect 447318 165452 447324 165464
rect 447376 165452 447382 165504
rect 56502 165384 56508 165436
rect 56560 165424 56566 165436
rect 129734 165424 129740 165436
rect 56560 165396 129740 165424
rect 56560 165384 56566 165396
rect 129734 165384 129740 165396
rect 129792 165384 129798 165436
rect 214558 165384 214564 165436
rect 214616 165424 214622 165436
rect 300854 165424 300860 165436
rect 214616 165396 300860 165424
rect 214616 165384 214622 165396
rect 300854 165384 300860 165396
rect 300912 165384 300918 165436
rect 371970 165384 371976 165436
rect 372028 165424 372034 165436
rect 455414 165424 455420 165436
rect 372028 165396 455420 165424
rect 372028 165384 372034 165396
rect 455414 165384 455420 165396
rect 455472 165384 455478 165436
rect 53282 165316 53288 165368
rect 53340 165356 53346 165368
rect 123478 165356 123484 165368
rect 53340 165328 123484 165356
rect 53340 165316 53346 165328
rect 123478 165316 123484 165328
rect 123536 165316 123542 165368
rect 211890 165316 211896 165368
rect 211948 165356 211954 165368
rect 280154 165356 280160 165368
rect 211948 165328 280160 165356
rect 211948 165316 211954 165328
rect 280154 165316 280160 165328
rect 280212 165316 280218 165368
rect 370682 165316 370688 165368
rect 370740 165356 370746 165368
rect 452654 165356 452660 165368
rect 370740 165328 452660 165356
rect 370740 165316 370746 165328
rect 452654 165316 452660 165328
rect 452712 165316 452718 165368
rect 56318 165248 56324 165300
rect 56376 165288 56382 165300
rect 125870 165288 125876 165300
rect 56376 165260 125876 165288
rect 56376 165248 56382 165260
rect 125870 165248 125876 165260
rect 125928 165248 125934 165300
rect 218974 165248 218980 165300
rect 219032 165288 219038 165300
rect 283374 165288 283380 165300
rect 219032 165260 283380 165288
rect 219032 165248 219038 165260
rect 283374 165248 283380 165260
rect 283432 165248 283438 165300
rect 369118 165248 369124 165300
rect 369176 165288 369182 165300
rect 449894 165288 449900 165300
rect 369176 165260 449900 165288
rect 369176 165248 369182 165260
rect 449894 165248 449900 165260
rect 449952 165248 449958 165300
rect 54938 165180 54944 165232
rect 54996 165220 55002 165232
rect 120902 165220 120908 165232
rect 54996 165192 120908 165220
rect 54996 165180 55002 165192
rect 120902 165180 120908 165192
rect 120960 165180 120966 165232
rect 183278 165180 183284 165232
rect 183336 165220 183342 165232
rect 197354 165220 197360 165232
rect 183336 165192 197360 165220
rect 183336 165180 183342 165192
rect 197354 165180 197360 165192
rect 197412 165180 197418 165232
rect 206370 165180 206376 165232
rect 206428 165220 206434 165232
rect 267918 165220 267924 165232
rect 206428 165192 267924 165220
rect 206428 165180 206434 165192
rect 267918 165180 267924 165192
rect 267976 165180 267982 165232
rect 366450 165180 366456 165232
rect 366508 165220 366514 165232
rect 442994 165220 443000 165232
rect 366508 165192 443000 165220
rect 366508 165180 366514 165192
rect 442994 165180 443000 165192
rect 443052 165180 443058 165232
rect 53190 165112 53196 165164
rect 53248 165152 53254 165164
rect 115934 165152 115940 165164
rect 53248 165124 115940 165152
rect 53248 165112 53254 165124
rect 115934 165112 115940 165124
rect 115992 165112 115998 165164
rect 218790 165112 218796 165164
rect 218848 165152 218854 165164
rect 277394 165152 277400 165164
rect 218848 165124 277400 165152
rect 218848 165112 218854 165124
rect 277394 165112 277400 165124
rect 277452 165112 277458 165164
rect 365070 165112 365076 165164
rect 365128 165152 365134 165164
rect 438026 165152 438032 165164
rect 365128 165124 438032 165152
rect 365128 165112 365134 165124
rect 438026 165112 438032 165124
rect 438084 165112 438090 165164
rect 503254 165112 503260 165164
rect 503312 165152 503318 165164
rect 517606 165152 517612 165164
rect 503312 165124 517612 165152
rect 503312 165112 503318 165124
rect 517606 165112 517612 165124
rect 517664 165112 517670 165164
rect 56042 165044 56048 165096
rect 56100 165084 56106 165096
rect 118326 165084 118332 165096
rect 56100 165056 118332 165084
rect 56100 165044 56106 165056
rect 118326 165044 118332 165056
rect 118384 165044 118390 165096
rect 183370 165044 183376 165096
rect 183428 165084 183434 165096
rect 197446 165084 197452 165096
rect 183428 165056 197452 165084
rect 183428 165044 183434 165056
rect 197446 165044 197452 165056
rect 197504 165044 197510 165096
rect 215938 165044 215944 165096
rect 215996 165084 216002 165096
rect 258074 165084 258080 165096
rect 215996 165056 258080 165084
rect 215996 165044 216002 165056
rect 258074 165044 258080 165056
rect 258132 165044 258138 165096
rect 369210 165044 369216 165096
rect 369268 165084 369274 165096
rect 434714 165084 434720 165096
rect 369268 165056 434720 165084
rect 369268 165044 369274 165056
rect 434714 165044 434720 165056
rect 434772 165044 434778 165096
rect 440234 165044 440240 165096
rect 440292 165084 440298 165096
rect 516594 165084 516600 165096
rect 440292 165056 516600 165084
rect 440292 165044 440298 165056
rect 516594 165044 516600 165056
rect 516652 165044 516658 165096
rect 54846 164976 54852 165028
rect 54904 165016 54910 165028
rect 113542 165016 113548 165028
rect 54904 164988 113548 165016
rect 54904 164976 54910 164988
rect 113542 164976 113548 164988
rect 113600 164976 113606 165028
rect 117314 164976 117320 165028
rect 117372 165016 117378 165028
rect 196802 165016 196808 165028
rect 117372 164988 196808 165016
rect 117372 164976 117378 164988
rect 196802 164976 196808 164988
rect 196860 164976 196866 165028
rect 210510 164976 210516 165028
rect 210568 165016 210574 165028
rect 252554 165016 252560 165028
rect 210568 164988 252560 165016
rect 210568 164976 210574 164988
rect 252554 164976 252560 164988
rect 252612 164976 252618 165028
rect 367830 164976 367836 165028
rect 367888 165016 367894 165028
rect 433334 165016 433340 165028
rect 367888 164988 433340 165016
rect 367888 164976 367894 164988
rect 433334 164976 433340 164988
rect 433392 164976 433398 165028
rect 503346 164976 503352 165028
rect 503404 165016 503410 165028
rect 517882 165016 517888 165028
rect 503404 164988 517888 165016
rect 503404 164976 503410 164988
rect 517882 164976 517888 164988
rect 517940 164976 517946 165028
rect 52178 164908 52184 164960
rect 52236 164948 52242 164960
rect 105722 164948 105728 164960
rect 52236 164920 105728 164948
rect 52236 164908 52242 164920
rect 105722 164908 105728 164920
rect 105780 164908 105786 164960
rect 115934 164908 115940 164960
rect 115992 164948 115998 164960
rect 196710 164948 196716 164960
rect 115992 164920 196716 164948
rect 115992 164908 115998 164920
rect 196710 164908 196716 164920
rect 196768 164908 196774 164960
rect 210418 164908 210424 164960
rect 210476 164948 210482 164960
rect 249794 164948 249800 164960
rect 210476 164920 249800 164948
rect 210476 164908 210482 164920
rect 249794 164908 249800 164920
rect 249852 164908 249858 164960
rect 374730 164908 374736 164960
rect 374788 164948 374794 164960
rect 374788 164920 418154 164948
rect 374788 164908 374794 164920
rect 49602 164840 49608 164892
rect 49660 164880 49666 164892
rect 92474 164880 92480 164892
rect 49660 164852 92480 164880
rect 49660 164840 49666 164852
rect 92474 164840 92480 164852
rect 92532 164840 92538 164892
rect 114554 164840 114560 164892
rect 114612 164880 114618 164892
rect 196618 164880 196624 164892
rect 114612 164852 196624 164880
rect 114612 164840 114618 164852
rect 196618 164840 196624 164852
rect 196676 164840 196682 164892
rect 218882 164840 218888 164892
rect 218940 164880 218946 164892
rect 247678 164880 247684 164892
rect 218940 164852 247684 164880
rect 218940 164840 218946 164852
rect 247678 164840 247684 164852
rect 247736 164840 247742 164892
rect 343450 164840 343456 164892
rect 343508 164880 343514 164892
rect 357618 164880 357624 164892
rect 343508 164852 357624 164880
rect 343508 164840 343514 164852
rect 357618 164840 357624 164852
rect 357676 164840 357682 164892
rect 373258 164840 373264 164892
rect 373316 164880 373322 164892
rect 416038 164880 416044 164892
rect 373316 164852 416044 164880
rect 373316 164840 373322 164852
rect 416038 164840 416044 164852
rect 416096 164840 416102 164892
rect 52086 164772 52092 164824
rect 52144 164812 52150 164824
rect 90266 164812 90272 164824
rect 52144 164784 90272 164812
rect 52144 164772 52150 164784
rect 90266 164772 90272 164784
rect 90324 164772 90330 164824
rect 376110 164772 376116 164824
rect 376168 164812 376174 164824
rect 409874 164812 409880 164824
rect 376168 164784 409880 164812
rect 376168 164772 376174 164784
rect 409874 164772 409880 164784
rect 409932 164772 409938 164824
rect 418126 164812 418154 164920
rect 510522 164908 510528 164960
rect 510580 164948 510586 164960
rect 517514 164948 517520 164960
rect 510580 164920 517520 164948
rect 510580 164908 510586 164920
rect 517514 164908 517520 164920
rect 517572 164908 517578 164960
rect 440326 164812 440332 164824
rect 418126 164784 440332 164812
rect 440326 164772 440332 164784
rect 440384 164772 440390 164824
rect 56410 164704 56416 164756
rect 56468 164744 56474 164756
rect 88334 164744 88340 164756
rect 56468 164716 88340 164744
rect 56468 164704 56474 164716
rect 88334 164704 88340 164716
rect 88392 164704 88398 164756
rect 378870 164704 378876 164756
rect 378928 164744 378934 164756
rect 412634 164744 412640 164756
rect 378928 164716 412640 164744
rect 378928 164704 378934 164716
rect 412634 164704 412640 164716
rect 412692 164704 412698 164756
rect 378962 164636 378968 164688
rect 379020 164676 379026 164688
rect 407114 164676 407120 164688
rect 379020 164648 407120 164676
rect 379020 164636 379026 164648
rect 407114 164636 407120 164648
rect 407172 164636 407178 164688
rect 428918 164568 428924 164620
rect 428976 164608 428982 164620
rect 433518 164608 433524 164620
rect 428976 164580 433524 164608
rect 428976 164568 428982 164580
rect 433518 164568 433524 164580
rect 433576 164568 433582 164620
rect 51626 164228 51632 164280
rect 51684 164268 51690 164280
rect 73798 164268 73804 164280
rect 51684 164240 73804 164268
rect 51684 164228 51690 164240
rect 73798 164228 73804 164240
rect 73856 164228 73862 164280
rect 87598 164228 87604 164280
rect 87656 164268 87662 164280
rect 108298 164268 108304 164280
rect 87656 164240 108304 164268
rect 87656 164228 87662 164240
rect 108298 164228 108304 164240
rect 108356 164228 108362 164280
rect 46566 164160 46572 164212
rect 46624 164200 46630 164212
rect 53282 164200 53288 164212
rect 46624 164172 53288 164200
rect 46624 164160 46630 164172
rect 53282 164160 53288 164172
rect 53340 164160 53346 164212
rect 58618 164160 58624 164212
rect 58676 164200 58682 164212
rect 59998 164200 60004 164212
rect 58676 164172 60004 164200
rect 58676 164160 58682 164172
rect 59998 164160 60004 164172
rect 60056 164160 60062 164212
rect 60090 164160 60096 164212
rect 60148 164200 60154 164212
rect 117866 164200 117872 164212
rect 60148 164172 117872 164200
rect 60148 164160 60154 164172
rect 117866 164160 117872 164172
rect 117924 164160 117930 164212
rect 211982 164160 211988 164212
rect 212040 164200 212046 164212
rect 323026 164200 323032 164212
rect 212040 164172 323032 164200
rect 212040 164160 212046 164172
rect 323026 164160 323032 164172
rect 323084 164160 323090 164212
rect 377398 164160 377404 164212
rect 377456 164200 377462 164212
rect 437750 164200 437756 164212
rect 377456 164172 437756 164200
rect 377456 164160 377462 164172
rect 437750 164160 437756 164172
rect 437808 164160 437814 164212
rect 46474 164092 46480 164144
rect 46532 164132 46538 164144
rect 52178 164132 52184 164144
rect 46532 164104 52184 164132
rect 46532 164092 46538 164104
rect 52178 164092 52184 164104
rect 52236 164092 52242 164144
rect 53374 164092 53380 164144
rect 53432 164132 53438 164144
rect 110966 164132 110972 164144
rect 53432 164104 110972 164132
rect 53432 164092 53438 164104
rect 110966 164092 110972 164104
rect 111024 164092 111030 164144
rect 219618 164092 219624 164144
rect 219676 164132 219682 164144
rect 264974 164132 264980 164144
rect 219676 164104 264980 164132
rect 219676 164092 219682 164104
rect 264974 164092 264980 164104
rect 265032 164092 265038 164144
rect 374546 164092 374552 164144
rect 374604 164132 374610 164144
rect 434714 164132 434720 164144
rect 374604 164104 434720 164132
rect 374604 164092 374610 164104
rect 434714 164092 434720 164104
rect 434772 164092 434778 164144
rect 55858 164024 55864 164076
rect 55916 164064 55922 164076
rect 57514 164064 57520 164076
rect 55916 164036 57520 164064
rect 55916 164024 55922 164036
rect 57514 164024 57520 164036
rect 57572 164024 57578 164076
rect 57698 164024 57704 164076
rect 57756 164064 57762 164076
rect 105170 164064 105176 164076
rect 57756 164036 105176 164064
rect 57756 164024 57762 164036
rect 105170 164024 105176 164036
rect 105228 164024 105234 164076
rect 216582 164024 216588 164076
rect 216640 164064 216646 164076
rect 236086 164064 236092 164076
rect 216640 164036 236092 164064
rect 216640 164024 216646 164036
rect 236086 164024 236092 164036
rect 236144 164024 236150 164076
rect 375006 164024 375012 164076
rect 375064 164064 375070 164076
rect 396166 164064 396172 164076
rect 375064 164036 396172 164064
rect 375064 164024 375070 164036
rect 396166 164024 396172 164036
rect 396224 164024 396230 164076
rect 54386 163956 54392 164008
rect 54444 163996 54450 164008
rect 55030 163996 55036 164008
rect 54444 163968 55036 163996
rect 54444 163956 54450 163968
rect 55030 163956 55036 163968
rect 55088 163996 55094 164008
rect 100846 163996 100852 164008
rect 55088 163968 100852 163996
rect 55088 163956 55094 163968
rect 100846 163956 100852 163968
rect 100904 163956 100910 164008
rect 216214 163956 216220 164008
rect 216272 163996 216278 164008
rect 235994 163996 236000 164008
rect 216272 163968 236000 163996
rect 216272 163956 216278 163968
rect 235994 163956 236000 163968
rect 236052 163956 236058 164008
rect 376202 163956 376208 164008
rect 376260 163996 376266 164008
rect 396074 163996 396080 164008
rect 376260 163968 396080 163996
rect 376260 163956 376266 163968
rect 396074 163956 396080 163968
rect 396132 163956 396138 164008
rect 52822 163888 52828 163940
rect 52880 163928 52886 163940
rect 56502 163928 56508 163940
rect 52880 163900 56508 163928
rect 52880 163888 52886 163900
rect 56502 163888 56508 163900
rect 56560 163928 56566 163940
rect 96614 163928 96620 163940
rect 56560 163900 96620 163928
rect 56560 163888 56566 163900
rect 96614 163888 96620 163900
rect 96672 163888 96678 163940
rect 52914 163820 52920 163872
rect 52972 163860 52978 163872
rect 55122 163860 55128 163872
rect 52972 163832 55128 163860
rect 52972 163820 52978 163832
rect 55122 163820 55128 163832
rect 55180 163860 55186 163872
rect 97994 163860 98000 163872
rect 55180 163832 98000 163860
rect 55180 163820 55186 163832
rect 97994 163820 98000 163832
rect 98052 163820 98058 163872
rect 59998 163752 60004 163804
rect 60056 163792 60062 163804
rect 106366 163792 106372 163804
rect 60056 163764 106372 163792
rect 60056 163752 60062 163764
rect 106366 163752 106372 163764
rect 106424 163752 106430 163804
rect 47854 163684 47860 163736
rect 47912 163724 47918 163736
rect 53374 163724 53380 163736
rect 47912 163696 53380 163724
rect 47912 163684 47918 163696
rect 53374 163684 53380 163696
rect 53432 163724 53438 163736
rect 109678 163724 109684 163736
rect 53432 163696 109684 163724
rect 53432 163684 53438 163696
rect 109678 163684 109684 163696
rect 109736 163684 109742 163736
rect 59354 163616 59360 163668
rect 59412 163656 59418 163668
rect 119062 163656 119068 163668
rect 59412 163628 119068 163656
rect 59412 163616 59418 163628
rect 119062 163616 119068 163628
rect 119120 163616 119126 163668
rect 375190 163616 375196 163668
rect 375248 163656 375254 163668
rect 422294 163656 422300 163668
rect 375248 163628 422300 163656
rect 375248 163616 375254 163628
rect 422294 163616 422300 163628
rect 422352 163616 422358 163668
rect 52178 163548 52184 163600
rect 52236 163588 52242 163600
rect 111886 163588 111892 163600
rect 52236 163560 111892 163588
rect 52236 163548 52242 163560
rect 111886 163548 111892 163560
rect 111944 163548 111950 163600
rect 372154 163548 372160 163600
rect 372212 163588 372218 163600
rect 375006 163588 375012 163600
rect 372212 163560 375012 163588
rect 372212 163548 372218 163560
rect 375006 163548 375012 163560
rect 375064 163588 375070 163600
rect 429286 163588 429292 163600
rect 375064 163560 429292 163588
rect 375064 163548 375070 163560
rect 429286 163548 429292 163560
rect 429344 163548 429350 163600
rect 53282 163480 53288 163532
rect 53340 163520 53346 163532
rect 113174 163520 113180 163532
rect 53340 163492 113180 163520
rect 53340 163480 53346 163492
rect 113174 163480 113180 163492
rect 113232 163480 113238 163532
rect 216674 163480 216680 163532
rect 216732 163520 216738 163532
rect 218882 163520 218888 163532
rect 216732 163492 218888 163520
rect 216732 163480 216738 163492
rect 218882 163480 218888 163492
rect 218940 163520 218946 163532
rect 263778 163520 263784 163532
rect 218940 163492 263784 163520
rect 218940 163480 218946 163492
rect 263778 163480 263784 163492
rect 263836 163480 263842 163532
rect 373166 163480 373172 163532
rect 373224 163520 373230 163532
rect 375098 163520 375104 163532
rect 373224 163492 375104 163520
rect 373224 163480 373230 163492
rect 375098 163480 375104 163492
rect 375156 163520 375162 163532
rect 431954 163520 431960 163532
rect 375156 163492 431960 163520
rect 375156 163480 375162 163492
rect 431954 163480 431960 163492
rect 432012 163480 432018 163532
rect 52362 163412 52368 163464
rect 52420 163452 52426 163464
rect 57238 163452 57244 163464
rect 52420 163424 57244 163452
rect 52420 163412 52426 163424
rect 57238 163412 57244 163424
rect 57296 163452 57302 163464
rect 95234 163452 95240 163464
rect 57296 163424 95240 163452
rect 57296 163412 57302 163424
rect 95234 163412 95240 163424
rect 95292 163412 95298 163464
rect 57514 163344 57520 163396
rect 57572 163384 57578 163396
rect 60090 163384 60096 163396
rect 57572 163356 60096 163384
rect 57572 163344 57578 163356
rect 60090 163344 60096 163356
rect 60148 163344 60154 163396
rect 375190 162868 375196 162920
rect 375248 162908 375254 162920
rect 375248 162880 376248 162908
rect 375248 162868 375254 162880
rect 49142 162800 49148 162852
rect 49200 162840 49206 162852
rect 53466 162840 53472 162852
rect 49200 162812 53472 162840
rect 49200 162800 49206 162812
rect 53466 162800 53472 162812
rect 53524 162800 53530 162852
rect 57054 162800 57060 162852
rect 57112 162840 57118 162852
rect 59170 162840 59176 162852
rect 57112 162812 59176 162840
rect 57112 162800 57118 162812
rect 59170 162800 59176 162812
rect 59228 162800 59234 162852
rect 216030 162800 216036 162852
rect 216088 162840 216094 162852
rect 217134 162840 217140 162852
rect 216088 162812 217140 162840
rect 216088 162800 216094 162812
rect 217134 162800 217140 162812
rect 217192 162800 217198 162852
rect 260834 162840 260840 162852
rect 217244 162812 260840 162840
rect 214466 162664 214472 162716
rect 214524 162704 214530 162716
rect 217244 162704 217272 162812
rect 260834 162800 260840 162812
rect 260892 162800 260898 162852
rect 259546 162772 259552 162784
rect 214524 162676 217272 162704
rect 217336 162744 259552 162772
rect 214524 162664 214530 162676
rect 214834 162596 214840 162648
rect 214892 162636 214898 162648
rect 217336 162636 217364 162744
rect 259546 162732 259552 162744
rect 259604 162732 259610 162784
rect 217870 162664 217876 162716
rect 217928 162704 217934 162716
rect 259454 162704 259460 162716
rect 217928 162676 259460 162704
rect 217928 162664 217934 162676
rect 259454 162664 259460 162676
rect 259512 162664 259518 162716
rect 376220 162648 376248 162880
rect 376294 162800 376300 162852
rect 376352 162840 376358 162852
rect 379790 162840 379796 162852
rect 376352 162812 379796 162840
rect 376352 162800 376358 162812
rect 379790 162800 379796 162812
rect 379848 162800 379854 162852
rect 379974 162800 379980 162852
rect 380032 162840 380038 162852
rect 436094 162840 436100 162852
rect 380032 162812 436100 162840
rect 380032 162800 380038 162812
rect 436094 162800 436100 162812
rect 436152 162800 436158 162852
rect 377214 162732 377220 162784
rect 377272 162772 377278 162784
rect 420914 162772 420920 162784
rect 377272 162744 420920 162772
rect 377272 162732 377278 162744
rect 420914 162732 420920 162744
rect 420972 162732 420978 162784
rect 376294 162664 376300 162716
rect 376352 162704 376358 162716
rect 418614 162704 418620 162716
rect 376352 162676 418620 162704
rect 376352 162664 376358 162676
rect 418614 162664 418620 162676
rect 418672 162664 418678 162716
rect 214892 162608 217364 162636
rect 214892 162596 214898 162608
rect 218514 162596 218520 162648
rect 218572 162636 218578 162648
rect 218974 162636 218980 162648
rect 218572 162608 218980 162636
rect 218572 162596 218578 162608
rect 218974 162596 218980 162608
rect 219032 162636 219038 162648
rect 258074 162636 258080 162648
rect 219032 162608 258080 162636
rect 219032 162596 219038 162608
rect 258074 162596 258080 162608
rect 258132 162596 258138 162648
rect 376202 162596 376208 162648
rect 376260 162596 376266 162648
rect 376386 162596 376392 162648
rect 376444 162636 376450 162648
rect 379146 162636 379152 162648
rect 376444 162608 379152 162636
rect 376444 162596 376450 162608
rect 379146 162596 379152 162608
rect 379204 162636 379210 162648
rect 419534 162636 419540 162648
rect 379204 162608 419540 162636
rect 379204 162596 379210 162608
rect 419534 162596 419540 162608
rect 419592 162596 419598 162648
rect 375926 162528 375932 162580
rect 375984 162568 375990 162580
rect 379974 162568 379980 162580
rect 375984 162540 379980 162568
rect 375984 162528 375990 162540
rect 379974 162528 379980 162540
rect 380032 162528 380038 162580
rect 374914 162460 374920 162512
rect 374972 162500 374978 162512
rect 379146 162500 379152 162512
rect 374972 162472 379152 162500
rect 374972 162460 374978 162472
rect 379146 162460 379152 162472
rect 379204 162460 379210 162512
rect 379790 162256 379796 162308
rect 379848 162296 379854 162308
rect 418154 162296 418160 162308
rect 379848 162268 418160 162296
rect 379848 162256 379854 162268
rect 418154 162256 418160 162268
rect 418212 162256 418218 162308
rect 59170 162188 59176 162240
rect 59228 162228 59234 162240
rect 89898 162228 89904 162240
rect 59228 162200 89904 162228
rect 59228 162188 59234 162200
rect 89898 162188 89904 162200
rect 89956 162188 89962 162240
rect 372246 162188 372252 162240
rect 372304 162228 372310 162240
rect 373718 162228 373724 162240
rect 372304 162200 373724 162228
rect 372304 162188 372310 162200
rect 373718 162188 373724 162200
rect 373776 162228 373782 162240
rect 428918 162228 428924 162240
rect 373776 162200 428924 162228
rect 373776 162188 373782 162200
rect 428918 162188 428924 162200
rect 428976 162188 428982 162240
rect 53466 162120 53472 162172
rect 53524 162160 53530 162172
rect 111150 162160 111156 162172
rect 53524 162132 111156 162160
rect 53524 162120 53530 162132
rect 111150 162120 111156 162132
rect 111208 162120 111214 162172
rect 218606 162120 218612 162172
rect 218664 162160 218670 162172
rect 219526 162160 219532 162172
rect 218664 162132 219532 162160
rect 218664 162120 218670 162132
rect 219526 162120 219532 162132
rect 219584 162160 219590 162172
rect 266354 162160 266360 162172
rect 219584 162132 266360 162160
rect 219584 162120 219590 162132
rect 266354 162120 266360 162132
rect 266412 162120 266418 162172
rect 372338 162120 372344 162172
rect 372396 162160 372402 162172
rect 374822 162160 374828 162172
rect 372396 162132 374828 162160
rect 372396 162120 372402 162132
rect 374822 162120 374828 162132
rect 374880 162160 374886 162172
rect 430574 162160 430580 162172
rect 374880 162132 430580 162160
rect 374880 162120 374886 162132
rect 430574 162120 430580 162132
rect 430632 162120 430638 162172
rect 376570 161916 376576 161968
rect 376628 161956 376634 161968
rect 377214 161956 377220 161968
rect 376628 161928 377220 161956
rect 376628 161916 376634 161928
rect 377214 161916 377220 161928
rect 377272 161916 377278 161968
rect 216214 161508 216220 161560
rect 216272 161548 216278 161560
rect 235258 161548 235264 161560
rect 216272 161520 235264 161548
rect 216272 161508 216278 161520
rect 235258 161508 235264 161520
rect 235316 161508 235322 161560
rect 217134 161440 217140 161492
rect 217192 161480 217198 161492
rect 236638 161480 236644 161492
rect 217192 161452 236644 161480
rect 217192 161440 217198 161452
rect 236638 161440 236644 161452
rect 236696 161440 236702 161492
rect 379146 161440 379152 161492
rect 379204 161480 379210 161492
rect 396718 161480 396724 161492
rect 379204 161452 396724 161480
rect 379204 161440 379210 161452
rect 396718 161440 396724 161452
rect 396776 161440 396782 161492
rect 357526 156612 357532 156664
rect 357584 156652 357590 156664
rect 357710 156652 357716 156664
rect 357584 156624 357716 156652
rect 357584 156612 357590 156624
rect 357710 156612 357716 156624
rect 357768 156612 357774 156664
rect 215754 148996 215760 149048
rect 215812 149036 215818 149048
rect 216490 149036 216496 149048
rect 215812 149008 216496 149036
rect 215812 148996 215818 149008
rect 216490 148996 216496 149008
rect 216548 149036 216554 149048
rect 278774 149036 278780 149048
rect 216548 149008 278780 149036
rect 216548 148996 216554 149008
rect 278774 148996 278780 149008
rect 278832 148996 278838 149048
rect 379698 148996 379704 149048
rect 379756 149036 379762 149048
rect 427906 149036 427912 149048
rect 379756 149008 427912 149036
rect 379756 148996 379762 149008
rect 427906 148996 427912 149008
rect 427964 148996 427970 149048
rect 215018 148928 215024 148980
rect 215076 148968 215082 148980
rect 276106 148968 276112 148980
rect 215076 148940 276112 148968
rect 215076 148928 215082 148940
rect 276106 148928 276112 148940
rect 276164 148928 276170 148980
rect 214926 148860 214932 148912
rect 214984 148900 214990 148912
rect 240134 148900 240140 148912
rect 214984 148872 240140 148900
rect 214984 148860 214990 148872
rect 240134 148860 240140 148872
rect 240192 148860 240198 148912
rect 46658 148656 46664 148708
rect 46716 148696 46722 148708
rect 59906 148696 59912 148708
rect 46716 148668 59912 148696
rect 46716 148656 46722 148668
rect 59906 148656 59912 148668
rect 59964 148696 59970 148708
rect 87598 148696 87604 148708
rect 59964 148668 87604 148696
rect 59964 148656 59970 148668
rect 87598 148656 87604 148668
rect 87656 148656 87662 148708
rect 213178 148656 213184 148708
rect 213236 148696 213242 148708
rect 238754 148696 238760 148708
rect 213236 148668 238760 148696
rect 213236 148656 213242 148668
rect 238754 148656 238760 148668
rect 238812 148656 238818 148708
rect 46750 148588 46756 148640
rect 46808 148628 46814 148640
rect 51994 148628 52000 148640
rect 46808 148600 52000 148628
rect 46808 148588 46814 148600
rect 51994 148588 52000 148600
rect 52052 148628 52058 148640
rect 80054 148628 80060 148640
rect 52052 148600 80060 148628
rect 52052 148588 52058 148600
rect 80054 148588 80060 148600
rect 80112 148588 80118 148640
rect 212258 148588 212264 148640
rect 212316 148628 212322 148640
rect 214558 148628 214564 148640
rect 212316 148600 214564 148628
rect 212316 148588 212322 148600
rect 214558 148588 214564 148600
rect 214616 148628 214622 148640
rect 241514 148628 241520 148640
rect 214616 148600 241520 148628
rect 214616 148588 214622 148600
rect 241514 148588 241520 148600
rect 241572 148588 241578 148640
rect 373902 148588 373908 148640
rect 373960 148628 373966 148640
rect 376018 148628 376024 148640
rect 373960 148600 376024 148628
rect 373960 148588 373966 148600
rect 376018 148588 376024 148600
rect 376076 148628 376082 148640
rect 398834 148628 398840 148640
rect 376076 148600 398840 148628
rect 376076 148588 376082 148600
rect 398834 148588 398840 148600
rect 398892 148588 398898 148640
rect 49234 148520 49240 148572
rect 49292 148560 49298 148572
rect 53190 148560 53196 148572
rect 49292 148532 53196 148560
rect 49292 148520 49298 148532
rect 53190 148520 53196 148532
rect 53248 148560 53254 148572
rect 81434 148560 81440 148572
rect 53248 148532 81440 148560
rect 53248 148520 53254 148532
rect 81434 148520 81440 148532
rect 81492 148520 81498 148572
rect 213362 148520 213368 148572
rect 213420 148560 213426 148572
rect 214650 148560 214656 148572
rect 213420 148532 214656 148560
rect 213420 148520 213426 148532
rect 214650 148520 214656 148532
rect 214708 148560 214714 148572
rect 270494 148560 270500 148572
rect 214708 148532 270500 148560
rect 214708 148520 214714 148532
rect 270494 148520 270500 148532
rect 270552 148520 270558 148572
rect 371694 148520 371700 148572
rect 371752 148560 371758 148572
rect 374638 148560 374644 148572
rect 371752 148532 374644 148560
rect 371752 148520 371758 148532
rect 374638 148520 374644 148532
rect 374696 148560 374702 148572
rect 397454 148560 397460 148572
rect 374696 148532 397460 148560
rect 374696 148520 374702 148532
rect 397454 148520 397460 148532
rect 397512 148520 397518 148572
rect 56226 148452 56232 148504
rect 56284 148492 56290 148504
rect 114554 148492 114560 148504
rect 56284 148464 114560 148492
rect 56284 148452 56290 148464
rect 114554 148452 114560 148464
rect 114612 148452 114618 148504
rect 215846 148452 215852 148504
rect 215904 148492 215910 148504
rect 271874 148492 271880 148504
rect 215904 148464 271880 148492
rect 215904 148452 215910 148464
rect 271874 148452 271880 148464
rect 271932 148452 271938 148504
rect 370958 148452 370964 148504
rect 371016 148492 371022 148504
rect 371970 148492 371976 148504
rect 371016 148464 371976 148492
rect 371016 148452 371022 148464
rect 371970 148452 371976 148464
rect 372028 148492 372034 148504
rect 400214 148492 400220 148504
rect 372028 148464 400220 148492
rect 372028 148452 372034 148464
rect 400214 148452 400220 148464
rect 400272 148452 400278 148504
rect 56318 148384 56324 148436
rect 56376 148424 56382 148436
rect 117314 148424 117320 148436
rect 56376 148396 117320 148424
rect 56376 148384 56382 148396
rect 117314 148384 117320 148396
rect 117372 148384 117378 148436
rect 212902 148384 212908 148436
rect 212960 148424 212966 148436
rect 214834 148424 214840 148436
rect 212960 148396 214840 148424
rect 212960 148384 212966 148396
rect 214834 148384 214840 148396
rect 214892 148424 214898 148436
rect 274634 148424 274640 148436
rect 214892 148396 274640 148424
rect 214892 148384 214898 148396
rect 274634 148384 274640 148396
rect 274692 148384 274698 148436
rect 372706 148384 372712 148436
rect 372764 148424 372770 148436
rect 401594 148424 401600 148436
rect 372764 148396 401600 148424
rect 372764 148384 372770 148396
rect 401594 148384 401600 148396
rect 401652 148384 401658 148436
rect 53006 148316 53012 148368
rect 53064 148356 53070 148368
rect 115934 148356 115940 148368
rect 53064 148328 115940 148356
rect 53064 148316 53070 148328
rect 115934 148316 115940 148328
rect 115992 148316 115998 148368
rect 212074 148316 212080 148368
rect 212132 148356 212138 148368
rect 213730 148356 213736 148368
rect 212132 148328 213736 148356
rect 212132 148316 212138 148328
rect 213730 148316 213736 148328
rect 213788 148356 213794 148368
rect 274726 148356 274732 148368
rect 213788 148328 274732 148356
rect 213788 148316 213794 148328
rect 274726 148316 274732 148328
rect 274784 148316 274790 148368
rect 372430 148316 372436 148368
rect 372488 148356 372494 148368
rect 379974 148356 379980 148368
rect 372488 148328 379980 148356
rect 372488 148316 372494 148328
rect 379974 148316 379980 148328
rect 380032 148356 380038 148368
rect 429194 148356 429200 148368
rect 380032 148328 429200 148356
rect 380032 148316 380038 148328
rect 429194 148316 429200 148328
rect 429252 148316 429258 148368
rect 212994 147704 213000 147756
rect 213052 147744 213058 147756
rect 215018 147744 215024 147756
rect 213052 147716 215024 147744
rect 213052 147704 213058 147716
rect 215018 147704 215024 147716
rect 215076 147704 215082 147756
rect 213638 147636 213644 147688
rect 213696 147676 213702 147688
rect 214926 147676 214932 147688
rect 213696 147648 214932 147676
rect 213696 147636 213702 147648
rect 214926 147636 214932 147648
rect 214984 147636 214990 147688
rect 379422 147636 379428 147688
rect 379480 147676 379486 147688
rect 379698 147676 379704 147688
rect 379480 147648 379704 147676
rect 379480 147636 379486 147648
rect 379698 147636 379704 147648
rect 379756 147636 379762 147688
rect 212166 147568 212172 147620
rect 212224 147608 212230 147620
rect 215846 147608 215852 147620
rect 212224 147580 215852 147608
rect 212224 147568 212230 147580
rect 215846 147568 215852 147580
rect 215904 147568 215910 147620
rect 369670 147568 369676 147620
rect 369728 147608 369734 147620
rect 372706 147608 372712 147620
rect 369728 147580 372712 147608
rect 369728 147568 369734 147580
rect 372706 147568 372712 147580
rect 372764 147608 372770 147620
rect 373258 147608 373264 147620
rect 372764 147580 373264 147608
rect 372764 147568 372770 147580
rect 373258 147568 373264 147580
rect 373316 147568 373322 147620
rect 210786 147500 210792 147552
rect 210844 147540 210850 147552
rect 213178 147540 213184 147552
rect 210844 147512 213184 147540
rect 210844 147500 210850 147512
rect 213178 147500 213184 147512
rect 213236 147500 213242 147552
rect 379256 146288 379744 146316
rect 47762 146208 47768 146260
rect 47820 146248 47826 146260
rect 51718 146248 51724 146260
rect 47820 146220 51724 146248
rect 47820 146208 47826 146220
rect 51718 146208 51724 146220
rect 51776 146208 51782 146260
rect 54754 146208 54760 146260
rect 54812 146248 54818 146260
rect 59722 146248 59728 146260
rect 54812 146220 59728 146248
rect 54812 146208 54818 146220
rect 59722 146208 59728 146220
rect 59780 146248 59786 146260
rect 99374 146248 99380 146260
rect 59780 146220 99380 146248
rect 59780 146208 59786 146220
rect 99374 146208 99380 146220
rect 99432 146208 99438 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197538 146248 197544 146260
rect 179104 146220 197544 146248
rect 179104 146208 179110 146220
rect 197538 146208 197544 146220
rect 197596 146208 197602 146260
rect 235258 146208 235264 146260
rect 235316 146248 235322 146260
rect 255314 146248 255320 146260
rect 235316 146220 255320 146248
rect 235316 146208 235322 146220
rect 255314 146208 255320 146220
rect 255372 146208 255378 146260
rect 276014 146208 276020 146260
rect 276072 146248 276078 146260
rect 356882 146248 356888 146260
rect 276072 146220 356888 146248
rect 276072 146208 276078 146220
rect 356882 146208 356888 146220
rect 356940 146208 356946 146260
rect 374730 146208 374736 146260
rect 374788 146248 374794 146260
rect 375558 146248 375564 146260
rect 374788 146220 375564 146248
rect 374788 146208 374794 146220
rect 375558 146208 375564 146220
rect 375616 146208 375622 146260
rect 376478 146208 376484 146260
rect 376536 146248 376542 146260
rect 377490 146248 377496 146260
rect 376536 146220 377496 146248
rect 376536 146208 376542 146220
rect 377490 146208 377496 146220
rect 377548 146208 377554 146260
rect 57054 146140 57060 146192
rect 57112 146180 57118 146192
rect 57974 146180 57980 146192
rect 57112 146152 57980 146180
rect 57112 146140 57118 146152
rect 57974 146140 57980 146152
rect 58032 146140 58038 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197630 146180 197636 146192
rect 179748 146152 197636 146180
rect 179748 146140 179754 146152
rect 197630 146140 197636 146152
rect 197688 146140 197694 146192
rect 219250 146140 219256 146192
rect 219308 146180 219314 146192
rect 219308 146152 229094 146180
rect 219308 146140 219314 146152
rect 52914 146072 52920 146124
rect 52972 146112 52978 146124
rect 53834 146112 53840 146124
rect 52972 146084 53840 146112
rect 52972 146072 52978 146084
rect 53834 146072 53840 146084
rect 53892 146112 53898 146124
rect 86954 146112 86960 146124
rect 53892 146084 86960 146112
rect 53892 146072 53898 146084
rect 86954 146072 86960 146084
rect 87012 146072 87018 146124
rect 229066 146112 229094 146152
rect 236638 146140 236644 146192
rect 236696 146180 236702 146192
rect 256694 146180 256700 146192
rect 236696 146152 256700 146180
rect 236696 146140 236702 146152
rect 256694 146140 256700 146152
rect 256752 146140 256758 146192
rect 338482 146140 338488 146192
rect 338540 146180 338546 146192
rect 360194 146180 360200 146192
rect 338540 146152 360200 146180
rect 338540 146140 338546 146152
rect 360194 146140 360200 146152
rect 360252 146140 360258 146192
rect 374454 146140 374460 146192
rect 374512 146180 374518 146192
rect 375190 146180 375196 146192
rect 374512 146152 375196 146180
rect 374512 146140 374518 146152
rect 375190 146140 375196 146152
rect 375248 146140 375254 146192
rect 375926 146140 375932 146192
rect 375984 146180 375990 146192
rect 378962 146180 378968 146192
rect 375984 146152 378968 146180
rect 375984 146140 375990 146152
rect 378962 146140 378968 146152
rect 379020 146180 379026 146192
rect 379256 146180 379284 146288
rect 379330 146208 379336 146260
rect 379388 146248 379394 146260
rect 379606 146248 379612 146260
rect 379388 146220 379612 146248
rect 379388 146208 379394 146220
rect 379606 146208 379612 146220
rect 379664 146208 379670 146260
rect 379716 146248 379744 146288
rect 404354 146248 404360 146260
rect 379716 146220 404360 146248
rect 404354 146208 404360 146220
rect 404412 146208 404418 146260
rect 379020 146152 379284 146180
rect 379020 146140 379026 146152
rect 251174 146112 251180 146124
rect 229066 146084 251180 146112
rect 251174 146072 251180 146084
rect 251232 146072 251238 146124
rect 340230 146072 340236 146124
rect 340288 146112 340294 146124
rect 357710 146112 357716 146124
rect 340288 146084 357716 146112
rect 340288 146072 340294 146084
rect 357710 146072 357716 146084
rect 357768 146072 357774 146124
rect 379624 146112 379652 146208
rect 396718 146140 396724 146192
rect 396776 146180 396782 146192
rect 416774 146180 416780 146192
rect 396776 146152 416780 146180
rect 396776 146140 396782 146152
rect 416774 146140 416780 146152
rect 416832 146140 416838 146192
rect 500218 146140 500224 146192
rect 500276 146180 500282 146192
rect 517514 146180 517520 146192
rect 500276 146152 517520 146180
rect 500276 146140 500282 146152
rect 517514 146140 517520 146152
rect 517572 146180 517578 146192
rect 517790 146180 517796 146192
rect 517572 146152 517796 146180
rect 517572 146140 517578 146152
rect 517790 146140 517796 146152
rect 517848 146140 517854 146192
rect 412726 146112 412732 146124
rect 379624 146084 412732 146112
rect 412726 146072 412732 146084
rect 412784 146072 412790 146124
rect 498654 146072 498660 146124
rect 498712 146112 498718 146124
rect 517698 146112 517704 146124
rect 498712 146084 517704 146112
rect 498712 146072 498718 146084
rect 517698 146072 517704 146084
rect 517756 146072 517762 146124
rect 57974 146004 57980 146056
rect 58032 146044 58038 146056
rect 91094 146044 91100 146056
rect 58032 146016 91100 146044
rect 58032 146004 58038 146016
rect 91094 146004 91100 146016
rect 91152 146004 91158 146056
rect 219066 146004 219072 146056
rect 219124 146044 219130 146056
rect 251266 146044 251272 146056
rect 219124 146016 251272 146044
rect 219124 146004 219130 146016
rect 251266 146004 251272 146016
rect 251324 146004 251330 146056
rect 378594 146004 378600 146056
rect 378652 146044 378658 146056
rect 411254 146044 411260 146056
rect 378652 146016 411260 146044
rect 378652 146004 378658 146016
rect 411254 146004 411260 146016
rect 411312 146004 411318 146056
rect 56134 145936 56140 145988
rect 56192 145976 56198 145988
rect 88426 145976 88432 145988
rect 56192 145948 88432 145976
rect 56192 145936 56198 145948
rect 88426 145936 88432 145948
rect 88484 145936 88490 145988
rect 217870 145936 217876 145988
rect 217928 145976 217934 145988
rect 249794 145976 249800 145988
rect 217928 145948 249800 145976
rect 217928 145936 217934 145948
rect 249794 145936 249800 145948
rect 249852 145936 249858 145988
rect 377858 145936 377864 145988
rect 377916 145976 377922 145988
rect 379238 145976 379244 145988
rect 377916 145948 379244 145976
rect 377916 145936 377922 145948
rect 379238 145936 379244 145948
rect 379296 145976 379302 145988
rect 409966 145976 409972 145988
rect 379296 145948 409972 145976
rect 379296 145936 379302 145948
rect 409966 145936 409972 145948
rect 410024 145936 410030 145988
rect 54938 145868 54944 145920
rect 54996 145908 55002 145920
rect 85574 145908 85580 145920
rect 54996 145880 85580 145908
rect 54996 145868 55002 145880
rect 85574 145868 85580 145880
rect 85632 145868 85638 145920
rect 219342 145868 219348 145920
rect 219400 145908 219406 145920
rect 248414 145908 248420 145920
rect 219400 145880 248420 145908
rect 219400 145868 219406 145880
rect 248414 145868 248420 145880
rect 248472 145868 248478 145920
rect 377490 145868 377496 145920
rect 377548 145908 377554 145920
rect 407206 145908 407212 145920
rect 377548 145880 407212 145908
rect 377548 145868 377554 145880
rect 407206 145868 407212 145880
rect 407264 145868 407270 145920
rect 46382 145800 46388 145852
rect 46440 145840 46446 145852
rect 52362 145840 52368 145852
rect 46440 145812 52368 145840
rect 46440 145800 46446 145812
rect 52362 145800 52368 145812
rect 52420 145840 52426 145852
rect 77294 145840 77300 145852
rect 52420 145812 77300 145840
rect 52420 145800 52426 145812
rect 77294 145800 77300 145812
rect 77352 145800 77358 145852
rect 215110 145800 215116 145852
rect 215168 145840 215174 145852
rect 244274 145840 244280 145852
rect 215168 145812 244280 145840
rect 215168 145800 215174 145812
rect 244274 145800 244280 145812
rect 244332 145800 244338 145852
rect 375650 145800 375656 145852
rect 375708 145840 375714 145852
rect 405734 145840 405740 145852
rect 375708 145812 405740 145840
rect 375708 145800 375714 145812
rect 405734 145800 405740 145812
rect 405792 145800 405798 145852
rect 51718 145732 51724 145784
rect 51776 145772 51782 145784
rect 78674 145772 78680 145784
rect 51776 145744 78680 145772
rect 51776 145732 51782 145744
rect 78674 145732 78680 145744
rect 78732 145732 78738 145784
rect 217962 145732 217968 145784
rect 218020 145772 218026 145784
rect 247034 145772 247040 145784
rect 218020 145744 247040 145772
rect 218020 145732 218026 145744
rect 247034 145732 247040 145744
rect 247092 145732 247098 145784
rect 375190 145732 375196 145784
rect 375248 145772 375254 145784
rect 403066 145772 403072 145784
rect 375248 145744 403072 145772
rect 375248 145732 375254 145744
rect 403066 145732 403072 145744
rect 403124 145732 403130 145784
rect 49326 145664 49332 145716
rect 49384 145704 49390 145716
rect 54570 145704 54576 145716
rect 49384 145676 54576 145704
rect 49384 145664 49390 145676
rect 54570 145664 54576 145676
rect 54628 145704 54634 145716
rect 82814 145704 82820 145716
rect 54628 145676 82820 145704
rect 54628 145664 54634 145676
rect 82814 145664 82820 145676
rect 82872 145664 82878 145716
rect 216122 145664 216128 145716
rect 216180 145704 216186 145716
rect 219342 145704 219348 145716
rect 216180 145676 219348 145704
rect 216180 145664 216186 145676
rect 219342 145664 219348 145676
rect 219400 145664 219406 145716
rect 219434 145664 219440 145716
rect 219492 145704 219498 145716
rect 244366 145704 244372 145716
rect 219492 145676 244372 145704
rect 219492 145664 219498 145676
rect 244366 145664 244372 145676
rect 244424 145664 244430 145716
rect 375558 145664 375564 145716
rect 375616 145704 375622 145716
rect 402974 145704 402980 145716
rect 375616 145676 402980 145704
rect 375616 145664 375622 145676
rect 402974 145664 402980 145676
rect 403032 145664 403038 145716
rect 56410 145596 56416 145648
rect 56468 145636 56474 145648
rect 84194 145636 84200 145648
rect 56468 145608 84200 145636
rect 56468 145596 56474 145608
rect 84194 145596 84200 145608
rect 84252 145596 84258 145648
rect 215662 145596 215668 145648
rect 215720 145636 215726 145648
rect 216306 145636 216312 145648
rect 215720 145608 216312 145636
rect 215720 145596 215726 145608
rect 216306 145596 216312 145608
rect 216364 145596 216370 145648
rect 216582 145596 216588 145648
rect 216640 145636 216646 145648
rect 242894 145636 242900 145648
rect 216640 145608 242900 145636
rect 216640 145596 216646 145608
rect 242894 145596 242900 145608
rect 242952 145596 242958 145648
rect 378778 145596 378784 145648
rect 378836 145636 378842 145648
rect 408494 145636 408500 145648
rect 378836 145608 408500 145636
rect 378836 145596 378842 145608
rect 408494 145596 408500 145608
rect 408552 145596 408558 145648
rect 517514 145596 517520 145648
rect 517572 145636 517578 145648
rect 580258 145636 580264 145648
rect 517572 145608 580264 145636
rect 517572 145596 517578 145608
rect 580258 145596 580264 145608
rect 580316 145596 580322 145648
rect 58618 145528 58624 145580
rect 58676 145568 58682 145580
rect 91186 145568 91192 145580
rect 58676 145540 91192 145568
rect 58676 145528 58682 145540
rect 91186 145528 91192 145540
rect 91244 145528 91250 145580
rect 191282 145528 191288 145580
rect 191340 145568 191346 145580
rect 202138 145568 202144 145580
rect 191340 145540 202144 145568
rect 191340 145528 191346 145540
rect 202138 145528 202144 145540
rect 202196 145568 202202 145580
rect 204898 145568 204904 145580
rect 202196 145540 204904 145568
rect 202196 145528 202202 145540
rect 204898 145528 204904 145540
rect 204956 145528 204962 145580
rect 217042 145528 217048 145580
rect 217100 145568 217106 145580
rect 219066 145568 219072 145580
rect 217100 145540 219072 145568
rect 217100 145528 217106 145540
rect 219066 145528 219072 145540
rect 219124 145528 219130 145580
rect 219342 145528 219348 145580
rect 219400 145568 219406 145580
rect 245654 145568 245660 145580
rect 219400 145540 245660 145568
rect 219400 145528 219406 145540
rect 245654 145528 245660 145540
rect 245712 145528 245718 145580
rect 280062 145528 280068 145580
rect 280120 145568 280126 145580
rect 307662 145568 307668 145580
rect 280120 145540 307668 145568
rect 280120 145528 280126 145540
rect 307662 145528 307668 145540
rect 307720 145528 307726 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358078 145568 358084 145580
rect 351696 145540 358084 145568
rect 351696 145528 351702 145540
rect 358078 145528 358084 145540
rect 358136 145568 358142 145580
rect 358722 145568 358728 145580
rect 358136 145540 358728 145568
rect 358136 145528 358142 145540
rect 358722 145528 358728 145540
rect 358780 145568 358786 145580
rect 510522 145568 510528 145580
rect 358780 145540 510528 145568
rect 358780 145528 358786 145540
rect 510522 145528 510528 145540
rect 510580 145528 510586 145580
rect 517698 145528 517704 145580
rect 517756 145568 517762 145580
rect 580350 145568 580356 145580
rect 517756 145540 580356 145568
rect 517756 145528 517762 145540
rect 580350 145528 580356 145540
rect 580408 145528 580414 145580
rect 58802 145460 58808 145512
rect 58860 145500 58866 145512
rect 84286 145500 84292 145512
rect 58860 145472 84292 145500
rect 58860 145460 58866 145472
rect 84286 145460 84292 145472
rect 84344 145460 84350 145512
rect 218514 145460 218520 145512
rect 218572 145500 218578 145512
rect 236086 145500 236092 145512
rect 218572 145472 236092 145500
rect 218572 145460 218578 145472
rect 236086 145460 236092 145472
rect 236144 145460 236150 145512
rect 378962 145460 378968 145512
rect 379020 145500 379026 145512
rect 396166 145500 396172 145512
rect 379020 145472 396172 145500
rect 379020 145460 379026 145472
rect 396166 145460 396172 145472
rect 396224 145460 396230 145512
rect 47670 145392 47676 145444
rect 47728 145432 47734 145444
rect 54662 145432 54668 145444
rect 47728 145404 54668 145432
rect 47728 145392 47734 145404
rect 54662 145392 54668 145404
rect 54720 145432 54726 145444
rect 76006 145432 76012 145444
rect 54720 145404 76012 145432
rect 54720 145392 54726 145404
rect 76006 145392 76012 145404
rect 76064 145392 76070 145444
rect 219066 145392 219072 145444
rect 219124 145432 219130 145444
rect 235994 145432 236000 145444
rect 219124 145404 236000 145432
rect 219124 145392 219130 145404
rect 235994 145392 236000 145404
rect 236052 145392 236058 145444
rect 378870 145392 378876 145444
rect 378928 145432 378934 145444
rect 396074 145432 396080 145444
rect 378928 145404 396080 145432
rect 378928 145392 378934 145404
rect 396074 145392 396080 145404
rect 396132 145392 396138 145444
rect 47486 145324 47492 145376
rect 47544 145364 47550 145376
rect 54846 145364 54852 145376
rect 47544 145336 54852 145364
rect 47544 145324 47550 145336
rect 54846 145324 54852 145336
rect 54904 145364 54910 145376
rect 75914 145364 75920 145376
rect 54904 145336 75920 145364
rect 54904 145324 54910 145336
rect 75914 145324 75920 145336
rect 75972 145324 75978 145376
rect 216306 145324 216312 145376
rect 216364 145364 216370 145376
rect 219434 145364 219440 145376
rect 216364 145336 219440 145364
rect 216364 145324 216370 145336
rect 219434 145324 219440 145336
rect 219492 145324 219498 145376
rect 219710 145324 219716 145376
rect 219768 145364 219774 145376
rect 253934 145364 253940 145376
rect 219768 145336 253940 145364
rect 219768 145324 219774 145336
rect 253934 145324 253940 145336
rect 253992 145324 253998 145376
rect 379882 145324 379888 145376
rect 379940 145364 379946 145376
rect 414014 145364 414020 145376
rect 379940 145336 414020 145364
rect 379940 145324 379946 145336
rect 414014 145324 414020 145336
rect 414072 145324 414078 145376
rect 59630 145256 59636 145308
rect 59688 145296 59694 145308
rect 93854 145296 93860 145308
rect 59688 145268 93860 145296
rect 59688 145256 59694 145268
rect 93854 145256 93860 145268
rect 93912 145256 93918 145308
rect 219802 145256 219808 145308
rect 219860 145296 219866 145308
rect 252554 145296 252560 145308
rect 219860 145268 252560 145296
rect 219860 145256 219866 145268
rect 252554 145256 252560 145268
rect 252612 145256 252618 145308
rect 378042 145256 378048 145308
rect 378100 145296 378106 145308
rect 411346 145296 411352 145308
rect 378100 145268 411352 145296
rect 378100 145256 378106 145268
rect 411346 145256 411352 145268
rect 411404 145256 411410 145308
rect 216766 145120 216772 145172
rect 216824 145160 216830 145172
rect 217870 145160 217876 145172
rect 216824 145132 217876 145160
rect 216824 145120 216830 145132
rect 217870 145120 217876 145132
rect 217928 145120 217934 145172
rect 218606 145052 218612 145104
rect 218664 145092 218670 145104
rect 219250 145092 219256 145104
rect 218664 145064 219256 145092
rect 218664 145052 218670 145064
rect 219250 145052 219256 145064
rect 219308 145052 219314 145104
rect 216398 144916 216404 144968
rect 216456 144956 216462 144968
rect 217962 144956 217968 144968
rect 216456 144928 217968 144956
rect 216456 144916 216462 144928
rect 217962 144916 217968 144928
rect 218020 144916 218026 144968
rect 219250 144916 219256 144968
rect 219308 144956 219314 144968
rect 219802 144956 219808 144968
rect 219308 144928 219808 144956
rect 219308 144916 219314 144928
rect 219802 144916 219808 144928
rect 219860 144916 219866 144968
rect 54478 144848 54484 144900
rect 54536 144888 54542 144900
rect 55858 144888 55864 144900
rect 54536 144860 55864 144888
rect 54536 144848 54542 144860
rect 55858 144848 55864 144860
rect 55916 144888 55922 144900
rect 56410 144888 56416 144900
rect 55916 144860 56416 144888
rect 55916 144848 55922 144860
rect 56410 144848 56416 144860
rect 56468 144848 56474 144900
rect 209314 144848 209320 144900
rect 209372 144888 209378 144900
rect 213270 144888 213276 144900
rect 209372 144860 213276 144888
rect 209372 144848 209378 144860
rect 213270 144848 213276 144860
rect 213328 144848 213334 144900
rect 213546 144848 213552 144900
rect 213604 144888 213610 144900
rect 216030 144888 216036 144900
rect 213604 144860 216036 144888
rect 213604 144848 213610 144860
rect 216030 144848 216036 144860
rect 216088 144888 216094 144900
rect 216582 144888 216588 144900
rect 216088 144860 216588 144888
rect 216088 144848 216094 144860
rect 216582 144848 216588 144860
rect 216640 144848 216646 144900
rect 307662 144848 307668 144900
rect 307720 144888 307726 144900
rect 356606 144888 356612 144900
rect 307720 144860 356612 144888
rect 307720 144848 307726 144860
rect 356606 144848 356612 144860
rect 356664 144848 356670 144900
rect 374362 144848 374368 144900
rect 374420 144888 374426 144900
rect 378778 144888 378784 144900
rect 374420 144860 378784 144888
rect 374420 144848 374426 144860
rect 378778 144848 378784 144860
rect 378836 144848 378842 144900
rect 51810 144780 51816 144832
rect 51868 144820 51874 144832
rect 58802 144820 58808 144832
rect 51868 144792 58808 144820
rect 51868 144780 51874 144792
rect 58802 144780 58808 144792
rect 58860 144780 58866 144832
rect 213454 144780 213460 144832
rect 213512 144820 213518 144832
rect 214926 144820 214932 144832
rect 213512 144792 214932 144820
rect 213512 144780 213518 144792
rect 214926 144780 214932 144792
rect 214984 144780 214990 144832
rect 51902 144712 51908 144764
rect 51960 144752 51966 144764
rect 58618 144752 58624 144764
rect 51960 144724 58624 144752
rect 51960 144712 51966 144724
rect 58618 144712 58624 144724
rect 58676 144712 58682 144764
rect 213086 144712 213092 144764
rect 213144 144752 213150 144764
rect 218790 144752 218796 144764
rect 213144 144724 218796 144752
rect 213144 144712 213150 144724
rect 218790 144712 218796 144724
rect 218848 144752 218854 144764
rect 219342 144752 219348 144764
rect 218848 144724 219348 144752
rect 218848 144712 218854 144724
rect 219342 144712 219348 144724
rect 219400 144712 219406 144764
rect 53098 144644 53104 144696
rect 53156 144684 53162 144696
rect 58894 144684 58900 144696
rect 53156 144656 58900 144684
rect 53156 144644 53162 144656
rect 58894 144644 58900 144656
rect 58952 144644 58958 144696
rect 50430 144576 50436 144628
rect 50488 144616 50494 144628
rect 58710 144616 58716 144628
rect 50488 144588 58716 144616
rect 50488 144576 50494 144588
rect 58710 144576 58716 144588
rect 58768 144576 58774 144628
rect 219894 143284 219900 143336
rect 219952 143324 219958 143336
rect 220078 143324 220084 143336
rect 219952 143296 220084 143324
rect 219952 143284 219958 143296
rect 220078 143284 220084 143296
rect 220136 143284 220142 143336
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 21358 97968 21364 97980
rect 3292 97940 21364 97968
rect 3292 97928 3298 97940
rect 21358 97928 21364 97940
rect 21416 97928 21422 97980
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 202230 70320 202236 70372
rect 202288 70360 202294 70372
rect 216674 70360 216680 70372
rect 202288 70332 216680 70360
rect 202288 70320 202294 70332
rect 216674 70320 216680 70332
rect 216732 70320 216738 70372
rect 363782 70320 363788 70372
rect 363840 70360 363846 70372
rect 376938 70360 376944 70372
rect 363840 70332 376944 70360
rect 363840 70320 363846 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 358078 68416 358084 68468
rect 358136 68456 358142 68468
rect 358722 68456 358728 68468
rect 358136 68428 358728 68456
rect 358136 68416 358142 68428
rect 358722 68416 358728 68428
rect 358780 68456 358786 68468
rect 358780 68428 364334 68456
rect 358780 68416 358786 68428
rect 364306 68320 364334 68428
rect 376938 68320 376944 68332
rect 364306 68292 376944 68320
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 204898 67600 204904 67652
rect 204956 67640 204962 67652
rect 216674 67640 216680 67652
rect 204956 67612 216680 67640
rect 204956 67600 204962 67612
rect 216674 67600 216680 67612
rect 216732 67600 216738 67652
rect 218330 61072 218336 61124
rect 218388 61112 218394 61124
rect 218606 61112 218612 61124
rect 218388 61084 218612 61112
rect 218388 61072 218394 61084
rect 218606 61072 218612 61084
rect 218664 61072 218670 61124
rect 378962 59712 378968 59764
rect 379020 59752 379026 59764
rect 396074 59752 396080 59764
rect 379020 59724 396080 59752
rect 379020 59712 379026 59724
rect 396074 59712 396080 59724
rect 396132 59712 396138 59764
rect 54662 59644 54668 59696
rect 54720 59684 54726 59696
rect 77110 59684 77116 59696
rect 54720 59656 77116 59684
rect 54720 59644 54726 59656
rect 77110 59644 77116 59656
rect 77168 59644 77174 59696
rect 218514 59644 218520 59696
rect 218572 59684 218578 59696
rect 237098 59684 237104 59696
rect 218572 59656 237104 59684
rect 218572 59644 218578 59656
rect 237098 59644 237104 59656
rect 237156 59644 237162 59696
rect 378870 59644 378876 59696
rect 378928 59684 378934 59696
rect 397086 59684 397092 59696
rect 378928 59656 397092 59684
rect 378928 59644 378934 59656
rect 397086 59644 397092 59656
rect 397144 59644 397150 59696
rect 55030 59576 55036 59628
rect 55088 59616 55094 59628
rect 100754 59616 100760 59628
rect 55088 59588 100760 59616
rect 55088 59576 55094 59588
rect 100754 59576 100760 59588
rect 100812 59576 100818 59628
rect 216214 59576 216220 59628
rect 216272 59616 216278 59628
rect 255866 59616 255872 59628
rect 216272 59588 255872 59616
rect 216272 59576 216278 59588
rect 255866 59576 255872 59588
rect 255924 59576 255930 59628
rect 379146 59576 379152 59628
rect 379204 59616 379210 59628
rect 416958 59616 416964 59628
rect 379204 59588 416964 59616
rect 379204 59576 379210 59588
rect 416958 59576 416964 59588
rect 417016 59576 417022 59628
rect 54570 59508 54576 59560
rect 54628 59548 54634 59560
rect 83090 59548 83096 59560
rect 54628 59520 83096 59548
rect 54628 59508 54634 59520
rect 83090 59508 83096 59520
rect 83148 59508 83154 59560
rect 217134 59508 217140 59560
rect 217192 59548 217198 59560
rect 256970 59548 256976 59560
rect 217192 59520 256976 59548
rect 217192 59508 217198 59520
rect 256970 59508 256976 59520
rect 257028 59508 257034 59560
rect 376202 59508 376208 59560
rect 376260 59548 376266 59560
rect 422846 59548 422852 59560
rect 376260 59520 422852 59548
rect 376260 59508 376266 59520
rect 422846 59508 422852 59520
rect 422904 59508 422910 59560
rect 54754 59440 54760 59492
rect 54812 59480 54818 59492
rect 99466 59480 99472 59492
rect 54812 59452 99472 59480
rect 54812 59440 54818 59452
rect 99466 59440 99472 59452
rect 99524 59440 99530 59492
rect 218882 59440 218888 59492
rect 218940 59480 218946 59492
rect 263870 59480 263876 59492
rect 218940 59452 263876 59480
rect 218940 59440 218946 59452
rect 263870 59440 263876 59452
rect 263928 59440 263934 59492
rect 377214 59440 377220 59492
rect 377272 59480 377278 59492
rect 423950 59480 423956 59492
rect 377272 59452 423956 59480
rect 377272 59440 377278 59452
rect 423950 59440 423956 59452
rect 424008 59440 424014 59492
rect 48222 59372 48228 59424
rect 48280 59412 48286 59424
rect 105906 59412 105912 59424
rect 48280 59384 105912 59412
rect 48280 59372 48286 59384
rect 105906 59372 105912 59384
rect 105964 59372 105970 59424
rect 215846 59372 215852 59424
rect 215904 59412 215910 59424
rect 262858 59412 262864 59424
rect 215904 59384 262864 59412
rect 215904 59372 215910 59384
rect 262858 59372 262864 59384
rect 262916 59372 262922 59424
rect 358170 59372 358176 59424
rect 358228 59412 358234 59424
rect 416038 59412 416044 59424
rect 358228 59384 416044 59412
rect 358228 59372 358234 59384
rect 416038 59372 416044 59384
rect 416096 59372 416102 59424
rect 55858 59304 55864 59356
rect 55916 59344 55922 59356
rect 84194 59344 84200 59356
rect 55916 59316 84200 59344
rect 55916 59304 55922 59316
rect 84194 59304 84200 59316
rect 84252 59304 84258 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 358078 59344 358084 59356
rect 218020 59316 358084 59344
rect 218020 59304 218026 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 375190 59304 375196 59356
rect 375248 59344 375254 59356
rect 403066 59344 403072 59356
rect 375248 59316 403072 59344
rect 375248 59304 375254 59316
rect 403066 59304 403072 59316
rect 403124 59304 403130 59356
rect 59170 59236 59176 59288
rect 59228 59276 59234 59288
rect 89990 59276 89996 59288
rect 59228 59248 89996 59276
rect 59228 59236 59234 59248
rect 89990 59236 89996 59248
rect 90048 59236 90054 59288
rect 218974 59236 218980 59288
rect 219032 59276 219038 59288
rect 258074 59276 258080 59288
rect 219032 59248 258080 59276
rect 219032 59236 219038 59248
rect 258074 59236 258080 59248
rect 258132 59236 258138 59288
rect 379790 59236 379796 59288
rect 379848 59276 379854 59288
rect 418154 59276 418160 59288
rect 379848 59248 418160 59276
rect 379848 59236 379854 59248
rect 418154 59236 418160 59248
rect 418212 59236 418218 59288
rect 59814 59168 59820 59220
rect 59872 59208 59878 59220
rect 94498 59208 94504 59220
rect 59872 59180 94504 59208
rect 59872 59168 59878 59180
rect 94498 59168 94504 59180
rect 94556 59168 94562 59220
rect 214742 59168 214748 59220
rect 214800 59208 214806 59220
rect 260650 59208 260656 59220
rect 214800 59180 260656 59208
rect 214800 59168 214806 59180
rect 260650 59168 260656 59180
rect 260708 59168 260714 59220
rect 374730 59168 374736 59220
rect 374788 59208 374794 59220
rect 404170 59208 404176 59220
rect 374788 59180 404176 59208
rect 374788 59168 374794 59180
rect 404170 59168 404176 59180
rect 404228 59168 404234 59220
rect 57238 59100 57244 59152
rect 57296 59140 57302 59152
rect 95878 59140 95884 59152
rect 57296 59112 95884 59140
rect 57296 59100 57302 59112
rect 95878 59100 95884 59112
rect 95936 59100 95942 59152
rect 214466 59100 214472 59152
rect 214524 59140 214530 59152
rect 261754 59140 261760 59152
rect 214524 59112 261760 59140
rect 214524 59100 214530 59112
rect 261754 59100 261760 59112
rect 261812 59100 261818 59152
rect 279234 59100 279240 59152
rect 279292 59140 279298 59152
rect 356606 59140 356612 59152
rect 279292 59112 356612 59140
rect 279292 59100 279298 59112
rect 356606 59100 356612 59112
rect 356664 59100 356670 59152
rect 376110 59100 376116 59152
rect 376168 59140 376174 59152
rect 419350 59140 419356 59152
rect 376168 59112 419356 59140
rect 376168 59100 376174 59112
rect 419350 59100 419356 59112
rect 419408 59100 419414 59152
rect 56502 59032 56508 59084
rect 56560 59072 56566 59084
rect 96982 59072 96988 59084
rect 56560 59044 96988 59072
rect 56560 59032 56566 59044
rect 96982 59032 96988 59044
rect 97040 59032 97046 59084
rect 212442 59032 212448 59084
rect 212500 59072 212506 59084
rect 290918 59072 290924 59084
rect 212500 59044 290924 59072
rect 212500 59032 212506 59044
rect 290918 59032 290924 59044
rect 290976 59032 290982 59084
rect 376386 59032 376392 59084
rect 376444 59072 376450 59084
rect 420638 59072 420644 59084
rect 376444 59044 420644 59072
rect 376444 59032 376450 59044
rect 420638 59032 420644 59044
rect 420696 59032 420702 59084
rect 56134 58964 56140 59016
rect 56192 59004 56198 59016
rect 102778 59004 102784 59016
rect 56192 58976 102784 59004
rect 56192 58964 56198 58976
rect 102778 58964 102784 58976
rect 102836 58964 102842 59016
rect 201310 58964 201316 59016
rect 201368 59004 201374 59016
rect 300854 59004 300860 59016
rect 201368 58976 300860 59004
rect 201368 58964 201374 58976
rect 300854 58964 300860 58976
rect 300912 58964 300918 59016
rect 376570 58964 376576 59016
rect 376628 59004 376634 59016
rect 421742 59004 421748 59016
rect 376628 58976 421748 59004
rect 376628 58964 376634 58976
rect 421742 58964 421748 58976
rect 421800 58964 421806 59016
rect 58894 58896 58900 58948
rect 58952 58936 58958 58948
rect 107562 58936 107568 58948
rect 58952 58908 107568 58936
rect 58952 58896 58958 58908
rect 107562 58896 107568 58908
rect 107620 58896 107626 58948
rect 212350 58896 212356 58948
rect 212408 58936 212414 58948
rect 315850 58936 315856 58948
rect 212408 58908 315856 58936
rect 212408 58896 212414 58908
rect 315850 58896 315856 58908
rect 315908 58896 315914 58948
rect 362218 58896 362224 58948
rect 362276 58936 362282 58948
rect 423490 58936 423496 58948
rect 362276 58908 423496 58936
rect 362276 58896 362282 58908
rect 423490 58896 423496 58908
rect 423548 58896 423554 58948
rect 51626 58828 51632 58880
rect 51684 58868 51690 58880
rect 101766 58868 101772 58880
rect 51684 58840 101772 58868
rect 51684 58828 51690 58840
rect 101766 58828 101772 58840
rect 101824 58828 101830 58880
rect 202782 58828 202788 58880
rect 202840 58868 202846 58880
rect 308490 58868 308496 58880
rect 202840 58840 308496 58868
rect 202840 58828 202846 58840
rect 308490 58828 308496 58840
rect 308548 58828 308554 58880
rect 356698 58828 356704 58880
rect 356756 58868 356762 58880
rect 425974 58868 425980 58880
rect 356756 58840 425980 58868
rect 356756 58828 356762 58840
rect 425974 58828 425980 58840
rect 426032 58828 426038 58880
rect 53650 58760 53656 58812
rect 53708 58800 53714 58812
rect 138382 58800 138388 58812
rect 53708 58772 138388 58800
rect 53708 58760 53714 58772
rect 138382 58760 138388 58772
rect 138440 58760 138446 58812
rect 206186 58760 206192 58812
rect 206244 58800 206250 58812
rect 320910 58800 320916 58812
rect 206244 58772 320916 58800
rect 206244 58760 206250 58772
rect 320910 58760 320916 58772
rect 320968 58760 320974 58812
rect 366358 58760 366364 58812
rect 366416 58800 366422 58812
rect 453390 58800 453396 58812
rect 366416 58772 453396 58800
rect 366416 58760 366422 58772
rect 453390 58760 453396 58772
rect 453448 58760 453454 58812
rect 50982 58692 50988 58744
rect 51040 58732 51046 58744
rect 148502 58732 148508 58744
rect 51040 58704 148508 58732
rect 51040 58692 51046 58704
rect 148502 58692 148508 58704
rect 148560 58692 148566 58744
rect 198642 58692 198648 58744
rect 198700 58732 198706 58744
rect 325878 58732 325884 58744
rect 198700 58704 325884 58732
rect 198700 58692 198706 58704
rect 325878 58692 325884 58704
rect 325936 58692 325942 58744
rect 364978 58692 364984 58744
rect 365036 58732 365042 58744
rect 475838 58732 475844 58744
rect 365036 58704 475844 58732
rect 365036 58692 365042 58704
rect 475838 58692 475844 58704
rect 475896 58692 475902 58744
rect 53558 58624 53564 58676
rect 53616 58664 53622 58676
rect 150894 58664 150900 58676
rect 53616 58636 150900 58664
rect 53616 58624 53622 58636
rect 150894 58624 150900 58636
rect 150952 58624 150958 58676
rect 219250 58624 219256 58676
rect 219308 58664 219314 58676
rect 428182 58664 428188 58676
rect 219308 58636 428188 58664
rect 219308 58624 219314 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 57238 57876 57244 57928
rect 57296 57916 57302 57928
rect 57882 57916 57888 57928
rect 57296 57888 57888 57916
rect 57296 57876 57302 57888
rect 57882 57876 57888 57888
rect 57940 57916 57946 57928
rect 204898 57916 204904 57928
rect 57940 57888 204904 57916
rect 57940 57876 57946 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 210970 57876 210976 57928
rect 211028 57916 211034 57928
rect 323302 57916 323308 57928
rect 211028 57888 323308 57916
rect 211028 57876 211034 57888
rect 323302 57876 323308 57888
rect 323360 57876 323366 57928
rect 343450 57876 343456 57928
rect 343508 57916 343514 57928
rect 357618 57916 357624 57928
rect 343508 57888 357624 57916
rect 343508 57876 343514 57888
rect 357618 57876 357624 57888
rect 357676 57876 357682 57928
rect 358630 57876 358636 57928
rect 358688 57916 358694 57928
rect 478414 57916 478420 57928
rect 358688 57888 478420 57916
rect 358688 57876 358694 57888
rect 478414 57876 478420 57888
rect 478472 57876 478478 57928
rect 503254 57876 503260 57928
rect 503312 57916 503318 57928
rect 517606 57916 517612 57928
rect 503312 57888 517612 57916
rect 503312 57876 503318 57888
rect 517606 57876 517612 57888
rect 517664 57876 517670 57928
rect 52270 57808 52276 57860
rect 52328 57848 52334 57860
rect 145558 57848 145564 57860
rect 52328 57820 145564 57848
rect 52328 57808 52334 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183462 57808 183468 57860
rect 183520 57848 183526 57860
rect 197446 57848 197452 57860
rect 183520 57820 197452 57848
rect 183520 57808 183526 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 209682 57808 209688 57860
rect 209740 57848 209746 57860
rect 310974 57848 310980 57860
rect 209740 57820 310980 57848
rect 209740 57808 209746 57820
rect 310974 57808 310980 57820
rect 311032 57808 311038 57860
rect 343174 57808 343180 57860
rect 343232 57848 343238 57860
rect 357434 57848 357440 57860
rect 343232 57820 357440 57848
rect 343232 57808 343238 57820
rect 357434 57808 357440 57820
rect 357492 57808 357498 57860
rect 376662 57808 376668 57860
rect 376720 57848 376726 57860
rect 485958 57848 485964 57860
rect 376720 57820 485964 57848
rect 376720 57808 376726 57820
rect 485958 57808 485964 57820
rect 486016 57808 486022 57860
rect 503530 57808 503536 57860
rect 503588 57848 503594 57860
rect 517882 57848 517888 57860
rect 503588 57820 517888 57848
rect 503588 57808 503594 57820
rect 517882 57808 517888 57820
rect 517940 57808 517946 57860
rect 41230 57740 41236 57792
rect 41288 57780 41294 57792
rect 123478 57780 123484 57792
rect 41288 57752 123484 57780
rect 41288 57740 41294 57752
rect 123478 57740 123484 57752
rect 123536 57740 123542 57792
rect 183186 57740 183192 57792
rect 183244 57780 183250 57792
rect 197354 57780 197360 57792
rect 183244 57752 197360 57780
rect 183244 57740 183250 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 215202 57740 215208 57792
rect 215260 57780 215266 57792
rect 313366 57780 313372 57792
rect 215260 57752 313372 57780
rect 215260 57740 215266 57752
rect 313366 57740 313372 57752
rect 313424 57740 313430 57792
rect 363690 57740 363696 57792
rect 363748 57780 363754 57792
rect 465902 57780 465908 57792
rect 363748 57752 465908 57780
rect 363748 57740 363754 57752
rect 465902 57740 465908 57752
rect 465960 57740 465966 57792
rect 53742 57672 53748 57724
rect 53800 57712 53806 57724
rect 130838 57712 130844 57724
rect 53800 57684 130844 57712
rect 53800 57672 53806 57684
rect 130838 57672 130844 57684
rect 130896 57672 130902 57724
rect 218698 57672 218704 57724
rect 218756 57712 218762 57724
rect 318334 57712 318340 57724
rect 218756 57684 318340 57712
rect 218756 57672 218762 57684
rect 318334 57672 318340 57684
rect 318392 57672 318398 57724
rect 360838 57672 360844 57724
rect 360896 57712 360902 57724
rect 445846 57712 445852 57724
rect 360896 57684 445852 57712
rect 360896 57672 360902 57684
rect 445846 57672 445852 57684
rect 445904 57672 445910 57724
rect 53282 57604 53288 57656
rect 53340 57644 53346 57656
rect 113174 57644 113180 57656
rect 53340 57616 113180 57644
rect 53340 57604 53346 57616
rect 113174 57604 113180 57616
rect 113232 57604 113238 57656
rect 205542 57604 205548 57656
rect 205600 57644 205606 57656
rect 295886 57644 295892 57656
rect 205600 57616 295892 57644
rect 205600 57604 205606 57616
rect 295886 57604 295892 57616
rect 295944 57604 295950 57656
rect 363598 57604 363604 57656
rect 363656 57644 363662 57656
rect 448238 57644 448244 57656
rect 363656 57616 448244 57644
rect 363656 57604 363662 57616
rect 448238 57604 448244 57616
rect 448296 57604 448302 57656
rect 59078 57536 59084 57588
rect 59136 57576 59142 57588
rect 103790 57576 103796 57588
rect 59136 57548 103796 57576
rect 59136 57536 59142 57548
rect 103790 57536 103796 57548
rect 103848 57536 103854 57588
rect 213822 57536 213828 57588
rect 213880 57576 213886 57588
rect 303430 57576 303436 57588
rect 213880 57548 303436 57576
rect 213880 57536 213886 57548
rect 303430 57536 303436 57548
rect 303488 57536 303494 57588
rect 362310 57536 362316 57588
rect 362368 57576 362374 57588
rect 443454 57576 443460 57588
rect 362368 57548 443460 57576
rect 362368 57536 362374 57548
rect 443454 57536 443460 57548
rect 443512 57536 443518 57588
rect 55122 57468 55128 57520
rect 55180 57508 55186 57520
rect 98086 57508 98092 57520
rect 55180 57480 98092 57508
rect 55180 57468 55186 57480
rect 98086 57468 98092 57480
rect 98144 57468 98150 57520
rect 215570 57468 215576 57520
rect 215628 57508 215634 57520
rect 305822 57508 305828 57520
rect 215628 57480 305828 57508
rect 215628 57468 215634 57480
rect 305822 57468 305828 57480
rect 305880 57468 305886 57520
rect 367738 57468 367744 57520
rect 367796 57508 367802 57520
rect 435910 57508 435916 57520
rect 367796 57480 435916 57508
rect 367796 57468 367802 57480
rect 435910 57468 435916 57480
rect 435968 57468 435974 57520
rect 51534 57400 51540 57452
rect 51592 57440 51598 57452
rect 88334 57440 88340 57452
rect 51592 57412 88340 57440
rect 51592 57400 51598 57412
rect 88334 57400 88340 57412
rect 88392 57400 88398 57452
rect 211062 57400 211068 57452
rect 211120 57440 211126 57452
rect 293310 57440 293316 57452
rect 211120 57412 293316 57440
rect 211120 57400 211126 57412
rect 293310 57400 293316 57412
rect 293368 57400 293374 57452
rect 371878 57400 371884 57452
rect 371936 57440 371942 57452
rect 438486 57440 438492 57452
rect 371936 57412 438492 57440
rect 371936 57400 371942 57412
rect 438486 57400 438492 57412
rect 438544 57400 438550 57452
rect 59262 57332 59268 57384
rect 59320 57372 59326 57384
rect 93670 57372 93676 57384
rect 59320 57344 93676 57372
rect 59320 57332 59326 57344
rect 93670 57332 93676 57344
rect 93728 57332 93734 57384
rect 218422 57332 218428 57384
rect 218480 57372 218486 57384
rect 298094 57372 298100 57384
rect 218480 57344 298100 57372
rect 218480 57332 218486 57344
rect 298094 57332 298100 57344
rect 298152 57332 298158 57384
rect 370590 57332 370596 57384
rect 370648 57372 370654 57384
rect 433518 57372 433524 57384
rect 370648 57344 433524 57372
rect 370648 57332 370654 57344
rect 433518 57332 433524 57344
rect 433576 57332 433582 57384
rect 52362 57264 52368 57316
rect 52420 57304 52426 57316
rect 78214 57304 78220 57316
rect 52420 57276 78220 57304
rect 52420 57264 52426 57276
rect 78214 57264 78220 57276
rect 78272 57264 78278 57316
rect 211798 57264 211804 57316
rect 211856 57304 211862 57316
rect 283466 57304 283472 57316
rect 211856 57276 283472 57304
rect 211856 57264 211862 57276
rect 283466 57264 283472 57276
rect 283524 57264 283530 57316
rect 370498 57264 370504 57316
rect 370556 57304 370562 57316
rect 418430 57304 418436 57316
rect 370556 57276 418436 57304
rect 370556 57264 370562 57276
rect 418430 57264 418436 57276
rect 418488 57264 418494 57316
rect 54846 57196 54852 57248
rect 54904 57236 54910 57248
rect 76006 57236 76012 57248
rect 54904 57208 76012 57236
rect 54904 57196 54910 57208
rect 76006 57196 76012 57208
rect 76064 57196 76070 57248
rect 218606 57196 218612 57248
rect 218664 57236 218670 57248
rect 258350 57236 258356 57248
rect 218664 57208 258356 57236
rect 218664 57196 218670 57208
rect 258350 57196 258356 57208
rect 258408 57196 258414 57248
rect 379054 57196 379060 57248
rect 379112 57236 379118 57248
rect 415486 57236 415492 57248
rect 379112 57208 415492 57236
rect 379112 57196 379118 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 77846 56584 77852 56636
rect 77904 56624 77910 56636
rect 117866 56624 117872 56636
rect 77904 56596 117872 56624
rect 77904 56584 77910 56596
rect 117866 56584 117872 56596
rect 117924 56584 117930 56636
rect 41322 56516 41328 56568
rect 41380 56556 41386 56568
rect 115934 56556 115940 56568
rect 41380 56528 115940 56556
rect 41380 56516 41386 56528
rect 115934 56516 115940 56528
rect 115992 56516 115998 56568
rect 214558 56516 214564 56568
rect 214616 56556 214622 56568
rect 241606 56556 241612 56568
rect 214616 56528 241612 56556
rect 214616 56516 214622 56528
rect 241606 56516 241612 56528
rect 241664 56516 241670 56568
rect 374638 56516 374644 56568
rect 374696 56556 374702 56568
rect 398190 56556 398196 56568
rect 374696 56528 398196 56556
rect 374696 56516 374702 56528
rect 398190 56516 398196 56528
rect 398248 56516 398254 56568
rect 52178 56448 52184 56500
rect 52236 56488 52242 56500
rect 112070 56488 112076 56500
rect 52236 56460 112076 56488
rect 52236 56448 52242 56460
rect 112070 56448 112076 56460
rect 112128 56448 112134 56500
rect 219066 56448 219072 56500
rect 219124 56488 219130 56500
rect 235994 56488 236000 56500
rect 219124 56460 236000 56488
rect 219124 56448 219130 56460
rect 235994 56448 236000 56460
rect 236052 56448 236058 56500
rect 374546 56448 374552 56500
rect 374604 56488 374610 56500
rect 435726 56488 435732 56500
rect 374604 56460 435732 56488
rect 374604 56448 374610 56460
rect 435726 56448 435732 56460
rect 435784 56448 435790 56500
rect 56318 56380 56324 56432
rect 56376 56420 56382 56432
rect 114094 56420 114100 56432
rect 56376 56392 114100 56420
rect 56376 56380 56382 56392
rect 114094 56380 114100 56392
rect 114152 56380 114158 56432
rect 215018 56380 215024 56432
rect 215076 56420 215082 56432
rect 273254 56420 273260 56432
rect 215076 56392 273260 56420
rect 215076 56380 215082 56392
rect 273254 56380 273260 56392
rect 273312 56380 273318 56432
rect 373810 56380 373816 56432
rect 373868 56420 373874 56432
rect 433334 56420 433340 56432
rect 373868 56392 433340 56420
rect 373868 56380 373874 56392
rect 433334 56380 433340 56392
rect 433392 56380 433398 56432
rect 53374 56312 53380 56364
rect 53432 56352 53438 56364
rect 109494 56352 109500 56364
rect 53432 56324 109500 56352
rect 53432 56312 53438 56324
rect 109494 56312 109500 56324
rect 109552 56312 109558 56364
rect 214650 56312 214656 56364
rect 214708 56352 214714 56364
rect 271046 56352 271052 56364
rect 214708 56324 271052 56352
rect 214708 56312 214714 56324
rect 271046 56312 271052 56324
rect 271104 56312 271110 56364
rect 374822 56312 374828 56364
rect 374880 56352 374886 56364
rect 431126 56352 431132 56364
rect 374880 56324 431132 56352
rect 374880 56312 374886 56324
rect 431126 56312 431132 56324
rect 431184 56312 431190 56364
rect 59906 56244 59912 56296
rect 59964 56284 59970 56296
rect 108574 56284 108580 56296
rect 59964 56256 108580 56284
rect 59964 56244 59970 56256
rect 108574 56244 108580 56256
rect 108632 56244 108638 56296
rect 219894 56244 219900 56296
rect 219952 56284 219958 56296
rect 268470 56284 268476 56296
rect 219952 56256 268476 56284
rect 219952 56244 219958 56256
rect 268470 56244 268476 56256
rect 268528 56244 268534 56296
rect 379422 56244 379428 56296
rect 379480 56284 379486 56296
rect 427630 56284 427636 56296
rect 379480 56256 427636 56284
rect 379480 56244 379486 56256
rect 427630 56244 427636 56256
rect 427688 56244 427694 56296
rect 58710 56176 58716 56228
rect 58768 56216 58774 56228
rect 93302 56216 93308 56228
rect 58768 56188 93308 56216
rect 58768 56176 58774 56188
rect 93302 56176 93308 56188
rect 93360 56176 93366 56228
rect 219158 56176 219164 56228
rect 219216 56216 219222 56228
rect 266354 56216 266360 56228
rect 219216 56188 266360 56216
rect 219216 56176 219222 56188
rect 266354 56176 266360 56188
rect 266412 56176 266418 56228
rect 379698 56176 379704 56228
rect 379756 56216 379762 56228
rect 426434 56216 426440 56228
rect 379756 56188 426440 56216
rect 379756 56176 379762 56188
rect 426434 56176 426440 56188
rect 426492 56176 426498 56228
rect 56226 56108 56232 56160
rect 56284 56148 56290 56160
rect 88702 56148 88708 56160
rect 56284 56120 88708 56148
rect 56284 56108 56290 56120
rect 88702 56108 88708 56120
rect 88760 56108 88766 56160
rect 219342 56108 219348 56160
rect 219400 56148 219406 56160
rect 253382 56148 253388 56160
rect 219400 56120 253388 56148
rect 219400 56108 219406 56120
rect 253382 56108 253388 56120
rect 253440 56108 253446 56160
rect 379882 56108 379888 56160
rect 379940 56148 379946 56160
rect 414566 56148 414572 56160
rect 379940 56120 414572 56148
rect 379940 56108 379946 56120
rect 414566 56108 414572 56120
rect 414624 56108 414630 56160
rect 54938 56040 54944 56092
rect 54996 56080 55002 56092
rect 86494 56080 86500 56092
rect 54996 56052 86500 56080
rect 54996 56040 55002 56052
rect 86494 56040 86500 56052
rect 86552 56040 86558 56092
rect 218330 56040 218336 56092
rect 218388 56080 218394 56092
rect 251174 56080 251180 56092
rect 218388 56052 251180 56080
rect 218388 56040 218394 56052
rect 251174 56040 251180 56052
rect 251232 56040 251238 56092
rect 379330 56040 379336 56092
rect 379388 56080 379394 56092
rect 412634 56080 412640 56092
rect 379388 56052 412640 56080
rect 379388 56040 379394 56052
rect 412634 56040 412640 56052
rect 412692 56040 412698 56092
rect 51994 55972 52000 56024
rect 52052 56012 52058 56024
rect 80422 56012 80428 56024
rect 52052 55984 80428 56012
rect 52052 55972 52058 55984
rect 80422 55972 80428 55984
rect 80480 55972 80486 56024
rect 216122 55972 216128 56024
rect 216180 56012 216186 56024
rect 248598 56012 248604 56024
rect 216180 55984 248604 56012
rect 216180 55972 216186 55984
rect 248598 55972 248604 55984
rect 248656 55972 248662 56024
rect 378594 55972 378600 56024
rect 378652 56012 378658 56024
rect 411254 56012 411260 56024
rect 378652 55984 411260 56012
rect 378652 55972 378658 55984
rect 411254 55972 411260 55984
rect 411312 55972 411318 56024
rect 58802 55904 58808 55956
rect 58860 55944 58866 55956
rect 85390 55944 85396 55956
rect 58860 55916 85396 55944
rect 58860 55904 58866 55916
rect 85390 55904 85396 55916
rect 85448 55904 85454 55956
rect 216306 55904 216312 55956
rect 216364 55944 216370 55956
rect 245286 55944 245292 55956
rect 216364 55916 245292 55944
rect 216364 55904 216370 55916
rect 245286 55904 245292 55916
rect 245344 55904 245350 55956
rect 378778 55904 378784 55956
rect 378836 55944 378842 55956
rect 408678 55944 408684 55956
rect 378836 55916 408684 55944
rect 378836 55904 378842 55916
rect 408678 55904 408684 55916
rect 408736 55904 408742 55956
rect 213178 55836 213184 55888
rect 213236 55876 213242 55888
rect 239122 55876 239128 55888
rect 213236 55848 239128 55876
rect 213236 55836 213242 55848
rect 239122 55836 239128 55848
rect 239180 55836 239186 55888
rect 371970 55836 371976 55888
rect 372028 55876 372034 55888
rect 400398 55876 400404 55888
rect 372028 55848 400404 55876
rect 372028 55836 372034 55848
rect 400398 55836 400404 55848
rect 400456 55836 400462 55888
rect 219986 55768 219992 55820
rect 220044 55808 220050 55820
rect 408310 55808 408316 55820
rect 220044 55780 408316 55808
rect 220044 55768 220050 55780
rect 408310 55768 408316 55780
rect 408368 55768 408374 55820
rect 212994 55700 213000 55752
rect 213052 55740 213058 55752
rect 275094 55740 275100 55752
rect 213052 55712 275100 55740
rect 213052 55700 213058 55712
rect 275094 55700 275100 55712
rect 275152 55700 275158 55752
rect 53006 55156 53012 55208
rect 53064 55196 53070 55208
rect 114554 55196 114560 55208
rect 53064 55168 114560 55196
rect 53064 55156 53070 55168
rect 114554 55156 114560 55168
rect 114612 55156 114618 55208
rect 216490 55156 216496 55208
rect 216548 55196 216554 55208
rect 277394 55196 277400 55208
rect 216548 55168 277400 55196
rect 216548 55156 216554 55168
rect 277394 55156 277400 55168
rect 277452 55156 277458 55208
rect 375834 55156 375840 55208
rect 375892 55196 375898 55208
rect 436094 55196 436100 55208
rect 375892 55168 436100 55196
rect 375892 55156 375898 55168
rect 436094 55156 436100 55168
rect 436152 55156 436158 55208
rect 56410 55088 56416 55140
rect 56468 55128 56474 55140
rect 116118 55128 116124 55140
rect 56468 55100 116124 55128
rect 56468 55088 56474 55100
rect 116118 55088 116124 55100
rect 116176 55088 116182 55140
rect 213730 55088 213736 55140
rect 213788 55128 213794 55140
rect 273346 55128 273352 55140
rect 213788 55100 273352 55128
rect 213788 55088 213794 55100
rect 273346 55088 273352 55100
rect 273404 55088 273410 55140
rect 376018 55088 376024 55140
rect 376076 55128 376082 55140
rect 398834 55128 398840 55140
rect 376076 55100 398840 55128
rect 376076 55088 376082 55100
rect 398834 55088 398840 55100
rect 398892 55088 398898 55140
rect 53466 55020 53472 55072
rect 53524 55060 53530 55072
rect 110414 55060 110420 55072
rect 53524 55032 110420 55060
rect 53524 55020 53530 55032
rect 110414 55020 110420 55032
rect 110472 55020 110478 55072
rect 215938 55020 215944 55072
rect 215996 55060 216002 55072
rect 271874 55060 271880 55072
rect 215996 55032 271880 55060
rect 215996 55020 216002 55032
rect 271874 55020 271880 55032
rect 271932 55020 271938 55072
rect 375098 55020 375104 55072
rect 375156 55060 375162 55072
rect 431954 55060 431960 55072
rect 375156 55032 431960 55060
rect 375156 55020 375162 55032
rect 431954 55020 431960 55032
rect 432012 55020 432018 55072
rect 42702 54952 42708 55004
rect 42760 54992 42766 55004
rect 89714 54992 89720 55004
rect 42760 54964 89720 54992
rect 42760 54952 42766 54964
rect 89714 54952 89720 54964
rect 89772 54952 89778 55004
rect 219526 54952 219532 55004
rect 219584 54992 219590 55004
rect 266446 54992 266452 55004
rect 219584 54964 266452 54992
rect 219584 54952 219590 54964
rect 266446 54952 266452 54964
rect 266504 54952 266510 55004
rect 375006 54952 375012 55004
rect 375064 54992 375070 55004
rect 429194 54992 429200 55004
rect 375064 54964 429200 54992
rect 375064 54952 375070 54964
rect 429194 54952 429200 54964
rect 429252 54952 429258 55004
rect 59998 54884 60004 54936
rect 60056 54924 60062 54936
rect 106274 54924 106280 54936
rect 60056 54896 106280 54924
rect 60056 54884 60062 54896
rect 106274 54884 106280 54896
rect 106332 54884 106338 54936
rect 219618 54884 219624 54936
rect 219676 54924 219682 54936
rect 264974 54924 264980 54936
rect 219676 54896 264980 54924
rect 219676 54884 219682 54896
rect 264974 54884 264980 54896
rect 265032 54884 265038 54936
rect 379974 54884 379980 54936
rect 380032 54924 380038 54936
rect 427814 54924 427820 54936
rect 380032 54896 427820 54924
rect 380032 54884 380038 54896
rect 427814 54884 427820 54896
rect 427872 54884 427878 54936
rect 57054 54816 57060 54868
rect 57112 54856 57118 54868
rect 91094 54856 91100 54868
rect 57112 54828 91100 54856
rect 57112 54816 57118 54828
rect 91094 54816 91100 54828
rect 91152 54816 91158 54868
rect 219710 54816 219716 54868
rect 219768 54856 219774 54868
rect 253934 54856 253940 54868
rect 219768 54828 253940 54856
rect 219768 54816 219774 54828
rect 253934 54816 253940 54828
rect 253992 54816 253998 54868
rect 378042 54816 378048 54868
rect 378100 54856 378106 54868
rect 411346 54856 411352 54868
rect 378100 54828 411352 54856
rect 378100 54816 378106 54828
rect 411346 54816 411352 54828
rect 411404 54816 411410 54868
rect 52914 54748 52920 54800
rect 52972 54788 52978 54800
rect 86954 54788 86960 54800
rect 52972 54760 86960 54788
rect 52972 54748 52978 54760
rect 86954 54748 86960 54760
rect 87012 54748 87018 54800
rect 217042 54748 217048 54800
rect 217100 54788 217106 54800
rect 251358 54788 251364 54800
rect 217100 54760 251364 54788
rect 217100 54748 217106 54760
rect 251358 54748 251364 54760
rect 251416 54748 251422 54800
rect 377858 54748 377864 54800
rect 377916 54788 377922 54800
rect 409874 54788 409880 54800
rect 377916 54760 409880 54788
rect 377916 54748 377922 54760
rect 409874 54748 409880 54760
rect 409932 54748 409938 54800
rect 58618 54680 58624 54732
rect 58676 54720 58682 54732
rect 91462 54720 91468 54732
rect 58676 54692 91468 54720
rect 58676 54680 58682 54692
rect 91462 54680 91468 54692
rect 91520 54680 91526 54732
rect 217870 54680 217876 54732
rect 217928 54720 217934 54732
rect 249794 54720 249800 54732
rect 217928 54692 249800 54720
rect 217928 54680 217934 54692
rect 249794 54680 249800 54692
rect 249852 54680 249858 54732
rect 376478 54680 376484 54732
rect 376536 54720 376542 54732
rect 407206 54720 407212 54732
rect 376536 54692 407212 54720
rect 376536 54680 376542 54692
rect 407206 54680 407212 54692
rect 407264 54680 407270 54732
rect 53190 54612 53196 54664
rect 53248 54652 53254 54664
rect 81434 54652 81440 54664
rect 53248 54624 81440 54652
rect 53248 54612 53254 54624
rect 81434 54612 81440 54624
rect 81492 54612 81498 54664
rect 216398 54612 216404 54664
rect 216456 54652 216462 54664
rect 247034 54652 247040 54664
rect 216456 54624 247040 54652
rect 216456 54612 216462 54624
rect 247034 54612 247040 54624
rect 247092 54612 247098 54664
rect 375282 54612 375288 54664
rect 375340 54652 375346 54664
rect 405826 54652 405832 54664
rect 375340 54624 405832 54652
rect 375340 54612 375346 54624
rect 405826 54612 405832 54624
rect 405884 54612 405890 54664
rect 51718 54544 51724 54596
rect 51776 54584 51782 54596
rect 78674 54584 78680 54596
rect 51776 54556 78680 54584
rect 51776 54544 51782 54556
rect 78674 54544 78680 54556
rect 78732 54544 78738 54596
rect 215110 54544 215116 54596
rect 215168 54584 215174 54596
rect 244366 54584 244372 54596
rect 215168 54556 244372 54584
rect 215168 54544 215174 54556
rect 244366 54544 244372 54556
rect 244424 54544 244430 54596
rect 375926 54544 375932 54596
rect 375984 54584 375990 54596
rect 404354 54584 404360 54596
rect 375984 54556 404360 54584
rect 375984 54544 375990 54556
rect 404354 54544 404360 54556
rect 404412 54544 404418 54596
rect 218790 54476 218796 54528
rect 218848 54516 218854 54528
rect 245654 54516 245660 54528
rect 218848 54488 245660 54516
rect 218848 54476 218854 54488
rect 245654 54476 245660 54488
rect 245712 54476 245718 54528
rect 373258 54476 373264 54528
rect 373316 54516 373322 54528
rect 401594 54516 401600 54528
rect 373316 54488 401600 54516
rect 373316 54476 373322 54488
rect 401594 54476 401600 54488
rect 401652 54476 401658 54528
rect 216030 54408 216036 54460
rect 216088 54448 216094 54460
rect 242894 54448 242900 54460
rect 216088 54420 242900 54448
rect 216088 54408 216094 54420
rect 242894 54408 242900 54420
rect 242952 54408 242958 54460
rect 373718 54408 373724 54460
rect 373776 54448 373782 54460
rect 433426 54448 433432 54460
rect 373776 54420 433432 54448
rect 373776 54408 373782 54420
rect 433426 54408 433432 54420
rect 433484 54408 433490 54460
rect 213270 54340 213276 54392
rect 213328 54380 213334 54392
rect 237374 54380 237380 54392
rect 213328 54352 237380 54380
rect 213328 54340 213334 54352
rect 237374 54340 237380 54352
rect 237432 54340 237438 54392
rect 213638 54272 213644 54324
rect 213696 54312 213702 54324
rect 240134 54312 240140 54324
rect 213696 54284 240140 54312
rect 213696 54272 213702 54284
rect 240134 54272 240140 54284
rect 240192 54272 240198 54324
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 125870 2796 125876 2848
rect 125928 2836 125934 2848
rect 367094 2836 367100 2848
rect 125928 2808 367100 2836
rect 125928 2796 125934 2808
rect 367094 2796 367100 2808
rect 367152 2796 367158 2848
<< via1 >>
rect 235172 700272 235224 700324
rect 304264 700272 304316 700324
rect 137744 683136 137796 683188
rect 580172 683136 580224 683188
rect 59084 649272 59136 649324
rect 542360 649272 542412 649324
rect 104900 647844 104952 647896
rect 429384 647844 429436 647896
rect 299480 646484 299532 646536
rect 401140 646484 401192 646536
rect 169760 645124 169812 645176
rect 430580 645124 430632 645176
rect 364340 643696 364392 643748
rect 423680 643696 423732 643748
rect 317052 643152 317104 643204
rect 430764 643152 430816 643204
rect 284944 643084 284996 643136
rect 430672 643084 430724 643136
rect 318800 642336 318852 642388
rect 494060 642336 494112 642388
rect 289820 641724 289872 641776
rect 435364 641724 435416 641776
rect 287704 641180 287756 641232
rect 378600 641180 378652 641232
rect 311256 641112 311308 641164
rect 332876 641112 332928 641164
rect 312636 641044 312688 641096
rect 337384 641044 337436 641096
rect 319628 640976 319680 641028
rect 355416 640976 355468 641028
rect 315304 640908 315356 640960
rect 359924 640908 359976 640960
rect 316684 640840 316736 640892
rect 364432 640840 364484 640892
rect 302884 640772 302936 640824
rect 350908 640772 350960 640824
rect 319812 640704 319864 640756
rect 373448 640704 373500 640756
rect 314016 640636 314068 640688
rect 368940 640636 368992 640688
rect 316868 640568 316920 640620
rect 387616 640568 387668 640620
rect 309784 640500 309836 640552
rect 383108 640500 383160 640552
rect 316960 640432 317012 640484
rect 396632 640432 396684 640484
rect 318156 640364 318208 640416
rect 428188 640364 428240 640416
rect 319536 640296 319588 640348
rect 323860 640296 323912 640348
rect 414664 640296 414716 640348
rect 457444 640296 457496 640348
rect 280712 639616 280764 639668
rect 341892 639616 341944 639668
rect 298100 639548 298152 639600
rect 428464 639548 428516 639600
rect 296720 639480 296772 639532
rect 432604 639480 432656 639532
rect 291200 639412 291252 639464
rect 429844 639412 429896 639464
rect 318340 639344 318392 639396
rect 457536 639344 457588 639396
rect 319444 639276 319496 639328
rect 470600 639276 470652 639328
rect 293960 639208 294012 639260
rect 512000 639208 512052 639260
rect 287060 639140 287112 639192
rect 510620 639140 510672 639192
rect 219164 639072 219216 639124
rect 580264 639072 580316 639124
rect 18604 639004 18656 639056
rect 409880 639004 409932 639056
rect 218704 638936 218756 638988
rect 414572 638936 414624 638988
rect 311164 637644 311216 637696
rect 317972 637644 318024 637696
rect 288440 637576 288492 637628
rect 512092 637576 512144 637628
rect 3424 636828 3476 636880
rect 316776 636828 316828 636880
rect 114192 634040 114244 634092
rect 121644 634040 121696 634092
rect 131120 634040 131172 634092
rect 151268 634040 151320 634092
rect 210424 634040 210476 634092
rect 219716 634040 219768 634092
rect 115664 633972 115716 634024
rect 124588 633972 124640 634024
rect 135260 633972 135312 634024
rect 183560 633972 183612 634024
rect 213920 633972 213972 634024
rect 225420 633972 225472 634024
rect 112536 633904 112588 633956
rect 123024 633904 123076 633956
rect 135168 633904 135220 633956
rect 160284 633904 160336 633956
rect 212540 633904 212592 633956
rect 271880 633904 271932 633956
rect 69296 633836 69348 633888
rect 127072 633836 127124 633888
rect 136548 633836 136600 633888
rect 162860 633836 162912 633888
rect 217876 633836 217928 633888
rect 242900 633836 242952 633888
rect 106648 633768 106700 633820
rect 121460 633768 121512 633820
rect 139124 633768 139176 633820
rect 166172 633768 166224 633820
rect 218888 633768 218940 633820
rect 251916 633768 251968 633820
rect 56508 633632 56560 633684
rect 77300 633632 77352 633684
rect 104072 633632 104124 633684
rect 114192 633632 114244 633684
rect 54852 633564 54904 633616
rect 88708 633564 88760 633616
rect 100668 633564 100720 633616
rect 122840 633700 122892 633752
rect 139216 633700 139268 633752
rect 174452 633700 174504 633752
rect 218796 633700 218848 633752
rect 263600 633700 263652 633752
rect 118240 633632 118292 633684
rect 124312 633632 124364 633684
rect 134892 633632 134944 633684
rect 180340 633632 180392 633684
rect 190000 633632 190052 633684
rect 204444 633632 204496 633684
rect 209780 633632 209832 633684
rect 260196 633632 260248 633684
rect 124220 633564 124272 633616
rect 171876 633564 171928 633616
rect 214012 633564 214064 633616
rect 269212 633564 269264 633616
rect 55128 633496 55180 633548
rect 91836 633496 91888 633548
rect 95056 633496 95108 633548
rect 120908 633496 120960 633548
rect 137652 633496 137704 633548
rect 109960 633428 110012 633480
rect 121000 633428 121052 633480
rect 133880 633428 133932 633480
rect 139676 633428 139728 633480
rect 140136 633496 140188 633548
rect 157524 633496 157576 633548
rect 192576 633496 192628 633548
rect 201684 633496 201736 633548
rect 219348 633496 219400 633548
rect 275100 633496 275152 633548
rect 186504 633428 186556 633480
rect 195704 633428 195756 633480
rect 200856 633428 200908 633480
rect 217324 633428 217376 633480
rect 231308 633428 231360 633480
rect 270408 633428 270460 633480
rect 277676 633428 277728 633480
rect 204260 632680 204312 632732
rect 270408 632680 270460 632732
rect 215300 632272 215352 632324
rect 234620 632272 234672 632324
rect 208400 632204 208452 632256
rect 240324 632204 240376 632256
rect 206284 632136 206336 632188
rect 254492 632136 254544 632188
rect 3424 632068 3476 632120
rect 313924 632068 313976 632120
rect 59360 631320 59412 631372
rect 97724 631320 97776 631372
rect 134984 631048 135036 631100
rect 142988 631048 143040 631100
rect 217968 631048 218020 631100
rect 228732 631048 228784 631100
rect 124864 630980 124916 631032
rect 178132 630980 178184 631032
rect 204352 630980 204404 631032
rect 222844 630980 222896 631032
rect 57796 630912 57848 630964
rect 80244 630912 80296 630964
rect 136456 630912 136508 630964
rect 149152 630912 149204 630964
rect 204904 630912 204956 630964
rect 237288 630912 237340 630964
rect 59268 630844 59320 630896
rect 65524 630844 65576 630896
rect 135076 630844 135128 630896
rect 154580 630844 154632 630896
rect 206376 630844 206428 630896
rect 248696 630844 248748 630896
rect 56416 630776 56468 630828
rect 71228 630776 71280 630828
rect 136640 630776 136692 630828
rect 168748 630776 168800 630828
rect 213184 630776 213236 630828
rect 257620 630776 257672 630828
rect 54944 630708 54996 630760
rect 74632 630708 74684 630760
rect 86776 630708 86828 630760
rect 124496 630708 124548 630760
rect 137836 630708 137888 630760
rect 145564 630708 145616 630760
rect 211804 630708 211856 630760
rect 266268 630708 266320 630760
rect 55036 630640 55088 630692
rect 62948 630640 63000 630692
rect 83464 630640 83516 630692
rect 124404 630640 124456 630692
rect 137928 630640 137980 630692
rect 218704 630640 218756 630692
rect 219440 630640 219492 630692
rect 246028 630640 246080 630692
rect 280712 630504 280764 630556
rect 139860 630368 139912 630420
rect 140136 630368 140188 630420
rect 198280 630368 198332 630420
rect 201592 630368 201644 630420
rect 280712 630300 280764 630352
rect 435364 630028 435416 630080
rect 483204 630028 483256 630080
rect 432604 629960 432656 630012
rect 494796 629960 494848 630012
rect 428464 629892 428516 629944
rect 501236 629892 501288 629944
rect 294604 627920 294656 627972
rect 317696 627920 317748 627972
rect 465448 627920 465500 627972
rect 580264 627920 580316 627972
rect 429844 627852 429896 627904
rect 456800 627852 456852 627904
rect 208492 625132 208544 625184
rect 216680 625132 216732 625184
rect 312544 623772 312596 623824
rect 317420 623772 317472 623824
rect 206468 619624 206520 619676
rect 216680 619624 216732 619676
rect 307024 618264 307076 618316
rect 317604 618264 317656 618316
rect 132500 615884 132552 615936
rect 136732 615884 136784 615936
rect 204996 615476 205048 615528
rect 216680 615476 216732 615528
rect 287796 614116 287848 614168
rect 317972 614116 318024 614168
rect 295984 608608 296036 608660
rect 317972 608608 318024 608660
rect 286324 604460 286376 604512
rect 317972 604460 318024 604512
rect 126244 597524 126296 597576
rect 136732 597524 136784 597576
rect 213276 597524 213328 597576
rect 216680 597524 216732 597576
rect 302240 596776 302292 596828
rect 318340 596776 318392 596828
rect 203248 596640 203300 596692
rect 204536 596640 204588 596692
rect 124128 596164 124180 596216
rect 134524 596164 134576 596216
rect 283656 596164 283708 596216
rect 302240 596164 302292 596216
rect 211160 594804 211212 594856
rect 216680 594804 216732 594856
rect 285036 594804 285088 594856
rect 317972 594804 318024 594856
rect 210516 590656 210568 590708
rect 216680 590656 216732 590708
rect 286416 589296 286468 589348
rect 317972 589296 318024 589348
rect 125600 585148 125652 585200
rect 136732 585148 136784 585200
rect 289084 585148 289136 585200
rect 317972 585148 318024 585200
rect 129004 582360 129056 582412
rect 136732 582360 136784 582412
rect 206560 582360 206612 582412
rect 216680 582360 216732 582412
rect 209044 579640 209096 579692
rect 216680 579640 216732 579692
rect 287888 579640 287940 579692
rect 317972 579640 318024 579692
rect 513012 579640 513064 579692
rect 560944 579640 560996 579692
rect 138572 572296 138624 572348
rect 139124 572296 139176 572348
rect 207020 570596 207072 570648
rect 217416 570596 217468 570648
rect 137376 569848 137428 569900
rect 139768 569848 139820 569900
rect 200948 569848 201000 569900
rect 202972 569848 203024 569900
rect 57888 569168 57940 569220
rect 138020 569168 138072 569220
rect 57244 569100 57296 569152
rect 59912 569100 59964 569152
rect 217692 568556 217744 568608
rect 219900 568556 219952 568608
rect 3424 568488 3476 568540
rect 286416 568488 286468 568540
rect 58716 568420 58768 568472
rect 60740 568420 60792 568472
rect 134524 568420 134576 568472
rect 204536 568420 204588 568472
rect 302240 568420 302292 568472
rect 57152 568352 57204 568404
rect 61384 568352 61436 568404
rect 106280 568216 106332 568268
rect 124588 568216 124640 568268
rect 164332 568216 164384 568268
rect 200856 568216 200908 568268
rect 99564 568148 99616 568200
rect 122196 568148 122248 568200
rect 137652 568148 137704 568200
rect 145288 568148 145340 568200
rect 182364 568148 182416 568200
rect 218888 568148 218940 568200
rect 96712 568080 96764 568132
rect 123024 568080 123076 568132
rect 139032 568080 139084 568132
rect 150624 568080 150676 568132
rect 154580 568080 154632 568132
rect 201684 568080 201736 568132
rect 54852 568012 54904 568064
rect 78772 568012 78824 568064
rect 93860 568012 93912 568064
rect 122840 568012 122892 568064
rect 134892 568012 134944 568064
rect 151820 568012 151872 568064
rect 156052 568012 156104 568064
rect 204444 568012 204496 568064
rect 219348 568012 219400 568064
rect 223580 568012 223632 568064
rect 242164 568012 242216 568064
rect 281080 568012 281132 568064
rect 58808 567944 58860 567996
rect 91100 567944 91152 567996
rect 98092 567944 98144 567996
rect 121000 567944 121052 567996
rect 122196 567944 122248 567996
rect 201776 567944 201828 567996
rect 217876 567944 217928 567996
rect 222200 567944 222252 567996
rect 260840 567944 260892 567996
rect 317052 567944 317104 567996
rect 58532 567876 58584 567928
rect 67640 567876 67692 567928
rect 78680 567876 78732 567928
rect 122288 567876 122340 567928
rect 139216 567876 139268 567928
rect 158720 567876 158772 567928
rect 194600 567876 194652 567928
rect 283564 567876 283616 567928
rect 64880 567808 64932 567860
rect 123392 567808 123444 567860
rect 138572 567808 138624 567860
rect 161664 567808 161716 567860
rect 179420 567808 179472 567860
rect 282184 567808 282236 567860
rect 139124 567604 139176 567656
rect 142160 567604 142212 567656
rect 87052 566788 87104 566840
rect 121460 566788 121512 566840
rect 157984 566788 158036 566840
rect 203156 566788 203208 566840
rect 111892 566720 111944 566772
rect 121552 566720 121604 566772
rect 125692 566720 125744 566772
rect 200764 566720 200816 566772
rect 58992 566652 59044 566704
rect 77300 566652 77352 566704
rect 84200 566652 84252 566704
rect 122104 566652 122156 566704
rect 200304 566652 200356 566704
rect 283472 566652 283524 566704
rect 57520 566584 57572 566636
rect 82912 566584 82964 566636
rect 86960 566584 87012 566636
rect 124312 566584 124364 566636
rect 187792 566584 187844 566636
rect 281724 566584 281776 566636
rect 69020 566516 69072 566568
rect 123484 566516 123536 566568
rect 180892 566516 180944 566568
rect 281908 566516 281960 566568
rect 67732 566448 67784 566500
rect 121920 566448 121972 566500
rect 137192 566448 137244 566500
rect 160100 566448 160152 566500
rect 180800 566448 180852 566500
rect 281816 566448 281868 566500
rect 137560 566244 137612 566296
rect 140780 566244 140832 566296
rect 139860 566040 139912 566092
rect 140872 566040 140924 566092
rect 59084 565972 59136 566024
rect 62120 565972 62172 566024
rect 267740 565836 267792 565888
rect 317972 565836 318024 565888
rect 151360 565632 151412 565684
rect 160744 565632 160796 565684
rect 148784 565564 148836 565616
rect 159364 565564 159416 565616
rect 143540 565496 143592 565548
rect 156420 565496 156472 565548
rect 159916 565496 159968 565548
rect 164884 565496 164936 565548
rect 82728 565428 82780 565480
rect 89812 565428 89864 565480
rect 147772 565428 147824 565480
rect 162308 565428 162360 565480
rect 231860 565428 231912 565480
rect 259644 565428 259696 565480
rect 74540 565360 74592 565412
rect 96988 565360 97040 565412
rect 100208 565360 100260 565412
rect 115204 565360 115256 565412
rect 154672 565360 154724 565412
rect 171324 565360 171376 565412
rect 182824 565360 182876 565412
rect 77024 565292 77076 565344
rect 84844 565292 84896 565344
rect 86040 565292 86092 565344
rect 108304 565292 108356 565344
rect 129740 565292 129792 565344
rect 153844 565292 153896 565344
rect 158812 565292 158864 565344
rect 182916 565292 182968 565344
rect 222384 565360 222436 565412
rect 253940 565360 253992 565412
rect 203340 565292 203392 565344
rect 212632 565292 212684 565344
rect 251272 565292 251324 565344
rect 252560 565292 252612 565344
rect 316960 565292 317012 565344
rect 68744 565224 68796 565276
rect 105544 565224 105596 565276
rect 118700 565224 118752 565276
rect 145104 565224 145156 565276
rect 147680 565224 147732 565276
rect 185492 565224 185544 565276
rect 190644 565224 190696 565276
rect 257068 565224 257120 565276
rect 269120 565224 269172 565276
rect 289084 565224 289136 565276
rect 71320 565156 71372 565208
rect 108396 565156 108448 565208
rect 110420 565156 110472 565208
rect 120724 565156 120776 565208
rect 133972 565156 134024 565208
rect 197452 565156 197504 565208
rect 227720 565156 227772 565208
rect 245660 565156 245712 565208
rect 247040 565156 247092 565208
rect 319812 565156 319864 565208
rect 62856 565088 62908 565140
rect 72424 565088 72476 565140
rect 75920 565088 75972 565140
rect 117412 565088 117464 565140
rect 132592 565088 132644 565140
rect 177028 565088 177080 565140
rect 191840 565088 191892 565140
rect 276940 565088 276992 565140
rect 60280 565020 60332 565072
rect 62580 565020 62632 565072
rect 94504 564884 94556 564936
rect 102784 564884 102836 564936
rect 187700 564884 187752 564936
rect 191196 564884 191248 564936
rect 113180 564476 113232 564528
rect 121184 564476 121236 564528
rect 71780 564408 71832 564460
rect 73804 564408 73856 564460
rect 100760 564408 100812 564460
rect 102876 564408 102928 564460
rect 106924 564408 106976 564460
rect 108580 564408 108632 564460
rect 116584 564408 116636 564460
rect 120172 564408 120224 564460
rect 173164 564408 173216 564460
rect 173992 564408 174044 564460
rect 198004 564408 198056 564460
rect 200212 564408 200264 564460
rect 225144 564408 225196 564460
rect 227996 564408 228048 564460
rect 260104 564408 260156 564460
rect 262772 564408 262824 564460
rect 264244 564408 264296 564460
rect 265348 564408 265400 564460
rect 267004 564408 267056 564460
rect 268660 564408 268712 564460
rect 269764 564408 269816 564460
rect 271236 564408 271288 564460
rect 278044 564408 278096 564460
rect 280252 564408 280304 564460
rect 274824 563932 274876 563984
rect 312636 563932 312688 563984
rect 57428 563864 57480 563916
rect 87604 563864 87656 563916
rect 128360 563864 128412 563916
rect 201960 563864 202012 563916
rect 226432 563864 226484 563916
rect 280804 563864 280856 563916
rect 85672 563796 85724 563848
rect 121828 563796 121880 563848
rect 122840 563796 122892 563848
rect 201040 563796 201092 563848
rect 219256 563796 219308 563848
rect 223672 563796 223724 563848
rect 255320 563796 255372 563848
rect 318248 563796 318300 563848
rect 59452 563728 59504 563780
rect 76012 563728 76064 563780
rect 80060 563728 80112 563780
rect 123300 563728 123352 563780
rect 195980 563728 196032 563780
rect 283288 563728 283340 563780
rect 63500 563660 63552 563712
rect 123668 563660 123720 563712
rect 138848 563660 138900 563712
rect 160192 563660 160244 563712
rect 179604 563660 179656 563712
rect 281540 563660 281592 563712
rect 266360 562572 266412 562624
rect 302884 562572 302936 562624
rect 120172 562504 120224 562556
rect 187700 562504 187752 562556
rect 198740 562504 198792 562556
rect 206468 562504 206520 562556
rect 215392 562504 215444 562556
rect 282092 562504 282144 562556
rect 80152 562436 80204 562488
rect 121092 562436 121144 562488
rect 126980 562436 127032 562488
rect 201500 562436 201552 562488
rect 234620 562436 234672 562488
rect 319720 562436 319772 562488
rect 57060 562368 57112 562420
rect 110512 562368 110564 562420
rect 138756 562368 138808 562420
rect 63592 562300 63644 562352
rect 122932 562300 122984 562352
rect 139400 562300 139452 562352
rect 139952 562300 140004 562352
rect 184940 562368 184992 562420
rect 274640 562368 274692 562420
rect 173900 562300 173952 562352
rect 186320 562300 186372 562352
rect 282000 562300 282052 562352
rect 281540 562232 281592 562284
rect 285036 562300 285088 562352
rect 190552 561144 190604 561196
rect 204996 561144 205048 561196
rect 88616 561076 88668 561128
rect 103520 561076 103572 561128
rect 193220 561076 193272 561128
rect 218796 561076 218848 561128
rect 59176 561008 59228 561060
rect 92572 561008 92624 561060
rect 142252 561008 142304 561060
rect 203248 561008 203300 561060
rect 217600 561008 217652 561060
rect 231952 561008 232004 561060
rect 263600 561008 263652 561060
rect 311256 561008 311308 561060
rect 70400 560940 70452 560992
rect 120816 560940 120868 560992
rect 138940 560940 138992 560992
rect 165712 560940 165764 560992
rect 201500 560940 201552 560992
rect 283012 560940 283064 560992
rect 21364 560260 21416 560312
rect 317972 560260 318024 560312
rect 266452 559784 266504 559836
rect 287704 559784 287756 559836
rect 88432 559716 88484 559768
rect 104900 559716 104952 559768
rect 176660 559716 176712 559768
rect 213276 559716 213328 559768
rect 273260 559716 273312 559768
rect 318156 559716 318208 559768
rect 129832 559648 129884 559700
rect 202880 559648 202932 559700
rect 240140 559648 240192 559700
rect 314016 559648 314068 559700
rect 62580 559580 62632 559632
rect 104992 559580 105044 559632
rect 122932 559580 122984 559632
rect 201868 559580 201920 559632
rect 233332 559580 233384 559632
rect 319628 559580 319680 559632
rect 65064 559512 65116 559564
rect 123116 559512 123168 559564
rect 138664 559512 138716 559564
rect 168472 559512 168524 559564
rect 196072 559512 196124 559564
rect 283380 559512 283432 559564
rect 219624 558424 219676 558476
rect 247132 558424 247184 558476
rect 279516 558424 279568 558476
rect 294604 558424 294656 558476
rect 176752 558356 176804 558408
rect 225052 558356 225104 558408
rect 256700 558356 256752 558408
rect 309784 558356 309836 558408
rect 57612 558288 57664 558340
rect 107752 558288 107804 558340
rect 134524 558288 134576 558340
rect 187884 558288 187936 558340
rect 197360 558288 197412 558340
rect 209044 558288 209096 558340
rect 227812 558288 227864 558340
rect 282920 558288 282972 558340
rect 70492 558220 70544 558272
rect 121736 558220 121788 558272
rect 124312 558220 124364 558272
rect 201224 558220 201276 558272
rect 245660 558220 245712 558272
rect 307024 558220 307076 558272
rect 66352 558152 66404 558204
rect 123576 558152 123628 558204
rect 137928 558152 137980 558204
rect 149152 558152 149204 558204
rect 186412 558152 186464 558204
rect 283104 558152 283156 558204
rect 40040 557472 40092 557524
rect 317420 557472 317472 557524
rect 192116 556996 192168 557048
rect 210424 556996 210476 557048
rect 188528 556928 188580 556980
rect 233240 556928 233292 556980
rect 260196 556928 260248 556980
rect 287888 556928 287940 556980
rect 78864 556860 78916 556912
rect 115388 556860 115440 556912
rect 152648 556860 152700 556912
rect 202052 556860 202104 556912
rect 229284 556860 229336 556912
rect 281264 556860 281316 556912
rect 58900 556792 58952 556844
rect 102508 556792 102560 556844
rect 140504 556792 140556 556844
rect 198004 556792 198056 556844
rect 245108 556792 245160 556844
rect 315304 556792 315356 556844
rect 124220 556452 124272 556504
rect 125416 556452 125468 556504
rect 126980 556316 127032 556368
rect 128268 556316 128320 556368
rect 217784 556180 217836 556232
rect 218612 556180 218664 556232
rect 219624 556044 219676 556096
rect 220728 556044 220780 556096
rect 222200 555772 222252 555824
rect 222844 555772 222896 555824
rect 193496 555636 193548 555688
rect 215944 555636 215996 555688
rect 217876 555636 217928 555688
rect 260104 555636 260156 555688
rect 94596 555568 94648 555620
rect 122012 555568 122064 555620
rect 142344 555568 142396 555620
rect 167736 555568 167788 555620
rect 178500 555568 178552 555620
rect 206560 555568 206612 555620
rect 250076 555568 250128 555620
rect 295984 555568 296036 555620
rect 58440 555500 58492 555552
rect 103244 555500 103296 555552
rect 144092 555500 144144 555552
rect 202236 555500 202288 555552
rect 208492 555500 208544 555552
rect 236000 555500 236052 555552
rect 236092 555500 236144 555552
rect 283196 555500 283248 555552
rect 63132 555432 63184 555484
rect 110604 555432 110656 555484
rect 121828 555432 121880 555484
rect 201132 555432 201184 555484
rect 205640 555432 205692 555484
rect 264244 555432 264296 555484
rect 270132 555432 270184 555484
rect 286324 555432 286376 555484
rect 58624 554208 58676 554260
rect 74540 554208 74592 554260
rect 189908 554208 189960 554260
rect 217324 554208 217376 554260
rect 73160 554140 73212 554192
rect 106924 554140 106976 554192
rect 157248 554140 157300 554192
rect 203064 554140 203116 554192
rect 250812 554140 250864 554192
rect 319536 554140 319588 554192
rect 72424 554072 72476 554124
rect 109684 554072 109736 554124
rect 136916 554072 136968 554124
rect 202328 554072 202380 554124
rect 206376 554072 206428 554124
rect 241520 554072 241572 554124
rect 242900 554072 242952 554124
rect 316868 554072 316920 554124
rect 69572 554004 69624 554056
rect 114560 554004 114612 554056
rect 179144 554004 179196 554056
rect 269764 554004 269816 554056
rect 57336 552916 57388 552968
rect 59544 552848 59596 552900
rect 70492 552848 70544 552900
rect 71688 552848 71740 552900
rect 81716 552780 81768 552832
rect 86960 552780 87012 552832
rect 88156 552780 88208 552832
rect 88432 552780 88484 552832
rect 89628 552780 89680 552832
rect 98092 552780 98144 552832
rect 123208 552916 123260 552968
rect 122932 552848 122984 552900
rect 124036 552848 124088 552900
rect 184940 552848 184992 552900
rect 216036 552916 216088 552968
rect 251548 552916 251600 552968
rect 202144 552848 202196 552900
rect 210700 552848 210752 552900
rect 139032 552780 139084 552832
rect 208400 552780 208452 552832
rect 209228 552780 209280 552832
rect 212540 552780 212592 552832
rect 213552 552780 213604 552832
rect 213920 552780 213972 552832
rect 215024 552780 215076 552832
rect 255320 552848 255372 552900
rect 256516 552848 256568 552900
rect 259460 552916 259512 552968
rect 311164 552916 311216 552968
rect 316684 552848 316736 552900
rect 280988 552780 281040 552832
rect 67640 552712 67692 552764
rect 68836 552712 68888 552764
rect 69020 552712 69072 552764
rect 70308 552712 70360 552764
rect 75920 552712 75972 552764
rect 76748 552712 76800 552764
rect 82452 552712 82504 552764
rect 116584 552712 116636 552764
rect 125600 552712 125652 552764
rect 126888 552712 126940 552764
rect 129740 552712 129792 552764
rect 130476 552712 130528 552764
rect 142160 552712 142212 552764
rect 143356 552712 143408 552764
rect 143540 552712 143592 552764
rect 144736 552712 144788 552764
rect 154580 552712 154632 552764
rect 155500 552712 155552 552764
rect 160100 552712 160152 552764
rect 161296 552712 161348 552764
rect 164332 552712 164384 552764
rect 165528 552712 165580 552764
rect 180800 552712 180852 552764
rect 181996 552712 182048 552764
rect 189172 552712 189224 552764
rect 267004 552712 267056 552764
rect 273260 552712 273312 552764
rect 274456 552712 274508 552764
rect 293960 552712 294012 552764
rect 295248 552712 295300 552764
rect 101036 552644 101088 552696
rect 106280 552644 106332 552696
rect 107568 552644 107620 552696
rect 127624 552644 127676 552696
rect 194692 552644 194744 552696
rect 198556 552644 198608 552696
rect 278044 552644 278096 552696
rect 238668 552576 238720 552628
rect 318524 552576 318576 552628
rect 256700 552508 256752 552560
rect 257988 552508 258040 552560
rect 293132 552508 293184 552560
rect 312912 552508 312964 552560
rect 289544 552440 289596 552492
rect 312728 552440 312780 552492
rect 285956 552372 286008 552424
rect 313004 552372 313056 552424
rect 283104 552304 283156 552356
rect 315396 552304 315448 552356
rect 284116 552236 284168 552288
rect 316868 552236 316920 552288
rect 242256 552168 242308 552220
rect 315304 552168 315356 552220
rect 237932 552100 237984 552152
rect 318432 552100 318484 552152
rect 283748 552032 283800 552084
rect 287796 552032 287848 552084
rect 293776 552032 293828 552084
rect 312636 552032 312688 552084
rect 137744 551964 137796 552016
rect 139768 551964 139820 552016
rect 171324 551420 171376 551472
rect 203432 551420 203484 551472
rect 252284 551420 252336 551472
rect 318064 551420 318116 551472
rect 137836 551352 137888 551404
rect 149060 551352 149112 551404
rect 168380 551352 168432 551404
rect 200764 551352 200816 551404
rect 219164 551352 219216 551404
rect 227168 551352 227220 551404
rect 271604 551352 271656 551404
rect 317972 551352 318024 551404
rect 57704 551284 57756 551336
rect 89720 551284 89772 551336
rect 120448 551284 120500 551336
rect 129096 551284 129148 551336
rect 139400 551284 139452 551336
rect 163412 551284 163464 551336
rect 184204 551284 184256 551336
rect 281632 551284 281684 551336
rect 285220 551284 285272 551336
rect 292488 551284 292540 551336
rect 244372 551216 244424 551268
rect 318248 551216 318300 551268
rect 287336 551148 287388 551200
rect 313096 551148 313148 551200
rect 207112 551080 207164 551132
rect 210516 551080 210568 551132
rect 291660 551080 291712 551132
rect 292396 551080 292448 551132
rect 292488 551080 292540 551132
rect 312820 551080 312872 551132
rect 273076 551012 273128 551064
rect 302884 551012 302936 551064
rect 272340 550944 272392 550996
rect 318340 550944 318392 550996
rect 263048 550876 263100 550928
rect 314016 550876 314068 550928
rect 264428 550808 264480 550860
rect 318156 550808 318208 550860
rect 255872 550740 255924 550792
rect 316684 550740 316736 550792
rect 291200 550672 291252 550724
rect 292396 550672 292448 550724
rect 292488 550672 292540 550724
rect 309784 550672 309836 550724
rect 278780 550604 278832 550656
rect 301412 550604 301464 550656
rect 84844 550536 84896 550588
rect 86776 550536 86828 550588
rect 87604 550536 87656 550588
rect 91008 550536 91060 550588
rect 108304 550536 108356 550588
rect 111800 550536 111852 550588
rect 115204 550536 115256 550588
rect 116124 550536 116176 550588
rect 135444 550536 135496 550588
rect 137284 550536 137336 550588
rect 154120 550536 154172 550588
rect 157248 550536 157300 550588
rect 165620 550536 165672 550588
rect 169852 550536 169904 550588
rect 174176 550536 174228 550588
rect 179512 550536 179564 550588
rect 201408 550536 201460 550588
rect 206284 550536 206336 550588
rect 217508 550536 217560 550588
rect 219256 550536 219308 550588
rect 219532 550536 219584 550588
rect 221464 550536 221516 550588
rect 222292 550536 222344 550588
rect 225788 550536 225840 550588
rect 105544 550468 105596 550520
rect 108948 550468 109000 550520
rect 134984 550468 135036 550520
rect 146944 550468 146996 550520
rect 162676 550468 162728 550520
rect 168472 550468 168524 550520
rect 202788 550468 202840 550520
rect 208492 550468 208544 550520
rect 55128 550400 55180 550452
rect 67364 550400 67416 550452
rect 91192 550400 91244 550452
rect 96804 550400 96856 550452
rect 139860 550400 139912 550452
rect 153384 550400 153436 550452
rect 164884 550400 164936 550452
rect 173440 550400 173492 550452
rect 55036 550332 55088 550384
rect 88892 550332 88944 550384
rect 89720 550332 89772 550384
rect 117596 550332 117648 550384
rect 135168 550332 135220 550384
rect 151268 550332 151320 550384
rect 159364 550332 159416 550384
rect 167000 550332 167052 550384
rect 57796 550264 57848 550316
rect 93216 550264 93268 550316
rect 96068 550264 96120 550316
rect 98092 550264 98144 550316
rect 118976 550264 119028 550316
rect 126244 550264 126296 550316
rect 135076 550264 135128 550316
rect 157708 550264 157760 550316
rect 164148 550264 164200 550316
rect 173164 550264 173216 550316
rect 199936 550264 199988 550316
rect 205088 550264 205140 550316
rect 262312 550264 262364 550316
rect 300492 550264 300544 550316
rect 60372 550196 60424 550248
rect 95332 550196 95384 550248
rect 114008 550196 114060 550248
rect 127072 550196 127124 550248
rect 138296 550196 138348 550248
rect 157984 550196 158036 550248
rect 160744 550196 160796 550248
rect 172704 550196 172756 550248
rect 257252 550196 257304 550248
rect 301964 550196 302016 550248
rect 56508 550128 56560 550180
rect 83924 550128 83976 550180
rect 85304 550128 85356 550180
rect 120908 550128 120960 550180
rect 137928 550128 137980 550180
rect 156972 550128 157024 550180
rect 158352 550128 158404 550180
rect 182824 550128 182876 550180
rect 195612 550128 195664 550180
rect 206468 550128 206520 550180
rect 270868 550128 270920 550180
rect 319720 550128 319772 550180
rect 59268 550060 59320 550112
rect 98920 550060 98972 550112
rect 106832 550060 106884 550112
rect 124404 550060 124456 550112
rect 136548 550060 136600 550112
rect 164884 550060 164936 550112
rect 170588 550060 170640 550112
rect 200948 550060 201000 550112
rect 212172 550060 212224 550112
rect 236092 550060 236144 550112
rect 252928 550060 252980 550112
rect 319812 550060 319864 550112
rect 56416 549992 56468 550044
rect 73804 549992 73856 550044
rect 78128 549992 78180 550044
rect 121644 549992 121696 550044
rect 136456 549992 136508 550044
rect 171968 549992 172020 550044
rect 176292 549992 176344 550044
rect 213184 549992 213236 550044
rect 217968 549992 218020 550044
rect 230020 549992 230072 550044
rect 231492 549992 231544 550044
rect 238760 549992 238812 550044
rect 239404 549992 239456 550044
rect 284944 549992 284996 550044
rect 54944 549924 54996 549976
rect 99656 549924 99708 549976
rect 103980 549924 104032 549976
rect 124496 549924 124548 549976
rect 146208 549924 146260 549976
rect 201592 549924 201644 549976
rect 220084 549924 220136 549976
rect 233608 549924 233660 549976
rect 237196 549924 237248 549976
rect 284116 549924 284168 549976
rect 299572 549924 299624 549976
rect 319444 549924 319496 549976
rect 61384 549856 61436 549908
rect 116860 549856 116912 549908
rect 139308 549856 139360 549908
rect 175556 549856 175608 549908
rect 182732 549856 182784 549908
rect 242164 549856 242216 549908
rect 245844 549856 245896 549908
rect 281172 549856 281224 549908
rect 281632 549856 281684 549908
rect 303160 549856 303212 549908
rect 278044 549788 278096 549840
rect 300676 549788 300728 549840
rect 277308 549720 277360 549772
rect 300400 549720 300452 549772
rect 276572 549652 276624 549704
rect 301688 549652 301740 549704
rect 273720 549584 273772 549636
rect 301872 549584 301924 549636
rect 296720 549516 296772 549568
rect 315488 549516 315540 549568
rect 240048 549448 240100 549500
rect 266360 549448 266412 549500
rect 275928 549448 275980 549500
rect 316960 549448 317012 549500
rect 280160 549380 280212 549432
rect 61660 549312 61712 549364
rect 64972 549312 65024 549364
rect 102784 549312 102836 549364
rect 106096 549312 106148 549364
rect 108396 549312 108448 549364
rect 114652 549312 114704 549364
rect 118240 549312 118292 549364
rect 124864 549312 124916 549364
rect 131212 549312 131264 549364
rect 134524 549312 134576 549364
rect 203524 549312 203576 549364
rect 211804 549312 211856 549364
rect 243636 549312 243688 549364
rect 273260 549312 273312 549364
rect 298836 549380 298888 549432
rect 319536 549380 319588 549432
rect 284484 549312 284536 549364
rect 300216 549312 300268 549364
rect 302056 549244 302108 549296
rect 295984 548768 296036 548820
rect 315672 548768 315724 548820
rect 268752 548700 268804 548752
rect 300124 548700 300176 548752
rect 265900 548632 265952 548684
rect 301780 548632 301832 548684
rect 273260 548564 273312 548616
rect 318708 548564 318760 548616
rect 266360 548496 266412 548548
rect 318616 548496 318668 548548
rect 265164 548428 265216 548480
rect 305644 548428 305696 548480
rect 260840 548360 260892 548412
rect 304448 548360 304500 548412
rect 254400 548292 254452 548344
rect 302976 548292 303028 548344
rect 236460 548224 236512 548276
rect 301228 548224 301280 548276
rect 249432 548156 249484 548208
rect 319628 548156 319680 548208
rect 235816 548088 235868 548140
rect 247224 548088 247276 548140
rect 319444 548088 319496 548140
rect 319720 548020 319772 548072
rect 301412 547816 301464 547868
rect 317972 547816 318024 547868
rect 301228 542308 301280 542360
rect 317972 542308 318024 542360
rect 302792 539588 302844 539640
rect 311164 539588 311216 539640
rect 313004 528504 313056 528556
rect 495440 528504 495492 528556
rect 313096 528436 313148 528488
rect 476120 528436 476172 528488
rect 315672 528368 315724 528420
rect 457444 528368 457496 528420
rect 300584 528300 300636 528352
rect 430580 528300 430632 528352
rect 300676 528232 300728 528284
rect 431224 528232 431276 528284
rect 301964 528164 302016 528216
rect 431316 528164 431368 528216
rect 302056 528096 302108 528148
rect 431408 528096 431460 528148
rect 318064 528028 318116 528080
rect 430672 528028 430724 528080
rect 319904 527960 319956 528012
rect 431132 527960 431184 528012
rect 319812 527892 319864 527944
rect 430856 527892 430908 527944
rect 318524 527824 318576 527876
rect 429568 527824 429620 527876
rect 318432 527756 318484 527808
rect 428372 527756 428424 527808
rect 304264 527212 304316 527264
rect 369308 527212 369360 527264
rect 301872 527144 301924 527196
rect 396908 527144 396960 527196
rect 312912 527076 312964 527128
rect 512276 527076 512328 527128
rect 315580 527008 315632 527060
rect 500960 527008 501012 527060
rect 309784 526940 309836 526992
rect 457812 526940 457864 526992
rect 315488 526872 315540 526924
rect 459560 526872 459612 526924
rect 319536 526804 319588 526856
rect 457628 526804 457680 526856
rect 300400 526736 300452 526788
rect 430948 526736 431000 526788
rect 300216 526668 300268 526720
rect 430764 526668 430816 526720
rect 303160 526600 303212 526652
rect 431040 526600 431092 526652
rect 315396 526532 315448 526584
rect 429476 526532 429528 526584
rect 301688 526464 301740 526516
rect 414940 526464 414992 526516
rect 324872 526396 324924 526448
rect 429200 526396 429252 526448
rect 316960 526328 317012 526380
rect 351276 526328 351328 526380
rect 313924 526260 313976 526312
rect 337660 526260 337712 526312
rect 300492 526192 300544 526244
rect 328644 526192 328696 526244
rect 319628 525716 319680 525768
rect 423956 525716 424008 525768
rect 319720 525648 319772 525700
rect 305644 525580 305696 525632
rect 320088 525580 320140 525632
rect 320456 525648 320508 525700
rect 419540 525648 419592 525700
rect 333244 525580 333296 525632
rect 318248 525512 318300 525564
rect 320272 525512 320324 525564
rect 320548 525512 320600 525564
rect 405924 525512 405976 525564
rect 300124 525444 300176 525496
rect 387892 525444 387944 525496
rect 316684 525376 316736 525428
rect 320364 525376 320416 525428
rect 320640 525376 320692 525428
rect 401600 525376 401652 525428
rect 301780 525308 301832 525360
rect 383660 525308 383712 525360
rect 302884 525240 302936 525292
rect 364708 525240 364760 525292
rect 318156 525172 318208 525224
rect 374460 525172 374512 525224
rect 301596 525104 301648 525156
rect 356244 525104 356296 525156
rect 319444 525036 319496 525088
rect 360292 525036 360344 525088
rect 302976 524968 303028 525020
rect 346676 524968 346728 525020
rect 304448 524900 304500 524952
rect 342260 524900 342312 524952
rect 318340 524832 318392 524884
rect 410524 524832 410576 524884
rect 314016 524764 314068 524816
rect 320640 524764 320692 524816
rect 304356 524356 304408 524408
rect 512184 524356 512236 524408
rect 301504 524288 301556 524340
rect 488540 524288 488592 524340
rect 312820 524220 312872 524272
rect 470600 524220 470652 524272
rect 302332 523676 302384 523728
rect 578884 523676 578936 523728
rect 312636 522928 312688 522980
rect 465080 522928 465132 522980
rect 312728 522860 312780 522912
rect 457720 522860 457772 522912
rect 315304 522792 315356 522844
rect 429660 522792 429712 522844
rect 316868 522724 316920 522776
rect 427820 522724 427872 522776
rect 44088 518168 44140 518220
rect 57888 518168 57940 518220
rect 311164 515380 311216 515432
rect 580264 515380 580316 515432
rect 560944 511912 560996 511964
rect 580172 511912 580224 511964
rect 302240 495456 302292 495508
rect 520924 495456 520976 495508
rect 201516 487772 201568 487824
rect 201776 487772 201828 487824
rect 274656 487772 274708 487824
rect 274824 487772 274876 487824
rect 128360 487024 128412 487076
rect 128636 487024 128688 487076
rect 178040 487024 178092 487076
rect 178316 487024 178368 487076
rect 248512 487024 248564 487076
rect 248788 487024 248840 487076
rect 140872 486480 140924 486532
rect 199016 486480 199068 486532
rect 14464 486412 14516 486464
rect 378140 486412 378192 486464
rect 53748 485732 53800 485784
rect 74264 485732 74316 485784
rect 74356 485732 74408 485784
rect 102876 485732 102928 485784
rect 152188 485732 152240 485784
rect 209780 485732 209832 485784
rect 209872 485732 209924 485784
rect 219900 485732 219952 485784
rect 56508 485664 56560 485716
rect 89168 485664 89220 485716
rect 150440 485664 150492 485716
rect 60004 485596 60056 485648
rect 91836 485596 91888 485648
rect 149520 485596 149572 485648
rect 205640 485596 205692 485648
rect 208216 485664 208268 485716
rect 217784 485664 217836 485716
rect 208400 485596 208452 485648
rect 209780 485596 209832 485648
rect 211252 485596 211304 485648
rect 56324 485528 56376 485580
rect 88340 485528 88392 485580
rect 151268 485528 151320 485580
rect 205732 485528 205784 485580
rect 50896 485460 50948 485512
rect 79324 485460 79376 485512
rect 157708 485460 157760 485512
rect 211160 485528 211212 485580
rect 244556 485528 244608 485580
rect 356796 485528 356848 485580
rect 239680 485460 239732 485512
rect 358268 485460 358320 485512
rect 56232 485392 56284 485444
rect 90548 485392 90600 485444
rect 149428 485392 149480 485444
rect 79232 485324 79284 485376
rect 104164 485324 104216 485376
rect 157432 485324 157484 485376
rect 188344 485324 188396 485376
rect 191196 485392 191248 485444
rect 205640 485392 205692 485444
rect 209320 485392 209372 485444
rect 219072 485392 219124 485444
rect 240048 485392 240100 485444
rect 358360 485392 358412 485444
rect 68284 485256 68336 485308
rect 105544 485256 105596 485308
rect 156696 485256 156748 485308
rect 157708 485256 157760 485308
rect 157800 485256 157852 485308
rect 189264 485256 189316 485308
rect 206928 485324 206980 485376
rect 219164 485324 219216 485376
rect 234528 485324 234580 485376
rect 364984 485324 365036 485376
rect 200304 485256 200356 485308
rect 200396 485256 200448 485308
rect 55956 485188 56008 485240
rect 103336 485188 103388 485240
rect 154304 485188 154356 485240
rect 200488 485188 200540 485240
rect 209504 485256 209556 485308
rect 221740 485256 221792 485308
rect 226064 485256 226116 485308
rect 356704 485256 356756 485308
rect 217508 485188 217560 485240
rect 224224 485188 224276 485240
rect 358176 485188 358228 485240
rect 61016 485120 61068 485172
rect 116584 485120 116636 485172
rect 139216 485120 139268 485172
rect 51632 485052 51684 485104
rect 100668 485052 100720 485104
rect 110328 485052 110380 485104
rect 180064 485052 180116 485104
rect 188344 485120 188396 485172
rect 191196 485120 191248 485172
rect 193864 485052 193916 485104
rect 195336 485052 195388 485104
rect 212356 485120 212408 485172
rect 230664 485120 230716 485172
rect 366364 485120 366416 485172
rect 199936 485052 199988 485104
rect 217416 485052 217468 485104
rect 225604 485052 225656 485104
rect 362224 485052 362276 485104
rect 56416 484984 56468 485036
rect 64144 484916 64196 484968
rect 72424 484916 72476 484968
rect 73804 484916 73856 484968
rect 78036 484916 78088 484968
rect 58532 484848 58584 484900
rect 79324 484984 79376 485036
rect 84384 484984 84436 485036
rect 139400 484984 139452 485036
rect 185584 484984 185636 485036
rect 189264 484984 189316 485036
rect 201500 484984 201552 485036
rect 78220 484916 78272 484968
rect 100208 484916 100260 484968
rect 158628 484916 158680 484968
rect 197452 484916 197504 484968
rect 81716 484848 81768 484900
rect 81256 484780 81308 484832
rect 155316 484780 155368 484832
rect 157800 484780 157852 484832
rect 68376 484712 68428 484764
rect 79232 484712 79284 484764
rect 166080 484712 166132 484764
rect 204904 484848 204956 484900
rect 50988 484372 51040 484424
rect 68468 484372 68520 484424
rect 195152 484372 195204 484424
rect 197084 484372 197136 484424
rect 205916 484372 205968 484424
rect 207664 484372 207716 484424
rect 211712 484372 211764 484424
rect 212816 484372 212868 484424
rect 213368 484372 213420 484424
rect 215024 484372 215076 484424
rect 217048 484372 217100 484424
rect 218152 484372 218204 484424
rect 220176 484372 220228 484424
rect 222660 484372 222712 484424
rect 285496 484304 285548 484356
rect 285864 484236 285916 484288
rect 286140 484236 286192 484288
rect 289728 484236 289780 484288
rect 291200 484236 291252 484288
rect 291936 484236 291988 484288
rect 358084 484304 358136 484356
rect 371148 484236 371200 484288
rect 62120 484168 62172 484220
rect 62948 484168 63000 484220
rect 78680 484168 78732 484220
rect 79692 484168 79744 484220
rect 92572 484168 92624 484220
rect 93308 484168 93360 484220
rect 140780 484168 140832 484220
rect 141700 484168 141752 484220
rect 142252 484168 142304 484220
rect 142988 484168 143040 484220
rect 207112 484168 207164 484220
rect 207756 484168 207808 484220
rect 280068 484168 280120 484220
rect 366916 484168 366968 484220
rect 62212 484100 62264 484152
rect 62396 484100 62448 484152
rect 67732 484100 67784 484152
rect 68192 484100 68244 484152
rect 69020 484100 69072 484152
rect 69572 484100 69624 484152
rect 70400 484100 70452 484152
rect 70860 484100 70912 484152
rect 71872 484100 71924 484152
rect 72608 484100 72660 484152
rect 74540 484100 74592 484152
rect 74724 484100 74776 484152
rect 75920 484100 75972 484152
rect 76564 484100 76616 484152
rect 78772 484100 78824 484152
rect 78956 484100 79008 484152
rect 92480 484100 92532 484152
rect 92940 484100 92992 484152
rect 93860 484100 93912 484152
rect 94596 484100 94648 484152
rect 100760 484100 100812 484152
rect 101588 484100 101640 484152
rect 106280 484100 106332 484152
rect 106924 484100 106976 484152
rect 107660 484100 107712 484152
rect 108212 484100 108264 484152
rect 109040 484100 109092 484152
rect 109592 484100 109644 484152
rect 116032 484100 116084 484152
rect 116676 484100 116728 484152
rect 139400 484100 139452 484152
rect 140044 484100 140096 484152
rect 140872 484100 140924 484152
rect 141332 484100 141384 484152
rect 142160 484100 142212 484152
rect 142620 484100 142672 484152
rect 143540 484100 143592 484152
rect 143908 484100 143960 484152
rect 154580 484100 154632 484152
rect 155408 484100 155460 484152
rect 167092 484100 167144 484152
rect 167736 484100 167788 484152
rect 169852 484100 169904 484152
rect 170404 484100 170456 484152
rect 171140 484100 171192 484152
rect 171692 484100 171744 484152
rect 172520 484100 172572 484152
rect 173532 484100 173584 484152
rect 175280 484100 175332 484152
rect 176108 484100 176160 484152
rect 198740 484100 198792 484152
rect 198924 484100 198976 484152
rect 200212 484100 200264 484152
rect 201040 484100 201092 484152
rect 201500 484100 201552 484152
rect 202052 484100 202104 484152
rect 202880 484100 202932 484152
rect 203892 484100 203944 484152
rect 204352 484100 204404 484152
rect 205180 484100 205232 484152
rect 205732 484100 205784 484152
rect 206468 484100 206520 484152
rect 207204 484100 207256 484152
rect 207572 484100 207624 484152
rect 208400 484100 208452 484152
rect 209412 484100 209464 484152
rect 211252 484100 211304 484152
rect 211804 484100 211856 484152
rect 212632 484100 212684 484152
rect 213460 484100 213512 484152
rect 213920 484100 213972 484152
rect 214932 484100 214984 484152
rect 226340 484100 226392 484152
rect 226708 484100 226760 484152
rect 227812 484100 227864 484152
rect 228548 484100 228600 484152
rect 231860 484100 231912 484152
rect 232412 484100 232464 484152
rect 236000 484100 236052 484152
rect 236828 484100 236880 484152
rect 240232 484100 240284 484152
rect 240876 484100 240928 484152
rect 241520 484100 241572 484152
rect 242164 484100 242216 484152
rect 263692 484100 263744 484152
rect 264244 484100 264296 484152
rect 265072 484100 265124 484152
rect 265900 484100 265952 484152
rect 266360 484100 266412 484152
rect 266820 484100 266872 484152
rect 267740 484100 267792 484152
rect 268660 484100 268712 484152
rect 269212 484100 269264 484152
rect 269948 484100 270000 484152
rect 270500 484100 270552 484152
rect 271236 484100 271288 484152
rect 271972 484100 272024 484152
rect 272524 484100 272576 484152
rect 273260 484100 273312 484152
rect 273812 484100 273864 484152
rect 274640 484100 274692 484152
rect 275192 484100 275244 484152
rect 277400 484100 277452 484152
rect 278228 484100 278280 484152
rect 278780 484100 278832 484152
rect 279148 484100 279200 484152
rect 281632 484100 281684 484152
rect 282276 484100 282328 484152
rect 282920 484100 282972 484152
rect 283196 484100 283248 484152
rect 285772 484100 285824 484152
rect 286692 484100 286744 484152
rect 287060 484100 287112 484152
rect 287980 484100 288032 484152
rect 288440 484100 288492 484152
rect 288900 484100 288952 484152
rect 289912 484100 289964 484152
rect 290556 484100 290608 484152
rect 291292 484100 291344 484152
rect 291476 484100 291528 484152
rect 297364 484100 297416 484152
rect 379980 484100 380032 484152
rect 203800 484032 203852 484084
rect 209596 484032 209648 484084
rect 257988 484032 258040 484084
rect 363972 484032 364024 484084
rect 226432 483964 226484 484016
rect 227260 483964 227312 484016
rect 262128 483964 262180 484016
rect 376208 483964 376260 484016
rect 245200 483896 245252 483948
rect 369124 483896 369176 483948
rect 248328 483828 248380 483880
rect 378784 483828 378836 483880
rect 60648 483760 60700 483812
rect 80704 483760 80756 483812
rect 229744 483760 229796 483812
rect 363604 483760 363656 483812
rect 54760 483692 54812 483744
rect 117320 483692 117372 483744
rect 176936 483692 176988 483744
rect 206560 483692 206612 483744
rect 224776 483692 224828 483744
rect 370504 483692 370556 483744
rect 3424 483624 3476 483676
rect 316776 483624 316828 483676
rect 287428 483556 287480 483608
rect 297364 483556 297416 483608
rect 113272 483352 113324 483404
rect 113548 483352 113600 483404
rect 51908 482944 51960 482996
rect 98460 482944 98512 482996
rect 47860 482876 47912 482928
rect 97540 482876 97592 482928
rect 49240 482808 49292 482860
rect 98000 482808 98052 482860
rect 46664 482740 46716 482792
rect 111248 482740 111300 482792
rect 46572 482672 46624 482724
rect 111708 482672 111760 482724
rect 176016 482672 176068 482724
rect 210700 482672 210752 482724
rect 285128 482672 285180 482724
rect 359832 482672 359884 482724
rect 49332 482604 49384 482656
rect 115204 482604 115256 482656
rect 173440 482604 173492 482656
rect 209044 482604 209096 482656
rect 274824 482604 274876 482656
rect 361304 482604 361356 482656
rect 46388 482536 46440 482588
rect 112076 482536 112128 482588
rect 138480 482536 138532 482588
rect 196992 482536 197044 482588
rect 278136 482536 278188 482588
rect 369584 482536 369636 482588
rect 46296 482468 46348 482520
rect 112536 482468 112588 482520
rect 137192 482468 137244 482520
rect 198096 482468 198148 482520
rect 277308 482468 277360 482520
rect 368296 482468 368348 482520
rect 46848 482400 46900 482452
rect 115664 482400 115716 482452
rect 138848 482400 138900 482452
rect 200396 482400 200448 482452
rect 257712 482400 257764 482452
rect 362592 482400 362644 482452
rect 45928 482332 45980 482384
rect 119620 482332 119672 482384
rect 136548 482332 136600 482384
rect 203156 482332 203208 482384
rect 261760 482332 261812 482384
rect 373540 482332 373592 482384
rect 50160 482264 50212 482316
rect 131120 482264 131172 482316
rect 136272 482264 136324 482316
rect 204536 482264 204588 482316
rect 245016 482264 245068 482316
rect 360936 482264 360988 482316
rect 50436 482196 50488 482248
rect 97172 482196 97224 482248
rect 54668 482128 54720 482180
rect 96712 482128 96764 482180
rect 58808 482060 58860 482112
rect 96252 482060 96304 482112
rect 127164 482060 127216 482112
rect 127348 482060 127400 482112
rect 182364 481312 182416 481364
rect 283012 481312 283064 481364
rect 283564 481312 283616 481364
rect 294052 481312 294104 481364
rect 294236 481312 294288 481364
rect 281448 481244 281500 481296
rect 370412 481244 370464 481296
rect 192116 481176 192168 481228
rect 192300 481176 192352 481228
rect 281080 481176 281132 481228
rect 376484 481176 376536 481228
rect 180892 481108 180944 481160
rect 181076 481108 181128 481160
rect 182364 481108 182416 481160
rect 189356 481108 189408 481160
rect 203892 481108 203944 481160
rect 251180 481108 251232 481160
rect 251364 481108 251416 481160
rect 261208 481108 261260 481160
rect 366732 481108 366784 481160
rect 180524 481040 180576 481092
rect 214840 481040 214892 481092
rect 243084 481040 243136 481092
rect 365076 481040 365128 481092
rect 56876 480972 56928 481024
rect 114284 480972 114336 481024
rect 158720 480972 158772 481024
rect 159364 480972 159416 481024
rect 160284 480972 160336 481024
rect 210424 480972 210476 481024
rect 229560 480972 229612 481024
rect 360844 480972 360896 481024
rect 3608 480904 3660 480956
rect 429292 480904 429344 480956
rect 82820 480836 82872 480888
rect 83556 480836 83608 480888
rect 85580 480836 85632 480888
rect 86316 480836 86368 480888
rect 126980 480836 127032 480888
rect 127716 480836 127768 480888
rect 158812 480836 158864 480888
rect 158996 480836 159048 480888
rect 160100 480836 160152 480888
rect 160652 480836 160704 480888
rect 161572 480836 161624 480888
rect 162492 480836 162544 480888
rect 179420 480836 179472 480888
rect 179604 480836 179656 480888
rect 182272 480836 182324 480888
rect 183100 480836 183152 480888
rect 183652 480836 183704 480888
rect 184020 480836 184072 480888
rect 184940 480836 184992 480888
rect 185860 480836 185912 480888
rect 187700 480836 187752 480888
rect 188436 480836 188488 480888
rect 191932 480836 191984 480888
rect 192392 480836 192444 480888
rect 193312 480836 193364 480888
rect 193772 480836 193824 480888
rect 245660 480836 245712 480888
rect 246580 480836 246632 480888
rect 248420 480836 248472 480888
rect 249156 480836 249208 480888
rect 251272 480836 251324 480888
rect 251916 480836 251968 480888
rect 252652 480836 252704 480888
rect 253204 480836 253256 480888
rect 253940 480836 253992 480888
rect 254492 480836 254544 480888
rect 259460 480836 259512 480888
rect 259644 480836 259696 480888
rect 262220 480836 262272 480888
rect 262404 480836 262456 480888
rect 295432 480836 295484 480888
rect 295892 480836 295944 480888
rect 296720 480836 296772 480888
rect 297732 480836 297784 480888
rect 298100 480836 298152 480888
rect 298468 480836 298520 480888
rect 183560 480768 183612 480820
rect 184388 480768 184440 480820
rect 192024 480768 192076 480820
rect 192852 480768 192904 480820
rect 193220 480768 193272 480820
rect 194140 480768 194192 480820
rect 88432 480564 88484 480616
rect 89260 480564 89312 480616
rect 70492 480360 70544 480412
rect 71228 480360 71280 480412
rect 292672 480292 292724 480344
rect 293316 480292 293368 480344
rect 220820 480224 220872 480276
rect 221004 480224 221056 480276
rect 59728 480156 59780 480208
rect 130292 480156 130344 480208
rect 45468 480088 45520 480140
rect 118884 480088 118936 480140
rect 43904 480020 43956 480072
rect 117964 480020 118016 480072
rect 294604 480020 294656 480072
rect 371700 480020 371752 480072
rect 43812 479952 43864 480004
rect 117412 479952 117464 480004
rect 278872 479952 278924 480004
rect 361396 479952 361448 480004
rect 58624 479884 58676 479936
rect 132776 479884 132828 479936
rect 275652 479884 275704 479936
rect 372436 479884 372488 479936
rect 53564 479816 53616 479868
rect 131580 479816 131632 479868
rect 272064 479816 272116 479868
rect 370320 479816 370372 479868
rect 57336 479748 57388 479800
rect 135260 479748 135312 479800
rect 161664 479748 161716 479800
rect 161940 479748 161992 479800
rect 255780 479748 255832 479800
rect 356888 479748 356940 479800
rect 42524 479680 42576 479732
rect 123024 479680 123076 479732
rect 190552 479680 190604 479732
rect 191012 479680 191064 479732
rect 256700 479680 256752 479732
rect 361028 479680 361080 479732
rect 49056 479612 49108 479664
rect 130660 479612 130712 479664
rect 258448 479612 258500 479664
rect 370872 479612 370924 479664
rect 47768 479544 47820 479596
rect 129924 479544 129976 479596
rect 178316 479544 178368 479596
rect 200764 479544 200816 479596
rect 245936 479544 245988 479596
rect 371976 479544 372028 479596
rect 46112 479476 46164 479528
rect 128912 479476 128964 479528
rect 163044 479476 163096 479528
rect 206376 479476 206428 479528
rect 236460 479476 236512 479528
rect 363788 479476 363840 479528
rect 46480 479408 46532 479460
rect 116032 479408 116084 479460
rect 259460 479408 259512 479460
rect 260196 479408 260248 479460
rect 47952 479340 48004 479392
rect 116124 479340 116176 479392
rect 50344 479272 50396 479324
rect 115940 479272 115992 479324
rect 269212 478456 269264 478508
rect 357072 478456 357124 478508
rect 269396 478388 269448 478440
rect 359464 478388 359516 478440
rect 186412 478320 186464 478372
rect 216036 478320 216088 478372
rect 270868 478320 270920 478372
rect 373172 478320 373224 478372
rect 177028 478252 177080 478304
rect 209228 478252 209280 478304
rect 270592 478252 270644 478304
rect 377312 478252 377364 478304
rect 85672 478184 85724 478236
rect 85856 478184 85908 478236
rect 165068 478184 165120 478236
rect 211896 478184 211948 478236
rect 247408 478184 247460 478236
rect 376024 478184 376076 478236
rect 62304 478116 62356 478168
rect 199292 478116 199344 478168
rect 238208 478116 238260 478168
rect 378876 478116 378928 478168
rect 49148 477436 49200 477488
rect 125600 477436 125652 477488
rect 291292 477436 291344 477488
rect 362776 477436 362828 477488
rect 56600 477368 56652 477420
rect 134708 477368 134760 477420
rect 291384 477368 291436 477420
rect 368388 477368 368440 477420
rect 42616 477300 42668 477352
rect 120540 477300 120592 477352
rect 278780 477300 278832 477352
rect 364156 477300 364208 477352
rect 43996 477232 44048 477284
rect 123300 477232 123352 477284
rect 274732 477232 274784 477284
rect 364248 477232 364300 477284
rect 42432 477164 42484 477216
rect 121552 477164 121604 477216
rect 263692 477164 263744 477216
rect 366824 477164 366876 477216
rect 43628 477096 43680 477148
rect 124956 477096 125008 477148
rect 258908 477096 258960 477148
rect 365352 477096 365404 477148
rect 43720 477028 43772 477080
rect 125876 477028 125928 477080
rect 254860 477028 254912 477080
rect 365444 477028 365496 477080
rect 48964 476960 49016 477012
rect 133420 476960 133472 477012
rect 263784 476960 263836 477012
rect 376300 476960 376352 477012
rect 47676 476892 47728 476944
rect 132868 476892 132920 476944
rect 185032 476892 185084 476944
rect 212080 476892 212132 476944
rect 241704 476892 241756 476944
rect 367836 476892 367888 476944
rect 43260 476824 43312 476876
rect 143632 476824 143684 476876
rect 150440 476824 150492 476876
rect 211804 476824 211856 476876
rect 238760 476824 238812 476876
rect 373264 476824 373316 476876
rect 62212 476756 62264 476808
rect 199384 476756 199436 476808
rect 204444 476756 204496 476808
rect 217324 476756 217376 476808
rect 237472 476756 237524 476808
rect 376116 476756 376168 476808
rect 57060 476688 57112 476740
rect 128636 476688 128688 476740
rect 58440 476620 58492 476672
rect 128360 476620 128412 476672
rect 290188 475600 290240 475652
rect 363512 475600 363564 475652
rect 292764 475532 292816 475584
rect 376760 475532 376812 475584
rect 270500 475464 270552 475516
rect 375288 475464 375340 475516
rect 176660 475396 176712 475448
rect 205088 475396 205140 475448
rect 207664 475396 207716 475448
rect 217692 475396 217744 475448
rect 259644 475396 259696 475448
rect 372160 475396 372212 475448
rect 164240 475328 164292 475380
rect 218796 475328 218848 475380
rect 245752 475328 245804 475380
rect 362408 475328 362460 475380
rect 182180 474784 182232 474836
rect 182456 474784 182508 474836
rect 276020 474648 276072 474700
rect 357256 474648 357308 474700
rect 47584 474580 47636 474632
rect 65524 474580 65576 474632
rect 271972 474580 272024 474632
rect 367560 474580 367612 474632
rect 45100 474512 45152 474564
rect 68284 474512 68336 474564
rect 263600 474512 263652 474564
rect 364064 474512 364116 474564
rect 43536 474444 43588 474496
rect 68376 474444 68428 474496
rect 268108 474444 268160 474496
rect 375104 474444 375156 474496
rect 57428 474376 57480 474428
rect 103612 474376 103664 474428
rect 251364 474376 251416 474428
rect 366640 474376 366692 474428
rect 51816 474308 51868 474360
rect 99564 474308 99616 474360
rect 188068 474308 188120 474360
rect 207756 474308 207808 474360
rect 245660 474308 245712 474360
rect 366548 474308 366600 474360
rect 50252 474240 50304 474292
rect 98644 474240 98696 474292
rect 179512 474240 179564 474292
rect 214932 474240 214984 474292
rect 252744 474240 252796 474292
rect 374828 474240 374880 474292
rect 51724 474172 51776 474224
rect 99472 474172 99524 474224
rect 158904 474172 158956 474224
rect 202236 474172 202288 474224
rect 243452 474172 243504 474224
rect 366456 474172 366508 474224
rect 57796 474104 57848 474156
rect 113272 474104 113324 474156
rect 168472 474104 168524 474156
rect 214564 474104 214616 474156
rect 254032 474104 254084 474156
rect 379060 474104 379112 474156
rect 45192 474036 45244 474088
rect 104992 474036 105044 474088
rect 139492 474036 139544 474088
rect 207296 474036 207348 474088
rect 231860 474036 231912 474088
rect 363696 474036 363748 474088
rect 59360 473968 59412 474020
rect 180156 473968 180208 474020
rect 185584 473968 185636 474020
rect 205824 473968 205876 474020
rect 227812 473968 227864 474020
rect 362316 473968 362368 474020
rect 288532 473900 288584 473952
rect 369032 473900 369084 473952
rect 289912 473832 289964 473884
rect 365536 473832 365588 473884
rect 299020 473220 299072 473272
rect 367652 473220 367704 473272
rect 285956 473152 286008 473204
rect 361488 473152 361540 473204
rect 262864 473084 262916 473136
rect 370964 473084 371016 473136
rect 240140 473016 240192 473068
rect 362500 473016 362552 473068
rect 241612 472948 241664 473000
rect 374644 472948 374696 473000
rect 240232 472880 240284 472932
rect 373356 472880 373408 472932
rect 58716 472812 58768 472864
rect 110604 472812 110656 472864
rect 226432 472812 226484 472864
rect 367744 472812 367796 472864
rect 45008 472744 45060 472796
rect 105636 472744 105688 472796
rect 175372 472744 175424 472796
rect 202420 472744 202472 472796
rect 237380 472744 237432 472796
rect 378968 472744 379020 472796
rect 45284 472676 45336 472728
rect 106372 472676 106424 472728
rect 169944 472676 169996 472728
rect 214656 472676 214708 472728
rect 227720 472676 227772 472728
rect 371884 472676 371936 472728
rect 45376 472608 45428 472660
rect 106464 472608 106516 472660
rect 160376 472608 160428 472660
rect 210516 472608 210568 472660
rect 226340 472608 226392 472660
rect 370596 472608 370648 472660
rect 52276 471928 52328 471980
rect 82820 471928 82872 471980
rect 182272 471928 182324 471980
rect 205180 471928 205232 471980
rect 285772 471928 285824 471980
rect 357164 471928 357216 471980
rect 42340 471860 42392 471912
rect 74356 471860 74408 471912
rect 190644 471860 190696 471912
rect 216220 471860 216272 471912
rect 287520 471860 287572 471912
rect 359556 471860 359608 471912
rect 49608 471792 49660 471844
rect 82268 471792 82320 471844
rect 174820 471792 174872 471844
rect 200856 471792 200908 471844
rect 295524 471792 295576 471844
rect 368940 471792 368992 471844
rect 52184 471724 52236 471776
rect 84292 471724 84344 471776
rect 182364 471724 182416 471776
rect 209320 471724 209372 471776
rect 295432 471724 295484 471776
rect 370228 471724 370280 471776
rect 50068 471656 50120 471708
rect 82912 471656 82964 471708
rect 183744 471656 183796 471708
rect 210884 471656 210936 471708
rect 296260 471656 296312 471708
rect 373080 471656 373132 471708
rect 52920 471588 52972 471640
rect 85764 471588 85816 471640
rect 139400 471588 139452 471640
rect 196900 471588 196952 471640
rect 295340 471588 295392 471640
rect 376852 471588 376904 471640
rect 50804 471520 50856 471572
rect 84936 471520 84988 471572
rect 140964 471520 141016 471572
rect 200488 471520 200540 471572
rect 292672 471520 292724 471572
rect 376576 471520 376628 471572
rect 49516 471452 49568 471504
rect 83188 471452 83240 471504
rect 140872 471452 140924 471504
rect 204444 471452 204496 471504
rect 294052 471452 294104 471504
rect 379336 471452 379388 471504
rect 57704 471384 57756 471436
rect 113364 471384 113416 471436
rect 142344 471384 142396 471436
rect 207388 471384 207440 471436
rect 285864 471384 285916 471436
rect 374460 471384 374512 471436
rect 54576 471316 54628 471368
rect 102324 471316 102376 471368
rect 109224 471316 109276 471368
rect 197636 471316 197688 471368
rect 259552 471316 259604 471368
rect 369400 471316 369452 471368
rect 53104 471248 53156 471300
rect 101220 471248 101272 471300
rect 109132 471248 109184 471300
rect 201684 471248 201736 471300
rect 250536 471248 250588 471300
rect 365168 471248 365220 471300
rect 52092 471180 52144 471232
rect 81532 471180 81584 471232
rect 192300 471180 192352 471232
rect 213368 471180 213420 471232
rect 299480 471180 299532 471232
rect 368848 471180 368900 471232
rect 46204 471112 46256 471164
rect 64972 471112 65024 471164
rect 190552 471112 190604 471164
rect 211528 471112 211580 471164
rect 47492 471044 47544 471096
rect 64880 471044 64932 471096
rect 193864 470636 193916 470688
rect 201868 470636 201920 470688
rect 289820 470500 289872 470552
rect 366272 470500 366324 470552
rect 283104 470432 283156 470484
rect 359924 470432 359976 470484
rect 282920 470364 282972 470416
rect 360016 470364 360068 470416
rect 281540 470296 281592 470348
rect 359740 470296 359792 470348
rect 296812 470228 296864 470280
rect 375380 470228 375432 470280
rect 281724 470160 281776 470212
rect 367008 470160 367060 470212
rect 267832 470092 267884 470144
rect 357992 470092 358044 470144
rect 285680 470024 285732 470076
rect 377588 470024 377640 470076
rect 178040 469956 178092 470008
rect 210792 469956 210844 470008
rect 281632 469956 281684 470008
rect 373724 469956 373776 470008
rect 179420 469888 179472 469940
rect 219072 469888 219124 469940
rect 284300 469888 284352 469940
rect 377496 469888 377548 469940
rect 57612 469820 57664 469872
rect 111984 469820 112036 469872
rect 116584 469820 116636 469872
rect 199476 469820 199528 469872
rect 265256 469820 265308 469872
rect 361120 469820 361172 469872
rect 283012 469752 283064 469804
rect 357808 469752 357860 469804
rect 48228 469140 48280 469192
rect 80244 469140 80296 469192
rect 193404 469140 193456 469192
rect 215852 469140 215904 469192
rect 277492 469140 277544 469192
rect 365628 469140 365680 469192
rect 50712 469072 50764 469124
rect 78680 469072 78732 469124
rect 191932 469072 191984 469124
rect 217784 469072 217836 469124
rect 269120 469072 269172 469124
rect 358544 469072 358596 469124
rect 46020 469004 46072 469056
rect 63592 469004 63644 469056
rect 189172 469004 189224 469056
rect 215116 469004 215168 469056
rect 273444 469004 273496 469056
rect 364892 469004 364944 469056
rect 54852 468936 54904 468988
rect 85672 468936 85724 468988
rect 180984 468936 181036 468988
rect 210332 468936 210384 468988
rect 266360 468936 266412 468988
rect 359648 468936 359700 468988
rect 56048 468868 56100 468920
rect 86960 468868 87012 468920
rect 175280 468868 175332 468920
rect 212172 468868 212224 468920
rect 266452 468868 266504 468920
rect 361212 468868 361264 468920
rect 54944 468800 54996 468852
rect 87052 468800 87104 468852
rect 158812 468800 158864 468852
rect 207664 468800 207716 468852
rect 255320 468800 255372 468852
rect 358452 468800 358504 468852
rect 53196 468732 53248 468784
rect 85580 468732 85632 468784
rect 161480 468732 161532 468784
rect 215944 468732 215996 468784
rect 265164 468732 265216 468784
rect 371608 468732 371660 468784
rect 59912 468664 59964 468716
rect 92664 468664 92716 468716
rect 109040 468664 109092 468716
rect 197728 468664 197780 468716
rect 266544 468664 266596 468716
rect 375012 468664 375064 468716
rect 50620 468596 50672 468648
rect 92572 468596 92624 468648
rect 107752 468596 107804 468648
rect 199108 468596 199160 468648
rect 249800 468596 249852 468648
rect 367928 468596 367980 468648
rect 49424 468528 49476 468580
rect 93952 468528 94004 468580
rect 107844 468528 107896 468580
rect 200304 468528 200356 468580
rect 249892 468528 249944 468580
rect 372068 468528 372120 468580
rect 44824 468460 44876 468512
rect 103704 468460 103756 468512
rect 107660 468460 107712 468512
rect 203064 468460 203116 468512
rect 252652 468460 252704 468512
rect 374920 468460 374972 468512
rect 192024 468392 192076 468444
rect 214380 468392 214432 468444
rect 293960 468392 294012 468444
rect 377404 468392 377456 468444
rect 182180 468324 182232 468376
rect 202512 468324 202564 468376
rect 296720 468324 296772 468376
rect 378140 468324 378192 468376
rect 197268 468256 197320 468308
rect 211252 468256 211304 468308
rect 52920 467916 52972 467968
rect 53380 467916 53432 467968
rect 80704 467780 80756 467832
rect 178040 467780 178092 467832
rect 291200 467712 291252 467764
rect 358728 467712 358780 467764
rect 277400 467644 277452 467696
rect 362868 467644 362920 467696
rect 42708 467576 42760 467628
rect 66352 467576 66404 467628
rect 273260 467576 273312 467628
rect 362132 467576 362184 467628
rect 41328 467508 41380 467560
rect 70492 467508 70544 467560
rect 273352 467508 273404 467560
rect 369676 467508 369728 467560
rect 41236 467440 41288 467492
rect 71872 467440 71924 467492
rect 189080 467440 189132 467492
rect 202144 467440 202196 467492
rect 253940 467440 253992 467492
rect 362684 467440 362736 467492
rect 42248 467372 42300 467424
rect 73804 467372 73856 467424
rect 184940 467372 184992 467424
rect 213184 467372 213236 467424
rect 262312 467372 262364 467424
rect 372252 467372 372304 467424
rect 41144 467304 41196 467356
rect 73896 467304 73948 467356
rect 172520 467304 172572 467356
rect 204996 467304 205048 467356
rect 258080 467304 258132 467356
rect 368020 467304 368072 467356
rect 41052 467236 41104 467288
rect 93860 467236 93912 467288
rect 180156 467236 180208 467288
rect 218244 467236 218296 467288
rect 251180 467236 251232 467288
rect 363880 467236 363932 467288
rect 57520 467168 57572 467220
rect 114744 467168 114796 467220
rect 149060 467168 149112 467220
rect 212908 467168 212960 467220
rect 251272 467168 251324 467220
rect 368204 467168 368256 467220
rect 44916 467100 44968 467152
rect 106280 467100 106332 467152
rect 146300 467100 146352 467152
rect 218704 467100 218756 467152
rect 252560 467100 252612 467152
rect 379152 467100 379204 467152
rect 178040 466556 178092 466608
rect 208584 466556 208636 466608
rect 47400 466488 47452 466540
rect 190920 466420 190972 466472
rect 207020 466420 207072 466472
rect 207480 466420 207532 466472
rect 207940 466420 207992 466472
rect 339408 466556 339460 466608
rect 362960 466556 363012 466608
rect 498200 466556 498252 466608
rect 517796 466556 517848 466608
rect 218244 466488 218296 466540
rect 339776 466488 339828 466540
rect 356980 466488 357032 466540
rect 499764 466488 499816 466540
rect 338488 466420 338540 466472
rect 339408 466420 339460 466472
rect 351000 466420 351052 466472
rect 360200 466420 360252 466472
rect 362960 466420 363012 466472
rect 498200 466420 498252 466472
rect 510896 466488 510948 466540
rect 517520 466488 517572 466540
rect 517888 466420 517940 466472
rect 53656 466352 53708 466404
rect 77300 466352 77352 466404
rect 187792 466352 187844 466404
rect 206652 466352 206704 466404
rect 274640 466352 274692 466404
rect 366180 466352 366232 466404
rect 52368 466284 52420 466336
rect 75920 466284 75972 466336
rect 183560 466284 183612 466336
rect 207848 466284 207900 466336
rect 267740 466284 267792 466336
rect 371792 466284 371844 466336
rect 59268 466216 59320 466268
rect 67640 466216 67692 466268
rect 193220 466216 193272 466268
rect 217600 466216 217652 466268
rect 259460 466216 259512 466268
rect 369492 466216 369544 466268
rect 54484 466148 54536 466200
rect 63500 466148 63552 466200
rect 180892 466148 180944 466200
rect 205272 466148 205324 466200
rect 262220 466148 262272 466200
rect 376392 466148 376444 466200
rect 51540 466080 51592 466132
rect 66260 466080 66312 466132
rect 173900 466080 173952 466132
rect 203800 466080 203852 466132
rect 248604 466080 248656 466132
rect 369308 466080 369360 466132
rect 43444 466012 43496 466064
rect 60740 466012 60792 466064
rect 173992 466012 174044 466064
rect 216128 466012 216180 466064
rect 248512 466012 248564 466064
rect 370780 466012 370832 466064
rect 44732 465944 44784 465996
rect 62120 465944 62172 465996
rect 142160 465944 142212 465996
rect 197820 465944 197872 465996
rect 248420 465944 248472 465996
rect 373448 465944 373500 465996
rect 43352 465876 43404 465928
rect 60832 465876 60884 465928
rect 142252 465876 142304 465928
rect 200580 465876 200632 465928
rect 244280 465876 244332 465928
rect 370688 465876 370740 465928
rect 53656 465808 53708 465860
rect 74724 465808 74776 465860
rect 158720 465808 158772 465860
rect 218888 465808 218940 465860
rect 241520 465808 241572 465860
rect 369216 465808 369268 465860
rect 50068 465740 50120 465792
rect 50712 465740 50764 465792
rect 52000 465740 52052 465792
rect 52276 465740 52328 465792
rect 53012 465740 53064 465792
rect 100852 465740 100904 465792
rect 140780 465740 140832 465792
rect 205916 465740 205968 465792
rect 212448 465740 212500 465792
rect 220912 465740 220964 465792
rect 236000 465740 236052 465792
rect 365260 465740 365312 465792
rect 48228 465672 48280 465724
rect 69020 465672 69072 465724
rect 72424 465672 72476 465724
rect 198924 465672 198976 465724
rect 205456 465672 205508 465724
rect 221004 465672 221056 465724
rect 242900 465672 242952 465724
rect 374736 465672 374788 465724
rect 194600 465604 194652 465656
rect 213092 465604 213144 465656
rect 288440 465604 288492 465656
rect 357900 465604 357952 465656
rect 187700 465536 187752 465588
rect 200948 465536 201000 465588
rect 298100 465536 298152 465588
rect 360752 465536 360804 465588
rect 193312 465468 193364 465520
rect 203984 465468 204036 465520
rect 198924 465060 198976 465112
rect 358820 465060 358872 465112
rect 518900 465060 518952 465112
rect 196992 464992 197044 465044
rect 200672 464992 200724 465044
rect 58992 464788 59044 464840
rect 89904 464788 89956 464840
rect 191840 464788 191892 464840
rect 210240 464788 210292 464840
rect 58900 464720 58952 464772
rect 92480 464720 92532 464772
rect 190460 464720 190512 464772
rect 208952 464720 209004 464772
rect 52920 464652 52972 464704
rect 100760 464652 100812 464704
rect 127072 464652 127124 464704
rect 198004 464652 198056 464704
rect 55864 464584 55916 464636
rect 121460 464584 121512 464636
rect 126980 464584 127032 464636
rect 199568 464584 199620 464636
rect 55772 464516 55824 464568
rect 130016 464516 130068 464568
rect 180800 464516 180852 464568
rect 206744 464516 206796 464568
rect 57152 464448 57204 464500
rect 131304 464448 131356 464500
rect 186320 464448 186372 464500
rect 212264 464448 212316 464500
rect 287060 464448 287112 464500
rect 364800 464448 364852 464500
rect 54392 464380 54444 464432
rect 133972 464380 134024 464432
rect 136640 464380 136692 464432
rect 197912 464380 197964 464432
rect 271880 464380 271932 464432
rect 373632 464380 373684 464432
rect 52276 464312 52328 464364
rect 133880 464312 133932 464364
rect 136732 464312 136784 464364
rect 199200 464312 199252 464364
rect 264980 464312 265032 464364
rect 368112 464312 368164 464364
rect 207940 422900 207992 422952
rect 217968 422900 218020 422952
rect 47400 418072 47452 418124
rect 57888 418072 57940 418124
rect 207204 417392 207256 417444
rect 216680 417392 216732 417444
rect 358084 417392 358136 417444
rect 377220 417392 377272 417444
rect 44640 416780 44692 416832
rect 57244 416780 57296 416832
rect 205732 416712 205784 416764
rect 207204 416712 207256 416764
rect 208124 414808 208176 414860
rect 216864 414808 216916 414860
rect 198096 414672 198148 414724
rect 205640 414672 205692 414724
rect 207204 414672 207256 414724
rect 217048 414672 217100 414724
rect 359832 414672 359884 414724
rect 377680 414672 377732 414724
rect 48872 413992 48924 414044
rect 57888 413992 57940 414044
rect 55680 413924 55732 413976
rect 57060 413924 57112 413976
rect 204352 413924 204404 413976
rect 206836 413924 206888 413976
rect 206008 413244 206060 413296
rect 216864 413244 216916 413296
rect 48780 412768 48832 412820
rect 57888 412768 57940 412820
rect 54300 412700 54352 412752
rect 55864 412700 55916 412752
rect 357808 411884 357860 411936
rect 377128 411884 377180 411936
rect 217784 411408 217836 411460
rect 219256 411408 219308 411460
rect 47400 411272 47452 411324
rect 57888 411272 57940 411324
rect 2964 411204 3016 411256
rect 14464 411204 14516 411256
rect 51632 410796 51684 410848
rect 55864 410796 55916 410848
rect 206836 410524 206888 410576
rect 216680 410524 216732 410576
rect 216956 410524 217008 410576
rect 360016 410524 360068 410576
rect 377220 410524 377272 410576
rect 377404 410252 377456 410304
rect 379244 410252 379296 410304
rect 51632 409844 51684 409896
rect 56968 409844 57020 409896
rect 359924 409096 359976 409148
rect 377404 409096 377456 409148
rect 52368 408484 52420 408536
rect 57888 408484 57940 408536
rect 216680 407464 216732 407516
rect 217048 407464 217100 407516
rect 216772 398216 216824 398268
rect 216680 398012 216732 398064
rect 198096 397536 198148 397588
rect 199016 397536 199068 397588
rect 198188 396788 198240 396840
rect 199568 396788 199620 396840
rect 520924 396720 520976 396772
rect 580356 396720 580408 396772
rect 216680 392028 216732 392080
rect 217048 392028 217100 392080
rect 43260 391892 43312 391944
rect 57888 391892 57940 391944
rect 209504 391892 209556 391944
rect 216680 391892 216732 391944
rect 359740 391892 359792 391944
rect 376944 391892 376996 391944
rect 207020 390464 207072 390516
rect 216680 390464 216732 390516
rect 360200 390464 360252 390516
rect 376944 390464 376996 390516
rect 57428 390328 57480 390380
rect 57428 390056 57480 390108
rect 44088 389784 44140 389836
rect 57612 389784 57664 389836
rect 206284 389172 206336 389224
rect 207020 389172 207072 389224
rect 358084 389172 358136 389224
rect 360200 389172 360252 389224
rect 46112 389104 46164 389156
rect 57612 389104 57664 389156
rect 203892 389104 203944 389156
rect 216680 389104 216732 389156
rect 359648 389104 359700 389156
rect 376944 389104 376996 389156
rect 56784 388764 56836 388816
rect 59544 388764 59596 388816
rect 57888 388424 57940 388476
rect 58440 388424 58492 388476
rect 57336 388356 57388 388408
rect 57520 388356 57572 388408
rect 216772 388356 216824 388408
rect 217048 388356 217100 388408
rect 57244 387744 57296 387796
rect 58532 387744 58584 387796
rect 372988 382236 373040 382288
rect 376760 382236 376812 382288
rect 57428 381896 57480 381948
rect 59360 381896 59412 381948
rect 55956 380944 56008 380996
rect 59452 380944 59504 380996
rect 197176 380944 197228 380996
rect 198188 380944 198240 380996
rect 57888 380876 57940 380928
rect 60740 380876 60792 380928
rect 196992 380876 197044 380928
rect 198004 380876 198056 380928
rect 198280 380876 198332 380928
rect 199108 380876 199160 380928
rect 217600 380876 217652 380928
rect 276020 380876 276072 380928
rect 376760 380876 376812 380928
rect 421748 380876 421800 380928
rect 54300 380808 54352 380860
rect 56600 380808 56652 380860
rect 48872 380740 48924 380792
rect 216680 380808 216732 380860
rect 48780 380604 48832 380656
rect 216864 380740 216916 380792
rect 364800 380740 364852 380792
rect 379520 380740 379572 380792
rect 51632 380536 51684 380588
rect 216956 380672 217008 380724
rect 373816 380672 373868 380724
rect 378140 380672 378192 380724
rect 434352 380672 434404 380724
rect 155960 380604 156012 380656
rect 204444 380604 204496 380656
rect 360752 380604 360804 380656
rect 376668 380604 376720 380656
rect 377312 380604 377364 380656
rect 425980 380604 426032 380656
rect 158536 380536 158588 380588
rect 205916 380536 205968 380588
rect 207020 380536 207072 380588
rect 213736 380536 213788 380588
rect 373632 380536 373684 380588
rect 433616 380536 433668 380588
rect 58624 380468 58676 380520
rect 105820 380468 105872 380520
rect 138480 380468 138532 380520
rect 200396 380468 200448 380520
rect 202880 380468 202932 380520
rect 213828 380468 213880 380520
rect 359464 380468 359516 380520
rect 421104 380468 421156 380520
rect 59544 380400 59596 380452
rect 118332 380400 118384 380452
rect 135904 380400 135956 380452
rect 200672 380400 200724 380452
rect 202972 380400 203024 380452
rect 274640 380400 274692 380452
rect 370320 380400 370372 380452
rect 436008 380400 436060 380452
rect 52276 380332 52328 380384
rect 113548 380332 113600 380384
rect 123576 380332 123628 380384
rect 204536 380332 204588 380384
rect 208400 380332 208452 380384
rect 218152 380332 218204 380384
rect 367560 380332 367612 380384
rect 438492 380332 438544 380384
rect 48964 380264 49016 380316
rect 110972 380264 111024 380316
rect 148600 380264 148652 380316
rect 196900 380264 196952 380316
rect 201040 380264 201092 380316
rect 295340 380264 295392 380316
rect 369676 380264 369728 380316
rect 440884 380264 440936 380316
rect 58532 380196 58584 380248
rect 120908 380196 120960 380248
rect 133512 380196 133564 380248
rect 199200 380196 199252 380248
rect 200212 380196 200264 380248
rect 301504 380196 301556 380248
rect 364892 380196 364944 380248
rect 443460 380196 443512 380248
rect 54392 380128 54444 380180
rect 115940 380128 115992 380180
rect 128360 380128 128412 380180
rect 197912 380128 197964 380180
rect 201776 380128 201828 380180
rect 311808 380128 311860 380180
rect 365628 380128 365680 380180
rect 465908 380128 465960 380180
rect 160928 380060 160980 380112
rect 207388 380060 207440 380112
rect 166080 379992 166132 380044
rect 200580 379992 200632 380044
rect 213828 379992 213880 380044
rect 236000 379992 236052 380044
rect 366272 379992 366324 380044
rect 55680 379924 55732 379976
rect 59636 379924 59688 379976
rect 163504 379924 163556 379976
rect 197820 379924 197872 379976
rect 215300 379924 215352 379976
rect 216404 379924 216456 379976
rect 237104 379924 237156 379976
rect 239956 379924 240008 379976
rect 259460 379924 259512 379976
rect 212540 379856 212592 379908
rect 217784 379856 217836 379908
rect 218152 379856 218204 379908
rect 218336 379856 218388 379908
rect 244280 379856 244332 379908
rect 213736 379788 213788 379840
rect 243084 379788 243136 379840
rect 215024 379720 215076 379772
rect 207020 379652 207072 379704
rect 208308 379652 208360 379704
rect 209412 379652 209464 379704
rect 212724 379652 212776 379704
rect 220728 379720 220780 379772
rect 254492 379720 254544 379772
rect 379520 379788 379572 379840
rect 379888 379788 379940 379840
rect 408684 379788 408736 379840
rect 381084 379720 381136 379772
rect 413468 379720 413520 379772
rect 204260 379516 204312 379568
rect 215300 379516 215352 379568
rect 216956 379516 217008 379568
rect 217600 379516 217652 379568
rect 256976 379652 257028 379704
rect 371056 379652 371108 379704
rect 376852 379652 376904 379704
rect 377404 379652 377456 379704
rect 379244 379652 379296 379704
rect 380900 379652 380952 379704
rect 425244 379652 425296 379704
rect 217784 379584 217836 379636
rect 219716 379584 219768 379636
rect 220728 379584 220780 379636
rect 255872 379584 255924 379636
rect 376576 379584 376628 379636
rect 422852 379584 422904 379636
rect 221832 379516 221884 379568
rect 265256 379516 265308 379568
rect 376668 379516 376720 379568
rect 436928 379516 436980 379568
rect 86592 379448 86644 379500
rect 208400 379448 208452 379500
rect 220636 379448 220688 379500
rect 47768 379380 47820 379432
rect 88340 379380 88392 379432
rect 92388 379380 92440 379432
rect 212816 379380 212868 379432
rect 213828 379380 213880 379432
rect 215392 379380 215444 379432
rect 219440 379380 219492 379432
rect 273260 379380 273312 379432
rect 274640 379448 274692 379500
rect 323308 379448 323360 379500
rect 368848 379448 368900 379500
rect 439044 379448 439096 379500
rect 275652 379380 275704 379432
rect 295340 379380 295392 379432
rect 310980 379380 311032 379432
rect 311808 379380 311860 379432
rect 315764 379380 315816 379432
rect 377404 379380 377456 379432
rect 427452 379380 427504 379432
rect 88800 379312 88852 379364
rect 209780 379312 209832 379364
rect 211068 379312 211120 379364
rect 220728 379312 220780 379364
rect 274364 379312 274416 379364
rect 301504 379312 301556 379364
rect 313372 379312 313424 379364
rect 375012 379312 375064 379364
rect 408316 379312 408368 379364
rect 55772 379244 55824 379296
rect 90640 379244 90692 379296
rect 90732 379244 90784 379296
rect 209872 379244 209924 379296
rect 219624 379244 219676 379296
rect 220544 379244 220596 379296
rect 91376 379176 91428 379228
rect 59728 379108 59780 379160
rect 93492 379108 93544 379160
rect 93584 379108 93636 379160
rect 195980 379108 196032 379160
rect 47676 379040 47728 379092
rect 108212 379040 108264 379092
rect 112352 379040 112404 379092
rect 205916 379040 205968 379092
rect 213828 379176 213880 379228
rect 220820 379176 220872 379228
rect 221924 379176 221976 379228
rect 211068 379108 211120 379160
rect 219440 379108 219492 379160
rect 220176 379108 220228 379160
rect 220452 379108 220504 379160
rect 211436 379040 211488 379092
rect 221556 379040 221608 379092
rect 53564 378972 53616 379024
rect 101036 378972 101088 379024
rect 195980 378972 196032 379024
rect 197268 378972 197320 379024
rect 220912 378972 220964 379024
rect 222108 378972 222160 379024
rect 57152 378904 57204 378956
rect 103520 378904 103572 378956
rect 205732 378904 205784 378956
rect 206836 378904 206888 378956
rect 219532 378904 219584 378956
rect 220728 378904 220780 378956
rect 371148 378972 371200 379024
rect 381268 378972 381320 379024
rect 247592 378904 247644 378956
rect 357900 378904 357952 378956
rect 379520 378904 379572 378956
rect 50160 378836 50212 378888
rect 98184 378836 98236 378888
rect 111248 378836 111300 378888
rect 199016 378836 199068 378888
rect 219164 378836 219216 378888
rect 245384 378836 245436 378888
rect 373724 378836 373776 378888
rect 396172 378836 396224 378888
rect 108856 378768 108908 378820
rect 208216 378768 208268 378820
rect 268660 378768 268712 378820
rect 359556 378768 359608 378820
rect 375196 378768 375248 378820
rect 379704 378768 379756 378820
rect 379980 378768 380032 378820
rect 405740 378768 405792 378820
rect 49056 378632 49108 378684
rect 96068 378632 96120 378684
rect 115848 378632 115900 378684
rect 213460 378700 213512 378752
rect 219808 378700 219860 378752
rect 220636 378700 220688 378752
rect 220176 378632 220228 378684
rect 248604 378632 248656 378684
rect 46204 378564 46256 378616
rect 46940 378564 46992 378616
rect 85488 378564 85540 378616
rect 213644 378564 213696 378616
rect 219164 378564 219216 378616
rect 221096 378564 221148 378616
rect 221556 378564 221608 378616
rect 251180 378564 251232 378616
rect 47584 378496 47636 378548
rect 49056 378496 49108 378548
rect 114468 378496 114520 378548
rect 205732 378496 205784 378548
rect 220544 378496 220596 378548
rect 250076 378496 250128 378548
rect 374552 378496 374604 378548
rect 375012 378496 375064 378548
rect 396080 378496 396132 378548
rect 199016 378428 199068 378480
rect 209596 378428 209648 378480
rect 271052 378428 271104 378480
rect 381268 378428 381320 378480
rect 412364 378428 412416 378480
rect 208400 378360 208452 378412
rect 211620 378360 211672 378412
rect 245660 378360 245712 378412
rect 379520 378360 379572 378412
rect 379796 378360 379848 378412
rect 411260 378360 411312 378412
rect 113456 378292 113508 378344
rect 215392 378292 215444 378344
rect 221924 378292 221976 378344
rect 252284 378292 252336 378344
rect 342260 378292 342312 378344
rect 343180 378292 343232 378344
rect 359372 378292 359424 378344
rect 49056 378224 49108 378276
rect 81440 378224 81492 378276
rect 205916 378224 205968 378276
rect 206928 378224 206980 378276
rect 211712 378224 211764 378276
rect 271972 378224 272024 378276
rect 276020 378224 276072 378276
rect 277032 378224 277084 378276
rect 356612 378224 356664 378276
rect 375196 378292 375248 378344
rect 407580 378292 407632 378344
rect 439044 378292 439096 378344
rect 516600 378292 516652 378344
rect 503076 378224 503128 378276
rect 517612 378224 517664 378276
rect 580264 378224 580316 378276
rect 46940 378156 46992 378208
rect 80336 378156 80388 378208
rect 87696 378156 87748 378208
rect 219808 378156 219860 378208
rect 220452 378156 220504 378208
rect 222108 378156 222160 378208
rect 253388 378156 253440 378208
rect 273260 378156 273312 378208
rect 303068 378156 303120 378208
rect 343548 378156 343600 378208
rect 503536 378156 503588 378208
rect 517704 378156 517756 378208
rect 580172 378156 580224 378208
rect 196716 378088 196768 378140
rect 287612 378088 287664 378140
rect 367008 378088 367060 378140
rect 374552 378088 374604 378140
rect 216772 378020 216824 378072
rect 217324 378020 217376 378072
rect 217508 378020 217560 378072
rect 308404 378020 308456 378072
rect 357256 378020 357308 378072
rect 458364 378020 458416 378072
rect 43352 377952 43404 378004
rect 199660 377952 199712 378004
rect 201592 377952 201644 378004
rect 318340 377952 318392 378004
rect 366180 377952 366232 378004
rect 452752 377952 452804 378004
rect 44732 377884 44784 377936
rect 183468 377884 183520 377936
rect 198832 377884 198884 377936
rect 300860 377884 300912 377936
rect 361304 377884 361356 377936
rect 448152 377884 448204 377936
rect 54484 377816 54536 377868
rect 182272 377816 182324 377868
rect 197544 377816 197596 377868
rect 298100 377816 298152 377868
rect 364248 377816 364300 377868
rect 451004 377816 451056 377868
rect 197452 377748 197504 377800
rect 295892 377748 295944 377800
rect 362132 377748 362184 377800
rect 445852 377748 445904 377800
rect 197360 377680 197412 377732
rect 293316 377680 293368 377732
rect 372436 377680 372488 377732
rect 455512 377680 455564 377732
rect 196808 377612 196860 377664
rect 290924 377612 290976 377664
rect 357072 377612 357124 377664
rect 423404 377612 423456 377664
rect 196624 377544 196676 377596
rect 285956 377544 286008 377596
rect 357992 377544 358044 377596
rect 410616 377544 410668 377596
rect 143632 377476 143684 377528
rect 205824 377476 205876 377528
rect 217416 377476 217468 377528
rect 305736 377476 305788 377528
rect 361488 377476 361540 377528
rect 371148 377476 371200 377528
rect 375104 377476 375156 377528
rect 413100 377476 413152 377528
rect 197084 377408 197136 377460
rect 277860 377408 277912 377460
rect 363512 377408 363564 377460
rect 379980 377408 380032 377460
rect 414572 377408 414624 377460
rect 146024 377340 146076 377392
rect 207296 377340 207348 377392
rect 212356 377340 212408 377392
rect 280804 377340 280856 377392
rect 371148 377340 371200 377392
rect 402980 377340 403032 377392
rect 44640 377272 44692 377324
rect 217324 377272 217376 377324
rect 369032 377272 369084 377324
rect 379244 377272 379296 377324
rect 409972 377272 410024 377324
rect 141056 377204 141108 377256
rect 201868 377204 201920 377256
rect 364156 377204 364208 377256
rect 474740 377204 474792 377256
rect 153568 377136 153620 377188
rect 200488 377136 200540 377188
rect 150992 377068 151044 377120
rect 198188 377068 198240 377120
rect 47400 377000 47452 377052
rect 217692 377000 217744 377052
rect 77208 376660 77260 376712
rect 204260 376660 204312 376712
rect 213092 376660 213144 376712
rect 283012 376660 283064 376712
rect 361396 376660 361448 376712
rect 473452 376660 473504 376712
rect 201500 376592 201552 376644
rect 320916 376592 320968 376644
rect 366916 376592 366968 376644
rect 477592 376592 477644 376644
rect 125968 376524 126020 376576
rect 203156 376524 203208 376576
rect 203984 376524 204036 376576
rect 273444 376524 273496 376576
rect 362868 376524 362920 376576
rect 470876 376524 470928 376576
rect 97724 376456 97776 376508
rect 214472 376456 214524 376508
rect 215024 376456 215076 376508
rect 215852 376456 215904 376508
rect 270960 376456 271012 376508
rect 376484 376456 376536 376508
rect 483388 376456 483440 376508
rect 210240 376388 210292 376440
rect 263600 376388 263652 376440
rect 369584 376388 369636 376440
rect 467932 376388 467984 376440
rect 214380 376320 214432 376372
rect 268108 376320 268160 376372
rect 368296 376320 368348 376372
rect 463516 376320 463568 376372
rect 131028 376252 131080 376304
rect 205640 376252 205692 376304
rect 213368 376252 213420 376304
rect 260932 376252 260984 376304
rect 358544 376252 358596 376304
rect 418252 376252 418304 376304
rect 211528 376184 211580 376236
rect 258356 376184 258408 376236
rect 375288 376184 375340 376236
rect 430672 376184 430724 376236
rect 94688 376116 94740 376168
rect 212540 376116 212592 376168
rect 214012 376116 214064 376168
rect 216312 376116 216364 376168
rect 219256 376116 219308 376168
rect 265348 376116 265400 376168
rect 373172 376116 373224 376168
rect 428188 376116 428240 376168
rect 202144 376048 202196 376100
rect 248236 376048 248288 376100
rect 371792 376048 371844 376100
rect 416044 376048 416096 376100
rect 216220 375980 216272 376032
rect 255964 375980 256016 376032
rect 365536 375980 365588 376032
rect 374552 375980 374604 376032
rect 415400 375980 415452 376032
rect 208952 375912 209004 375964
rect 253572 375912 253624 375964
rect 374460 375912 374512 375964
rect 377312 375912 377364 375964
rect 403624 375912 403676 375964
rect 99472 375844 99524 375896
rect 214012 375844 214064 375896
rect 215116 375844 215168 375896
rect 250628 375844 250680 375896
rect 104072 375708 104124 375760
rect 216588 375708 216640 375760
rect 217232 375708 217284 375760
rect 100760 375640 100812 375692
rect 216496 375640 216548 375692
rect 216312 375572 216364 375624
rect 239956 375776 240008 375828
rect 101956 375300 102008 375352
rect 213920 375300 213972 375352
rect 218060 375300 218112 375352
rect 218244 375300 218296 375352
rect 219348 375300 219400 375352
rect 266360 375300 266412 375352
rect 215116 375232 215168 375284
rect 215484 375232 215536 375284
rect 262772 375232 262824 375284
rect 107568 375164 107620 375216
rect 207020 375164 207072 375216
rect 208308 375164 208360 375216
rect 279148 375164 279200 375216
rect 357072 375368 357124 375420
rect 374368 375368 374420 375420
rect 375472 375368 375524 375420
rect 368940 375300 368992 375352
rect 369584 375300 369636 375352
rect 428280 375300 428332 375352
rect 373080 375232 373132 375284
rect 431132 375232 431184 375284
rect 367652 375164 367704 375216
rect 370044 375164 370096 375216
rect 375472 375164 375524 375216
rect 432236 375164 432288 375216
rect 213920 375096 213972 375148
rect 217508 375096 217560 375148
rect 261668 375096 261720 375148
rect 379336 375096 379388 375148
rect 423956 375096 424008 375148
rect 106464 375028 106516 375080
rect 218060 375028 218112 375080
rect 375564 375028 375616 375080
rect 376576 375028 376628 375080
rect 405372 375028 405424 375080
rect 368388 374960 368440 375012
rect 375748 374960 375800 375012
rect 416964 374960 417016 375012
rect 362776 374892 362828 374944
rect 377128 374892 377180 374944
rect 418160 374892 418212 374944
rect 358728 374824 358780 374876
rect 376484 374824 376536 374876
rect 418344 374824 418396 374876
rect 207020 374756 207072 374808
rect 208124 374756 208176 374808
rect 217876 374756 217928 374808
rect 102968 374688 103020 374740
rect 215116 374688 215168 374740
rect 357164 374756 357216 374808
rect 375564 374756 375616 374808
rect 267556 374688 267608 374740
rect 371700 374688 371752 374740
rect 378140 374756 378192 374808
rect 426440 374756 426492 374808
rect 183468 374620 183520 374672
rect 197360 374620 197412 374672
rect 342260 374620 342312 374672
rect 370228 374620 370280 374672
rect 372436 374620 372488 374672
rect 429384 374688 429436 374740
rect 370044 374484 370096 374536
rect 370412 374484 370464 374536
rect 437756 374620 437808 374672
rect 199384 371832 199436 371884
rect 199936 371832 199988 371884
rect 359188 371832 359240 371884
rect 359188 371220 359240 371272
rect 359464 371220 359516 371272
rect 199476 370472 199528 370524
rect 359096 370472 359148 370524
rect 359832 370472 359884 370524
rect 518992 370472 519044 370524
rect 199660 369112 199712 369164
rect 199844 369112 199896 369164
rect 359096 369112 359148 369164
rect 359832 369112 359884 369164
rect 199568 366324 199620 366376
rect 359004 366324 359056 366376
rect 519268 366324 519320 366376
rect 519636 366324 519688 366376
rect 359188 364964 359240 365016
rect 359556 364964 359608 365016
rect 518900 364964 518952 365016
rect 519084 364964 519136 365016
rect 359464 363604 359516 363656
rect 519176 363604 519228 363656
rect 199752 362176 199804 362228
rect 358912 362176 358964 362228
rect 359188 362176 359240 362228
rect 519452 362176 519504 362228
rect 202604 360204 202656 360256
rect 206284 360204 206336 360256
rect 500776 359660 500828 359712
rect 518072 359660 518124 359712
rect 197452 359524 197504 359576
rect 208584 359524 208636 359576
rect 339868 359524 339920 359576
rect 356980 359524 357032 359576
rect 357164 359524 357216 359576
rect 498936 359524 498988 359576
rect 517980 359524 518032 359576
rect 190920 359456 190972 359508
rect 201500 359456 201552 359508
rect 202604 359456 202656 359508
rect 351736 359456 351788 359508
rect 358084 359456 358136 359508
rect 360200 359252 360252 359304
rect 362960 359252 363012 359304
rect 179696 358844 179748 358896
rect 178592 358776 178644 358828
rect 197452 358776 197504 358828
rect 3332 358708 3384 358760
rect 18604 358708 18656 358760
rect 55956 358708 56008 358760
rect 59452 358708 59504 358760
rect 342260 358844 342312 358896
rect 343548 358844 343600 358896
rect 358544 358844 358596 358896
rect 338488 358776 338540 358828
rect 360200 358776 360252 358828
rect 510896 358776 510948 358828
rect 517520 358776 517572 358828
rect 198096 358708 198148 358760
rect 203892 358708 203944 358760
rect 218520 358708 218572 358760
rect 221372 358708 221424 358760
rect 379428 358708 379480 358760
rect 380992 358708 381044 358760
rect 219256 358640 219308 358692
rect 220912 358640 220964 358692
rect 375288 358640 375340 358692
rect 381084 358640 381136 358692
rect 217048 358572 217100 358624
rect 220820 358572 220872 358624
rect 214380 358504 214432 358556
rect 221004 358504 221056 358556
rect 219164 358232 219216 358284
rect 221096 358232 221148 358284
rect 215668 358096 215720 358148
rect 221188 358096 221240 358148
rect 182824 358028 182876 358080
rect 201592 358028 201644 358080
rect 342260 358028 342312 358080
rect 377036 357960 377088 358012
rect 381268 357960 381320 358012
rect 57152 357824 57204 357876
rect 59360 357824 59412 357876
rect 378692 357824 378744 357876
rect 380900 357824 380952 357876
rect 215852 357484 215904 357536
rect 221280 357484 221332 357536
rect 375840 357484 375892 357536
rect 381176 357484 381228 357536
rect 58624 357348 58676 357400
rect 60740 357348 60792 357400
rect 55128 303900 55180 303952
rect 56600 303900 56652 303952
rect 46296 303560 46348 303612
rect 57336 303560 57388 303612
rect 57612 303560 57664 303612
rect 46388 300772 46440 300824
rect 56968 300772 57020 300824
rect 57428 300772 57480 300824
rect 520188 288396 520240 288448
rect 580264 288396 580316 288448
rect 518992 287036 519044 287088
rect 519452 287036 519504 287088
rect 580356 287036 580408 287088
rect 200948 284248 201000 284300
rect 216680 284248 216732 284300
rect 361212 284248 361264 284300
rect 376944 284248 376996 284300
rect 201500 282820 201552 282872
rect 216680 282820 216732 282872
rect 368204 282820 368256 282872
rect 376760 282820 376812 282872
rect 203800 282752 203852 282804
rect 216772 282752 216824 282804
rect 55128 282208 55180 282260
rect 58716 282208 58768 282260
rect 51632 282140 51684 282192
rect 58532 282140 58584 282192
rect 358084 282140 358136 282192
rect 376944 282140 376996 282192
rect 44088 281460 44140 281512
rect 57244 281460 57296 281512
rect 57520 281460 57572 281512
rect 374460 274728 374512 274780
rect 375012 274728 375064 274780
rect 212908 274660 212960 274712
rect 215392 274660 215444 274712
rect 219348 273572 219400 273624
rect 219900 273572 219952 273624
rect 266360 273572 266412 273624
rect 55864 273504 55916 273556
rect 110972 273504 111024 273556
rect 200856 273504 200908 273556
rect 250720 273504 250772 273556
rect 44824 273436 44876 273488
rect 133420 273436 133472 273488
rect 215392 273436 215444 273488
rect 273352 273436 273404 273488
rect 370320 273436 370372 273488
rect 379336 273436 379388 273488
rect 45192 273368 45244 273420
rect 135904 273368 135956 273420
rect 213460 273368 213512 273420
rect 215024 273368 215076 273420
rect 275744 273368 275796 273420
rect 369032 273368 369084 273420
rect 378140 273368 378192 273420
rect 378600 273368 378652 273420
rect 45100 273300 45152 273352
rect 138480 273300 138532 273352
rect 215760 273300 215812 273352
rect 278044 273300 278096 273352
rect 362684 273300 362736 273352
rect 421104 273300 421156 273352
rect 45008 273232 45060 273284
rect 140872 273232 140924 273284
rect 205272 273232 205324 273284
rect 283472 273232 283524 273284
rect 369400 273232 369452 273284
rect 451004 273232 451056 273284
rect 371148 273164 371200 273216
rect 375196 273164 375248 273216
rect 379336 273164 379388 273216
rect 423772 273164 423824 273216
rect 53840 273096 53892 273148
rect 100760 273096 100812 273148
rect 378600 273096 378652 273148
rect 426440 273096 426492 273148
rect 365444 273028 365496 273080
rect 423404 273028 423456 273080
rect 42524 272824 42576 272876
rect 60832 272960 60884 273012
rect 210332 272960 210384 273012
rect 288164 272960 288216 273012
rect 372344 272960 372396 273012
rect 373172 272960 373224 273012
rect 431132 272960 431184 273012
rect 58624 272892 58676 272944
rect 61108 272892 61160 272944
rect 61476 272892 61528 272944
rect 206744 272892 206796 272944
rect 285956 272892 286008 272944
rect 358452 272892 358504 272944
rect 425980 272892 426032 272944
rect 59636 272824 59688 272876
rect 60740 272824 60792 272876
rect 61752 272824 61804 272876
rect 209320 272824 209372 272876
rect 290924 272824 290976 272876
rect 356888 272824 356940 272876
rect 428188 272824 428240 272876
rect 50436 272756 50488 272808
rect 90732 272756 90784 272808
rect 210884 272756 210936 272808
rect 300860 272756 300912 272808
rect 370964 272756 371016 272808
rect 468484 272756 468536 272808
rect 47860 272688 47912 272740
rect 93676 272688 93728 272740
rect 202512 272688 202564 272740
rect 293316 272688 293368 272740
rect 376300 272688 376352 272740
rect 473452 272688 473504 272740
rect 49240 272620 49292 272672
rect 95884 272620 95936 272672
rect 205180 272620 205232 272672
rect 298468 272620 298520 272672
rect 364064 272620 364116 272672
rect 470876 272620 470928 272672
rect 51908 272552 51960 272604
rect 98460 272552 98512 272604
rect 207848 272552 207900 272604
rect 305828 272552 305880 272604
rect 366824 272552 366876 272604
rect 475844 272552 475896 272604
rect 45284 272484 45336 272536
rect 143540 272484 143592 272536
rect 208216 272484 208268 272536
rect 210884 272484 210936 272536
rect 212264 272484 212316 272536
rect 320916 272484 320968 272536
rect 368112 272484 368164 272536
rect 478420 272484 478472 272536
rect 46664 272416 46716 272468
rect 47492 272416 47544 272468
rect 46572 272348 46624 272400
rect 47676 272348 47728 272400
rect 58532 272416 58584 272468
rect 59728 272416 59780 272468
rect 99380 272416 99432 272468
rect 374552 272416 374604 272468
rect 396724 272416 396776 272468
rect 76012 272348 76064 272400
rect 65340 272280 65392 272332
rect 95976 272280 96028 272332
rect 67364 272212 67416 272264
rect 96988 272212 97040 272264
rect 46756 272144 46808 272196
rect 46940 272144 46992 272196
rect 60832 272144 60884 272196
rect 94228 272144 94280 272196
rect 53932 272076 53984 272128
rect 86960 272076 87012 272128
rect 49332 272008 49384 272060
rect 82820 272008 82872 272060
rect 83464 272008 83516 272060
rect 98000 272008 98052 272060
rect 47676 271940 47728 271992
rect 75920 271940 75972 271992
rect 213736 271940 213788 271992
rect 216220 271940 216272 271992
rect 236000 271940 236052 271992
rect 421564 271940 421616 271992
rect 437940 271940 437992 271992
rect 98644 271872 98696 271924
rect 100760 271872 100812 271924
rect 114468 271872 114520 271924
rect 127624 271872 127676 271924
rect 210884 271872 210936 271924
rect 268200 271872 268252 271924
rect 356980 271872 357032 271924
rect 359372 271872 359424 271924
rect 43536 271804 43588 271856
rect 129740 271804 129792 271856
rect 151360 271804 151412 271856
rect 198004 271804 198056 271856
rect 213184 271804 213236 271856
rect 313280 271804 313332 271856
rect 343548 271804 343600 271856
rect 358544 271804 358596 271856
rect 360292 271872 360344 271924
rect 374460 271872 374512 271924
rect 375196 271872 375248 271924
rect 402980 271872 403032 271924
rect 366732 271804 366784 271856
rect 455788 271804 455840 271856
rect 42340 271736 42392 271788
rect 123208 271736 123260 271788
rect 157248 271736 157300 271788
rect 203064 271736 203116 271788
rect 212080 271736 212132 271788
rect 307760 271736 307812 271788
rect 373540 271736 373592 271788
rect 458180 271736 458232 271788
rect 42432 271668 42484 271720
rect 53840 271668 53892 271720
rect 54392 271668 54444 271720
rect 57152 271668 57204 271720
rect 128360 271668 128412 271720
rect 154488 271668 154540 271720
rect 200304 271668 200356 271720
rect 200764 271668 200816 271720
rect 268016 271668 268068 271720
rect 369492 271668 369544 271720
rect 452660 271668 452712 271720
rect 46480 271600 46532 271652
rect 53932 271600 53984 271652
rect 55956 271600 56008 271652
rect 125600 271600 125652 271652
rect 158628 271600 158680 271652
rect 201684 271600 201736 271652
rect 214840 271600 214892 271652
rect 280160 271600 280212 271652
rect 365352 271600 365404 271652
rect 445760 271600 445812 271652
rect 54576 271532 54628 271584
rect 120080 271532 120132 271584
rect 161296 271532 161348 271584
rect 197636 271532 197688 271584
rect 214932 271532 214984 271584
rect 276020 271532 276072 271584
rect 372160 271532 372212 271584
rect 447140 271532 447192 271584
rect 52920 271464 52972 271516
rect 117320 271464 117372 271516
rect 164148 271464 164200 271516
rect 197728 271464 197780 271516
rect 205088 271464 205140 271516
rect 264980 271464 265032 271516
rect 363972 271464 364024 271516
rect 437480 271464 437532 271516
rect 48136 271396 48188 271448
rect 51908 271396 51960 271448
rect 53104 271396 53156 271448
rect 115940 271396 115992 271448
rect 210792 271396 210844 271448
rect 270500 271396 270552 271448
rect 361028 271396 361080 271448
rect 433340 271396 433392 271448
rect 48044 271328 48096 271380
rect 52460 271328 52512 271380
rect 53012 271328 53064 271380
rect 113548 271328 113600 271380
rect 219072 271328 219124 271380
rect 277676 271328 277728 271380
rect 368020 271328 368072 271380
rect 440240 271328 440292 271380
rect 503628 271328 503680 271380
rect 517612 271328 517664 271380
rect 51816 271260 51868 271312
rect 104900 271260 104952 271312
rect 183468 271260 183520 271312
rect 197360 271260 197412 271312
rect 209228 271260 209280 271312
rect 263600 271260 263652 271312
rect 362592 271260 362644 271312
rect 434720 271260 434772 271312
rect 51724 271192 51776 271244
rect 103520 271192 103572 271244
rect 206560 271192 206612 271244
rect 260840 271192 260892 271244
rect 343548 271192 343600 271244
rect 356980 271192 357032 271244
rect 370872 271192 370924 271244
rect 443000 271192 443052 271244
rect 503628 271192 503680 271244
rect 517704 271192 517756 271244
rect 50252 271124 50304 271176
rect 100760 271124 100812 271176
rect 183468 271124 183520 271176
rect 201592 271124 201644 271176
rect 202420 271124 202472 271176
rect 252560 271124 252612 271176
rect 277124 271124 277176 271176
rect 356612 271124 356664 271176
rect 356888 271124 356940 271176
rect 374920 271124 374972 271176
rect 413100 271124 413152 271176
rect 440148 271124 440200 271176
rect 516600 271124 516652 271176
rect 54668 271056 54720 271108
rect 88340 271056 88392 271108
rect 212172 271056 212224 271108
rect 258264 271056 258316 271108
rect 379060 271056 379112 271108
rect 416044 271056 416096 271108
rect 46112 270988 46164 271040
rect 77300 270988 77352 271040
rect 210700 270988 210752 271040
rect 255320 270988 255372 271040
rect 374828 270988 374880 271040
rect 409880 270988 409932 271040
rect 47768 270920 47820 270972
rect 78680 270920 78732 270972
rect 216128 270920 216180 270972
rect 247040 270920 247092 270972
rect 379152 270920 379204 270972
rect 407120 270920 407172 270972
rect 50344 270444 50396 270496
rect 51816 270444 51868 270496
rect 59820 270444 59872 270496
rect 107660 270444 107712 270496
rect 115848 270444 115900 270496
rect 196992 270444 197044 270496
rect 211712 270444 211764 270496
rect 212172 270444 212224 270496
rect 215116 270444 215168 270496
rect 216404 270444 216456 270496
rect 219808 270444 219860 270496
rect 220636 270444 220688 270496
rect 247040 270444 247092 270496
rect 280068 270444 280120 270496
rect 356612 270444 356664 270496
rect 357072 270444 357124 270496
rect 369768 270444 369820 270496
rect 371700 270444 371752 270496
rect 377036 270444 377088 270496
rect 378048 270444 378100 270496
rect 411260 270444 411312 270496
rect 81440 270376 81492 270428
rect 109040 270376 109092 270428
rect 117228 270376 117280 270428
rect 197176 270376 197228 270428
rect 211620 270376 211672 270428
rect 213092 270376 213144 270428
rect 213644 270376 213696 270428
rect 215668 270376 215720 270428
rect 216680 270376 216732 270428
rect 217232 270376 217284 270428
rect 263600 270376 263652 270428
rect 369676 270376 369728 270428
rect 401692 270376 401744 270428
rect 63500 270308 63552 270360
rect 92480 270308 92532 270360
rect 219164 270308 219216 270360
rect 251180 270308 251232 270360
rect 376300 270308 376352 270360
rect 377128 270308 377180 270360
rect 411352 270308 411404 270360
rect 53932 270240 53984 270292
rect 84200 270240 84252 270292
rect 220728 270240 220780 270292
rect 249800 270240 249852 270292
rect 375104 270240 375156 270292
rect 377496 270240 377548 270292
rect 378600 270240 378652 270292
rect 379796 270240 379848 270292
rect 379888 270240 379940 270292
rect 408500 270240 408552 270292
rect 53840 270172 53892 270224
rect 85580 270172 85632 270224
rect 219348 270172 219400 270224
rect 248512 270172 248564 270224
rect 370964 270172 371016 270224
rect 373632 270172 373684 270224
rect 400220 270172 400272 270224
rect 80060 270104 80112 270156
rect 111800 270104 111852 270156
rect 216772 270104 216824 270156
rect 219624 270104 219676 270156
rect 220728 270104 220780 270156
rect 224224 270104 224276 270156
rect 245660 270104 245712 270156
rect 375656 270104 375708 270156
rect 379704 270104 379756 270156
rect 405740 270104 405792 270156
rect 51816 270036 51868 270088
rect 84660 270036 84712 270088
rect 217048 270036 217100 270088
rect 219072 270036 219124 270088
rect 251272 270036 251324 270088
rect 371700 270036 371752 270088
rect 397460 270036 397512 270088
rect 55956 269968 56008 270020
rect 88340 269968 88392 270020
rect 219256 269968 219308 270020
rect 252560 269968 252612 270020
rect 372528 269968 372580 270020
rect 373908 269968 373960 270020
rect 398840 269968 398892 270020
rect 57980 269900 58032 269952
rect 91100 269900 91152 269952
rect 215668 269900 215720 269952
rect 224132 269900 224184 269952
rect 224408 269900 224460 269952
rect 265164 269900 265216 269952
rect 377496 269900 377548 269952
rect 407120 269900 407172 269952
rect 57060 269832 57112 269884
rect 89720 269832 89772 269884
rect 213092 269832 213144 269884
rect 224224 269832 224276 269884
rect 224316 269832 224368 269884
rect 262220 269832 262272 269884
rect 374368 269832 374420 269884
rect 379888 269832 379940 269884
rect 389272 269832 389324 269884
rect 420920 269832 420972 269884
rect 46664 269764 46716 269816
rect 59820 269764 59872 269816
rect 77852 269764 77904 269816
rect 113180 269764 113232 269816
rect 217876 269764 217928 269816
rect 218612 269764 218664 269816
rect 266360 269764 266412 269816
rect 371792 269764 371844 269816
rect 379152 269764 379204 269816
rect 379612 269764 379664 269816
rect 412916 269764 412968 269816
rect 209412 269696 209464 269748
rect 210792 269696 210844 269748
rect 239128 269696 239180 269748
rect 373724 269696 373776 269748
rect 376208 269696 376260 269748
rect 396080 269696 396132 269748
rect 224132 269628 224184 269680
rect 244280 269628 244332 269680
rect 377128 269628 377180 269680
rect 391940 269628 391992 269680
rect 212172 269560 212224 269612
rect 271880 269560 271932 269612
rect 216404 269492 216456 269544
rect 224316 269492 224368 269544
rect 217968 269424 218020 269476
rect 220636 269424 220688 269476
rect 219256 269288 219308 269340
rect 219808 269288 219860 269340
rect 54760 269220 54812 269272
rect 55956 269220 56008 269272
rect 218520 269220 218572 269272
rect 219624 269220 219676 269272
rect 224408 269220 224460 269272
rect 379152 269152 379204 269204
rect 389180 269152 389232 269204
rect 376484 269084 376536 269136
rect 390560 269084 390612 269136
rect 47952 269016 48004 269068
rect 53840 269016 53892 269068
rect 54576 269016 54628 269068
rect 214472 269016 214524 269068
rect 216036 269016 216088 269068
rect 219716 269016 219768 269068
rect 253940 269016 253992 269068
rect 376576 269016 376628 269068
rect 379060 269016 379112 269068
rect 383568 269016 383620 269068
rect 436192 269016 436244 269068
rect 45376 268948 45428 269000
rect 144920 268948 144972 269000
rect 213552 268948 213604 269000
rect 242900 268948 242952 269000
rect 372252 268948 372304 269000
rect 373816 268948 373868 269000
rect 433340 268948 433392 269000
rect 42248 268880 42300 268932
rect 107752 268880 107804 268932
rect 213276 268880 213328 268932
rect 215852 268880 215904 268932
rect 231860 268880 231912 268932
rect 259460 268880 259512 268932
rect 375932 268880 375984 268932
rect 376760 268880 376812 268932
rect 383384 268880 383436 268932
rect 383476 268880 383528 268932
rect 416780 268880 416832 268932
rect 49148 268812 49200 268864
rect 110420 268812 110472 268864
rect 216496 268812 216548 268864
rect 230480 268812 230532 268864
rect 259552 268812 259604 268864
rect 379980 268812 380032 268864
rect 414020 268812 414072 268864
rect 43904 268744 43956 268796
rect 57980 268744 58032 268796
rect 229192 268744 229244 268796
rect 260840 268744 260892 268796
rect 379244 268744 379296 268796
rect 409880 268744 409932 268796
rect 43812 268676 43864 268728
rect 57060 268676 57112 268728
rect 215852 268676 215904 268728
rect 255320 268676 255372 268728
rect 389180 268676 389232 268728
rect 419540 268676 419592 268728
rect 46848 268608 46900 268660
rect 53932 268608 53984 268660
rect 54484 268608 54536 268660
rect 207940 268608 207992 268660
rect 218520 268608 218572 268660
rect 258080 268608 258132 268660
rect 374920 268608 374972 268660
rect 375748 268608 375800 268660
rect 383476 268608 383528 268660
rect 390560 268608 390612 268660
rect 418252 268608 418304 268660
rect 50436 268540 50488 268592
rect 63500 268540 63552 268592
rect 216036 268540 216088 268592
rect 256700 268540 256752 268592
rect 377312 268540 377364 268592
rect 403532 268540 403584 268592
rect 43720 268472 43772 268524
rect 46480 268472 46532 268524
rect 80060 268472 80112 268524
rect 209504 268472 209556 268524
rect 213460 268472 213512 268524
rect 269120 268472 269172 268524
rect 391940 268472 391992 268524
rect 418160 268472 418212 268524
rect 43628 268404 43680 268456
rect 47860 268404 47912 268456
rect 81440 268404 81492 268456
rect 209596 268404 209648 268456
rect 213368 268404 213420 268456
rect 270500 268404 270552 268456
rect 45468 268336 45520 268388
rect 50436 268336 50488 268388
rect 53104 268336 53156 268388
rect 106372 268336 106424 268388
rect 206836 268336 206888 268388
rect 212080 268336 212132 268388
rect 273168 268336 273220 268388
rect 379060 268336 379112 268388
rect 404360 268336 404412 268388
rect 44916 268268 44968 268320
rect 147680 268268 147732 268320
rect 216312 268268 216364 268320
rect 231860 268268 231912 268320
rect 215116 268200 215168 268252
rect 218336 268200 218388 268252
rect 244372 268200 244424 268252
rect 375564 268200 375616 268252
rect 377312 268200 377364 268252
rect 191748 253852 191800 253904
rect 201408 253852 201460 253904
rect 202880 253852 202932 253904
rect 340788 253852 340840 253904
rect 357164 253920 357216 253972
rect 357532 253920 357584 253972
rect 500868 253308 500920 253360
rect 517796 253308 517848 253360
rect 180524 253240 180576 253292
rect 197636 253240 197688 253292
rect 198096 253240 198148 253292
rect 339408 253240 339460 253292
rect 360200 253240 360252 253292
rect 499212 253240 499264 253292
rect 517704 253240 517756 253292
rect 517980 253240 518032 253292
rect 179328 253172 179380 253224
rect 197544 253172 197596 253224
rect 351828 253172 351880 253224
rect 358084 253172 358136 253224
rect 517796 253172 517848 253224
rect 518072 253172 518124 253224
rect 510896 252560 510948 252612
rect 517520 252560 517572 252612
rect 58716 252492 58768 252544
rect 60832 252492 60884 252544
rect 374828 252492 374880 252544
rect 375288 252492 375340 252544
rect 436100 252492 436152 252544
rect 373632 252424 373684 252476
rect 375840 252424 375892 252476
rect 434720 252424 434772 252476
rect 372160 252356 372212 252408
rect 372436 252356 372488 252408
rect 429200 252356 429252 252408
rect 55864 252152 55916 252204
rect 60740 252152 60792 252204
rect 75828 252016 75880 252068
rect 98644 252016 98696 252068
rect 377128 252016 377180 252068
rect 389180 252016 389232 252068
rect 52920 251948 52972 252000
rect 83464 251948 83516 252000
rect 371056 251948 371108 252000
rect 379704 251948 379756 252000
rect 425704 251948 425756 252000
rect 58624 251880 58676 251932
rect 106280 251880 106332 251932
rect 214472 251880 214524 251932
rect 229100 251880 229152 251932
rect 370412 251880 370464 251932
rect 373540 251880 373592 251932
rect 421564 251880 421616 251932
rect 57612 251812 57664 251864
rect 104900 251812 104952 251864
rect 214840 251812 214892 251864
rect 230480 251812 230532 251864
rect 369584 251812 369636 251864
rect 372436 251812 372488 251864
rect 427084 251812 427136 251864
rect 50528 251132 50580 251184
rect 75828 251132 75880 251184
rect 43996 251064 44048 251116
rect 56876 251064 56928 251116
rect 57612 251064 57664 251116
rect 42616 250996 42668 251048
rect 52920 250996 52972 251048
rect 519452 183540 519504 183592
rect 520188 183540 520240 183592
rect 580264 183540 580316 183592
rect 520096 183472 520148 183524
rect 580356 183472 580408 183524
rect 204996 177964 205048 178016
rect 217048 177964 217100 178016
rect 363880 177964 363932 178016
rect 377036 177964 377088 178016
rect 216772 176808 216824 176860
rect 217048 176808 217100 176860
rect 202880 176604 202932 176656
rect 216680 176604 216732 176656
rect 202144 176128 202196 176180
rect 202880 176128 202932 176180
rect 358084 175924 358136 175976
rect 376944 175924 376996 175976
rect 207664 175176 207716 175228
rect 217140 175176 217192 175228
rect 365260 175176 365312 175228
rect 377404 175176 377456 175228
rect 216772 175108 216824 175160
rect 217048 175108 217100 175160
rect 52000 166948 52052 167000
rect 101036 166948 101088 167000
rect 197452 166948 197504 167000
rect 201500 166948 201552 167000
rect 362500 166948 362552 167000
rect 423404 166948 423456 167000
rect 50896 166880 50948 166932
rect 103520 166880 103572 166932
rect 358268 166880 358320 166932
rect 418436 166880 418488 166932
rect 50804 166812 50856 166864
rect 108304 166812 108356 166864
rect 214748 166812 214800 166864
rect 260932 166812 260984 166864
rect 358360 166812 358412 166864
rect 421012 166812 421064 166864
rect 58992 166744 59044 166796
rect 140872 166744 140924 166796
rect 203524 166744 203576 166796
rect 265900 166744 265952 166796
rect 356796 166744 356848 166796
rect 445852 166744 445904 166796
rect 56232 166676 56284 166728
rect 138480 166676 138532 166728
rect 203708 166676 203760 166728
rect 270868 166676 270920 166728
rect 369308 166676 369360 166728
rect 470968 166676 471020 166728
rect 60004 166608 60056 166660
rect 145932 166608 145984 166660
rect 204904 166608 204956 166660
rect 285956 166608 286008 166660
rect 373448 166608 373500 166660
rect 475844 166608 475896 166660
rect 59176 166540 59228 166592
rect 148508 166540 148560 166592
rect 210608 166540 210660 166592
rect 295892 166540 295944 166592
rect 370780 166540 370832 166592
rect 473452 166540 473504 166592
rect 59912 166472 59964 166524
rect 150900 166472 150952 166524
rect 206468 166472 206520 166524
rect 293408 166472 293460 166524
rect 372068 166472 372120 166524
rect 480904 166472 480956 166524
rect 58900 166404 58952 166456
rect 153292 166404 153344 166456
rect 203616 166404 203668 166456
rect 291016 166404 291068 166456
rect 367928 166404 367980 166456
rect 478420 166404 478472 166456
rect 41052 166336 41104 166388
rect 163320 166336 163372 166388
rect 209136 166336 209188 166388
rect 298468 166336 298520 166388
rect 365168 166336 365220 166388
rect 483388 166336 483440 166388
rect 41144 166268 41196 166320
rect 165896 166268 165948 166320
rect 202328 166268 202380 166320
rect 305920 166268 305972 166320
rect 366640 166268 366692 166320
rect 485964 166268 486016 166320
rect 49516 166200 49568 166252
rect 98460 166200 98512 166252
rect 374644 166200 374696 166252
rect 430948 166200 431000 166252
rect 50712 166132 50764 166184
rect 96068 166132 96120 166184
rect 373356 166132 373408 166184
rect 428188 166132 428240 166184
rect 357624 165588 357676 165640
rect 360292 165588 360344 165640
rect 373632 165588 373684 165640
rect 373816 165588 373868 165640
rect 433340 165588 433392 165640
rect 50528 165520 50580 165572
rect 51632 165520 51684 165572
rect 54208 165520 54260 165572
rect 132500 165520 132552 165572
rect 209044 165520 209096 165572
rect 325884 165520 325936 165572
rect 343272 165520 343324 165572
rect 356980 165520 357032 165572
rect 357440 165520 357492 165572
rect 362408 165520 362460 165572
rect 458364 165520 458416 165572
rect 55036 165452 55088 165504
rect 128360 165452 128412 165504
rect 214656 165452 214708 165504
rect 308404 165452 308456 165504
rect 360936 165452 360988 165504
rect 447324 165452 447376 165504
rect 56508 165384 56560 165436
rect 129740 165384 129792 165436
rect 214564 165384 214616 165436
rect 300860 165384 300912 165436
rect 371976 165384 372028 165436
rect 455420 165384 455472 165436
rect 53288 165316 53340 165368
rect 123484 165316 123536 165368
rect 211896 165316 211948 165368
rect 280160 165316 280212 165368
rect 370688 165316 370740 165368
rect 452660 165316 452712 165368
rect 56324 165248 56376 165300
rect 125876 165248 125928 165300
rect 218980 165248 219032 165300
rect 283380 165248 283432 165300
rect 369124 165248 369176 165300
rect 449900 165248 449952 165300
rect 54944 165180 54996 165232
rect 120908 165180 120960 165232
rect 183284 165180 183336 165232
rect 197360 165180 197412 165232
rect 206376 165180 206428 165232
rect 267924 165180 267976 165232
rect 366456 165180 366508 165232
rect 443000 165180 443052 165232
rect 53196 165112 53248 165164
rect 115940 165112 115992 165164
rect 218796 165112 218848 165164
rect 277400 165112 277452 165164
rect 365076 165112 365128 165164
rect 438032 165112 438084 165164
rect 503260 165112 503312 165164
rect 517612 165112 517664 165164
rect 56048 165044 56100 165096
rect 118332 165044 118384 165096
rect 183376 165044 183428 165096
rect 197452 165044 197504 165096
rect 215944 165044 215996 165096
rect 258080 165044 258132 165096
rect 369216 165044 369268 165096
rect 434720 165044 434772 165096
rect 440240 165044 440292 165096
rect 516600 165044 516652 165096
rect 54852 164976 54904 165028
rect 113548 164976 113600 165028
rect 117320 164976 117372 165028
rect 196808 164976 196860 165028
rect 210516 164976 210568 165028
rect 252560 164976 252612 165028
rect 367836 164976 367888 165028
rect 433340 164976 433392 165028
rect 503352 164976 503404 165028
rect 517888 164976 517940 165028
rect 52184 164908 52236 164960
rect 105728 164908 105780 164960
rect 115940 164908 115992 164960
rect 196716 164908 196768 164960
rect 210424 164908 210476 164960
rect 249800 164908 249852 164960
rect 374736 164908 374788 164960
rect 49608 164840 49660 164892
rect 92480 164840 92532 164892
rect 114560 164840 114612 164892
rect 196624 164840 196676 164892
rect 218888 164840 218940 164892
rect 247684 164840 247736 164892
rect 343456 164840 343508 164892
rect 357624 164840 357676 164892
rect 373264 164840 373316 164892
rect 416044 164840 416096 164892
rect 52092 164772 52144 164824
rect 90272 164772 90324 164824
rect 376116 164772 376168 164824
rect 409880 164772 409932 164824
rect 510528 164908 510580 164960
rect 517520 164908 517572 164960
rect 440332 164772 440384 164824
rect 56416 164704 56468 164756
rect 88340 164704 88392 164756
rect 378876 164704 378928 164756
rect 412640 164704 412692 164756
rect 378968 164636 379020 164688
rect 407120 164636 407172 164688
rect 428924 164568 428976 164620
rect 433524 164568 433576 164620
rect 51632 164228 51684 164280
rect 73804 164228 73856 164280
rect 87604 164228 87656 164280
rect 108304 164228 108356 164280
rect 46572 164160 46624 164212
rect 53288 164160 53340 164212
rect 58624 164160 58676 164212
rect 60004 164160 60056 164212
rect 60096 164160 60148 164212
rect 117872 164160 117924 164212
rect 211988 164160 212040 164212
rect 323032 164160 323084 164212
rect 377404 164160 377456 164212
rect 437756 164160 437808 164212
rect 46480 164092 46532 164144
rect 52184 164092 52236 164144
rect 53380 164092 53432 164144
rect 110972 164092 111024 164144
rect 219624 164092 219676 164144
rect 264980 164092 265032 164144
rect 374552 164092 374604 164144
rect 434720 164092 434772 164144
rect 55864 164024 55916 164076
rect 57520 164024 57572 164076
rect 57704 164024 57756 164076
rect 105176 164024 105228 164076
rect 216588 164024 216640 164076
rect 236092 164024 236144 164076
rect 375012 164024 375064 164076
rect 396172 164024 396224 164076
rect 54392 163956 54444 164008
rect 55036 163956 55088 164008
rect 100852 163956 100904 164008
rect 216220 163956 216272 164008
rect 236000 163956 236052 164008
rect 376208 163956 376260 164008
rect 396080 163956 396132 164008
rect 52828 163888 52880 163940
rect 56508 163888 56560 163940
rect 96620 163888 96672 163940
rect 52920 163820 52972 163872
rect 55128 163820 55180 163872
rect 98000 163820 98052 163872
rect 60004 163752 60056 163804
rect 106372 163752 106424 163804
rect 47860 163684 47912 163736
rect 53380 163684 53432 163736
rect 109684 163684 109736 163736
rect 59360 163616 59412 163668
rect 119068 163616 119120 163668
rect 375196 163616 375248 163668
rect 422300 163616 422352 163668
rect 52184 163548 52236 163600
rect 111892 163548 111944 163600
rect 372160 163548 372212 163600
rect 375012 163548 375064 163600
rect 429292 163548 429344 163600
rect 53288 163480 53340 163532
rect 113180 163480 113232 163532
rect 216680 163480 216732 163532
rect 218888 163480 218940 163532
rect 263784 163480 263836 163532
rect 373172 163480 373224 163532
rect 375104 163480 375156 163532
rect 431960 163480 432012 163532
rect 52368 163412 52420 163464
rect 57244 163412 57296 163464
rect 95240 163412 95292 163464
rect 57520 163344 57572 163396
rect 60096 163344 60148 163396
rect 375196 162868 375248 162920
rect 49148 162800 49200 162852
rect 53472 162800 53524 162852
rect 57060 162800 57112 162852
rect 59176 162800 59228 162852
rect 216036 162800 216088 162852
rect 217140 162800 217192 162852
rect 214472 162664 214524 162716
rect 260840 162800 260892 162852
rect 214840 162596 214892 162648
rect 259552 162732 259604 162784
rect 217876 162664 217928 162716
rect 259460 162664 259512 162716
rect 376300 162800 376352 162852
rect 379796 162800 379848 162852
rect 379980 162800 380032 162852
rect 436100 162800 436152 162852
rect 377220 162732 377272 162784
rect 420920 162732 420972 162784
rect 376300 162664 376352 162716
rect 418620 162664 418672 162716
rect 218520 162596 218572 162648
rect 218980 162596 219032 162648
rect 258080 162596 258132 162648
rect 376208 162596 376260 162648
rect 376392 162596 376444 162648
rect 379152 162596 379204 162648
rect 419540 162596 419592 162648
rect 375932 162528 375984 162580
rect 379980 162528 380032 162580
rect 374920 162460 374972 162512
rect 379152 162460 379204 162512
rect 379796 162256 379848 162308
rect 418160 162256 418212 162308
rect 59176 162188 59228 162240
rect 89904 162188 89956 162240
rect 372252 162188 372304 162240
rect 373724 162188 373776 162240
rect 428924 162188 428976 162240
rect 53472 162120 53524 162172
rect 111156 162120 111208 162172
rect 218612 162120 218664 162172
rect 219532 162120 219584 162172
rect 266360 162120 266412 162172
rect 372344 162120 372396 162172
rect 374828 162120 374880 162172
rect 430580 162120 430632 162172
rect 376576 161916 376628 161968
rect 377220 161916 377272 161968
rect 216220 161508 216272 161560
rect 235264 161508 235316 161560
rect 217140 161440 217192 161492
rect 236644 161440 236696 161492
rect 379152 161440 379204 161492
rect 396724 161440 396776 161492
rect 357532 156612 357584 156664
rect 357716 156612 357768 156664
rect 215760 148996 215812 149048
rect 216496 148996 216548 149048
rect 278780 148996 278832 149048
rect 379704 148996 379756 149048
rect 427912 148996 427964 149048
rect 215024 148928 215076 148980
rect 276112 148928 276164 148980
rect 214932 148860 214984 148912
rect 240140 148860 240192 148912
rect 46664 148656 46716 148708
rect 59912 148656 59964 148708
rect 87604 148656 87656 148708
rect 213184 148656 213236 148708
rect 238760 148656 238812 148708
rect 46756 148588 46808 148640
rect 52000 148588 52052 148640
rect 80060 148588 80112 148640
rect 212264 148588 212316 148640
rect 214564 148588 214616 148640
rect 241520 148588 241572 148640
rect 373908 148588 373960 148640
rect 376024 148588 376076 148640
rect 398840 148588 398892 148640
rect 49240 148520 49292 148572
rect 53196 148520 53248 148572
rect 81440 148520 81492 148572
rect 213368 148520 213420 148572
rect 214656 148520 214708 148572
rect 270500 148520 270552 148572
rect 371700 148520 371752 148572
rect 374644 148520 374696 148572
rect 397460 148520 397512 148572
rect 56232 148452 56284 148504
rect 114560 148452 114612 148504
rect 215852 148452 215904 148504
rect 271880 148452 271932 148504
rect 370964 148452 371016 148504
rect 371976 148452 372028 148504
rect 400220 148452 400272 148504
rect 56324 148384 56376 148436
rect 117320 148384 117372 148436
rect 212908 148384 212960 148436
rect 214840 148384 214892 148436
rect 274640 148384 274692 148436
rect 372712 148384 372764 148436
rect 401600 148384 401652 148436
rect 53012 148316 53064 148368
rect 115940 148316 115992 148368
rect 212080 148316 212132 148368
rect 213736 148316 213788 148368
rect 274732 148316 274784 148368
rect 372436 148316 372488 148368
rect 379980 148316 380032 148368
rect 429200 148316 429252 148368
rect 213000 147704 213052 147756
rect 215024 147704 215076 147756
rect 213644 147636 213696 147688
rect 214932 147636 214984 147688
rect 379428 147636 379480 147688
rect 379704 147636 379756 147688
rect 212172 147568 212224 147620
rect 215852 147568 215904 147620
rect 369676 147568 369728 147620
rect 372712 147568 372764 147620
rect 373264 147568 373316 147620
rect 210792 147500 210844 147552
rect 213184 147500 213236 147552
rect 47768 146208 47820 146260
rect 51724 146208 51776 146260
rect 54760 146208 54812 146260
rect 59728 146208 59780 146260
rect 99380 146208 99432 146260
rect 179052 146208 179104 146260
rect 197544 146208 197596 146260
rect 235264 146208 235316 146260
rect 255320 146208 255372 146260
rect 276020 146208 276072 146260
rect 356888 146208 356940 146260
rect 374736 146208 374788 146260
rect 375564 146208 375616 146260
rect 376484 146208 376536 146260
rect 377496 146208 377548 146260
rect 57060 146140 57112 146192
rect 57980 146140 58032 146192
rect 179696 146140 179748 146192
rect 197636 146140 197688 146192
rect 219256 146140 219308 146192
rect 52920 146072 52972 146124
rect 53840 146072 53892 146124
rect 86960 146072 87012 146124
rect 236644 146140 236696 146192
rect 256700 146140 256752 146192
rect 338488 146140 338540 146192
rect 360200 146140 360252 146192
rect 374460 146140 374512 146192
rect 375196 146140 375248 146192
rect 375932 146140 375984 146192
rect 378968 146140 379020 146192
rect 379336 146208 379388 146260
rect 379612 146208 379664 146260
rect 404360 146208 404412 146260
rect 251180 146072 251232 146124
rect 340236 146072 340288 146124
rect 357716 146072 357768 146124
rect 396724 146140 396776 146192
rect 416780 146140 416832 146192
rect 500224 146140 500276 146192
rect 517520 146140 517572 146192
rect 517796 146140 517848 146192
rect 412732 146072 412784 146124
rect 498660 146072 498712 146124
rect 517704 146072 517756 146124
rect 57980 146004 58032 146056
rect 91100 146004 91152 146056
rect 219072 146004 219124 146056
rect 251272 146004 251324 146056
rect 378600 146004 378652 146056
rect 411260 146004 411312 146056
rect 56140 145936 56192 145988
rect 88432 145936 88484 145988
rect 217876 145936 217928 145988
rect 249800 145936 249852 145988
rect 377864 145936 377916 145988
rect 379244 145936 379296 145988
rect 409972 145936 410024 145988
rect 54944 145868 54996 145920
rect 85580 145868 85632 145920
rect 219348 145868 219400 145920
rect 248420 145868 248472 145920
rect 377496 145868 377548 145920
rect 407212 145868 407264 145920
rect 46388 145800 46440 145852
rect 52368 145800 52420 145852
rect 77300 145800 77352 145852
rect 215116 145800 215168 145852
rect 244280 145800 244332 145852
rect 375656 145800 375708 145852
rect 405740 145800 405792 145852
rect 51724 145732 51776 145784
rect 78680 145732 78732 145784
rect 217968 145732 218020 145784
rect 247040 145732 247092 145784
rect 375196 145732 375248 145784
rect 403072 145732 403124 145784
rect 49332 145664 49384 145716
rect 54576 145664 54628 145716
rect 82820 145664 82872 145716
rect 216128 145664 216180 145716
rect 219348 145664 219400 145716
rect 219440 145664 219492 145716
rect 244372 145664 244424 145716
rect 375564 145664 375616 145716
rect 402980 145664 403032 145716
rect 56416 145596 56468 145648
rect 84200 145596 84252 145648
rect 215668 145596 215720 145648
rect 216312 145596 216364 145648
rect 216588 145596 216640 145648
rect 242900 145596 242952 145648
rect 378784 145596 378836 145648
rect 408500 145596 408552 145648
rect 517520 145596 517572 145648
rect 580264 145596 580316 145648
rect 58624 145528 58676 145580
rect 91192 145528 91244 145580
rect 191288 145528 191340 145580
rect 202144 145528 202196 145580
rect 204904 145528 204956 145580
rect 217048 145528 217100 145580
rect 219072 145528 219124 145580
rect 219348 145528 219400 145580
rect 245660 145528 245712 145580
rect 280068 145528 280120 145580
rect 307668 145528 307720 145580
rect 351644 145528 351696 145580
rect 358084 145528 358136 145580
rect 358728 145528 358780 145580
rect 510528 145528 510580 145580
rect 517704 145528 517756 145580
rect 580356 145528 580408 145580
rect 58808 145460 58860 145512
rect 84292 145460 84344 145512
rect 218520 145460 218572 145512
rect 236092 145460 236144 145512
rect 378968 145460 379020 145512
rect 396172 145460 396224 145512
rect 47676 145392 47728 145444
rect 54668 145392 54720 145444
rect 76012 145392 76064 145444
rect 219072 145392 219124 145444
rect 236000 145392 236052 145444
rect 378876 145392 378928 145444
rect 396080 145392 396132 145444
rect 47492 145324 47544 145376
rect 54852 145324 54904 145376
rect 75920 145324 75972 145376
rect 216312 145324 216364 145376
rect 219440 145324 219492 145376
rect 219716 145324 219768 145376
rect 253940 145324 253992 145376
rect 379888 145324 379940 145376
rect 414020 145324 414072 145376
rect 59636 145256 59688 145308
rect 93860 145256 93912 145308
rect 219808 145256 219860 145308
rect 252560 145256 252612 145308
rect 378048 145256 378100 145308
rect 411352 145256 411404 145308
rect 216772 145120 216824 145172
rect 217876 145120 217928 145172
rect 218612 145052 218664 145104
rect 219256 145052 219308 145104
rect 216404 144916 216456 144968
rect 217968 144916 218020 144968
rect 219256 144916 219308 144968
rect 219808 144916 219860 144968
rect 54484 144848 54536 144900
rect 55864 144848 55916 144900
rect 56416 144848 56468 144900
rect 209320 144848 209372 144900
rect 213276 144848 213328 144900
rect 213552 144848 213604 144900
rect 216036 144848 216088 144900
rect 216588 144848 216640 144900
rect 307668 144848 307720 144900
rect 356612 144848 356664 144900
rect 374368 144848 374420 144900
rect 378784 144848 378836 144900
rect 51816 144780 51868 144832
rect 58808 144780 58860 144832
rect 213460 144780 213512 144832
rect 214932 144780 214984 144832
rect 51908 144712 51960 144764
rect 58624 144712 58676 144764
rect 213092 144712 213144 144764
rect 218796 144712 218848 144764
rect 219348 144712 219400 144764
rect 53104 144644 53156 144696
rect 58900 144644 58952 144696
rect 50436 144576 50488 144628
rect 58716 144576 58768 144628
rect 219900 143284 219952 143336
rect 220084 143284 220136 143336
rect 3240 97928 3292 97980
rect 21364 97928 21416 97980
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 202236 70320 202288 70372
rect 216680 70320 216732 70372
rect 363788 70320 363840 70372
rect 376944 70320 376996 70372
rect 358084 68416 358136 68468
rect 358728 68416 358780 68468
rect 376944 68280 376996 68332
rect 204904 67600 204956 67652
rect 216680 67600 216732 67652
rect 218336 61072 218388 61124
rect 218612 61072 218664 61124
rect 378968 59712 379020 59764
rect 396080 59712 396132 59764
rect 54668 59644 54720 59696
rect 77116 59644 77168 59696
rect 218520 59644 218572 59696
rect 237104 59644 237156 59696
rect 378876 59644 378928 59696
rect 397092 59644 397144 59696
rect 55036 59576 55088 59628
rect 100760 59576 100812 59628
rect 216220 59576 216272 59628
rect 255872 59576 255924 59628
rect 379152 59576 379204 59628
rect 416964 59576 417016 59628
rect 54576 59508 54628 59560
rect 83096 59508 83148 59560
rect 217140 59508 217192 59560
rect 256976 59508 257028 59560
rect 376208 59508 376260 59560
rect 422852 59508 422904 59560
rect 54760 59440 54812 59492
rect 99472 59440 99524 59492
rect 218888 59440 218940 59492
rect 263876 59440 263928 59492
rect 377220 59440 377272 59492
rect 423956 59440 424008 59492
rect 48228 59372 48280 59424
rect 105912 59372 105964 59424
rect 215852 59372 215904 59424
rect 262864 59372 262916 59424
rect 358176 59372 358228 59424
rect 416044 59372 416096 59424
rect 55864 59304 55916 59356
rect 84200 59304 84252 59356
rect 217968 59304 218020 59356
rect 358084 59304 358136 59356
rect 375196 59304 375248 59356
rect 403072 59304 403124 59356
rect 59176 59236 59228 59288
rect 89996 59236 90048 59288
rect 218980 59236 219032 59288
rect 258080 59236 258132 59288
rect 379796 59236 379848 59288
rect 418160 59236 418212 59288
rect 59820 59168 59872 59220
rect 94504 59168 94556 59220
rect 214748 59168 214800 59220
rect 260656 59168 260708 59220
rect 374736 59168 374788 59220
rect 404176 59168 404228 59220
rect 57244 59100 57296 59152
rect 95884 59100 95936 59152
rect 214472 59100 214524 59152
rect 261760 59100 261812 59152
rect 279240 59100 279292 59152
rect 356612 59100 356664 59152
rect 376116 59100 376168 59152
rect 419356 59100 419408 59152
rect 56508 59032 56560 59084
rect 96988 59032 97040 59084
rect 212448 59032 212500 59084
rect 290924 59032 290976 59084
rect 376392 59032 376444 59084
rect 420644 59032 420696 59084
rect 56140 58964 56192 59016
rect 102784 58964 102836 59016
rect 201316 58964 201368 59016
rect 300860 58964 300912 59016
rect 376576 58964 376628 59016
rect 421748 58964 421800 59016
rect 58900 58896 58952 58948
rect 107568 58896 107620 58948
rect 212356 58896 212408 58948
rect 315856 58896 315908 58948
rect 362224 58896 362276 58948
rect 423496 58896 423548 58948
rect 51632 58828 51684 58880
rect 101772 58828 101824 58880
rect 202788 58828 202840 58880
rect 308496 58828 308548 58880
rect 356704 58828 356756 58880
rect 425980 58828 426032 58880
rect 53656 58760 53708 58812
rect 138388 58760 138440 58812
rect 206192 58760 206244 58812
rect 320916 58760 320968 58812
rect 366364 58760 366416 58812
rect 453396 58760 453448 58812
rect 50988 58692 51040 58744
rect 148508 58692 148560 58744
rect 198648 58692 198700 58744
rect 325884 58692 325936 58744
rect 364984 58692 365036 58744
rect 475844 58692 475896 58744
rect 53564 58624 53616 58676
rect 150900 58624 150952 58676
rect 219256 58624 219308 58676
rect 428188 58624 428240 58676
rect 57244 57876 57296 57928
rect 57888 57876 57940 57928
rect 204904 57876 204956 57928
rect 210976 57876 211028 57928
rect 323308 57876 323360 57928
rect 343456 57876 343508 57928
rect 357624 57876 357676 57928
rect 358636 57876 358688 57928
rect 478420 57876 478472 57928
rect 503260 57876 503312 57928
rect 517612 57876 517664 57928
rect 52276 57808 52328 57860
rect 145564 57808 145616 57860
rect 183468 57808 183520 57860
rect 197452 57808 197504 57860
rect 209688 57808 209740 57860
rect 310980 57808 311032 57860
rect 343180 57808 343232 57860
rect 357440 57808 357492 57860
rect 376668 57808 376720 57860
rect 485964 57808 486016 57860
rect 503536 57808 503588 57860
rect 517888 57808 517940 57860
rect 41236 57740 41288 57792
rect 123484 57740 123536 57792
rect 183192 57740 183244 57792
rect 197360 57740 197412 57792
rect 215208 57740 215260 57792
rect 313372 57740 313424 57792
rect 363696 57740 363748 57792
rect 465908 57740 465960 57792
rect 53748 57672 53800 57724
rect 130844 57672 130896 57724
rect 218704 57672 218756 57724
rect 318340 57672 318392 57724
rect 360844 57672 360896 57724
rect 445852 57672 445904 57724
rect 53288 57604 53340 57656
rect 113180 57604 113232 57656
rect 205548 57604 205600 57656
rect 295892 57604 295944 57656
rect 363604 57604 363656 57656
rect 448244 57604 448296 57656
rect 59084 57536 59136 57588
rect 103796 57536 103848 57588
rect 213828 57536 213880 57588
rect 303436 57536 303488 57588
rect 362316 57536 362368 57588
rect 443460 57536 443512 57588
rect 55128 57468 55180 57520
rect 98092 57468 98144 57520
rect 215576 57468 215628 57520
rect 305828 57468 305880 57520
rect 367744 57468 367796 57520
rect 435916 57468 435968 57520
rect 51540 57400 51592 57452
rect 88340 57400 88392 57452
rect 211068 57400 211120 57452
rect 293316 57400 293368 57452
rect 371884 57400 371936 57452
rect 438492 57400 438544 57452
rect 59268 57332 59320 57384
rect 93676 57332 93728 57384
rect 218428 57332 218480 57384
rect 298100 57332 298152 57384
rect 370596 57332 370648 57384
rect 433524 57332 433576 57384
rect 52368 57264 52420 57316
rect 78220 57264 78272 57316
rect 211804 57264 211856 57316
rect 283472 57264 283524 57316
rect 370504 57264 370556 57316
rect 418436 57264 418488 57316
rect 54852 57196 54904 57248
rect 76012 57196 76064 57248
rect 218612 57196 218664 57248
rect 258356 57196 258408 57248
rect 379060 57196 379112 57248
rect 415492 57196 415544 57248
rect 77852 56584 77904 56636
rect 117872 56584 117924 56636
rect 41328 56516 41380 56568
rect 115940 56516 115992 56568
rect 214564 56516 214616 56568
rect 241612 56516 241664 56568
rect 374644 56516 374696 56568
rect 398196 56516 398248 56568
rect 52184 56448 52236 56500
rect 112076 56448 112128 56500
rect 219072 56448 219124 56500
rect 236000 56448 236052 56500
rect 374552 56448 374604 56500
rect 435732 56448 435784 56500
rect 56324 56380 56376 56432
rect 114100 56380 114152 56432
rect 215024 56380 215076 56432
rect 273260 56380 273312 56432
rect 373816 56380 373868 56432
rect 433340 56380 433392 56432
rect 53380 56312 53432 56364
rect 109500 56312 109552 56364
rect 214656 56312 214708 56364
rect 271052 56312 271104 56364
rect 374828 56312 374880 56364
rect 431132 56312 431184 56364
rect 59912 56244 59964 56296
rect 108580 56244 108632 56296
rect 219900 56244 219952 56296
rect 268476 56244 268528 56296
rect 379428 56244 379480 56296
rect 427636 56244 427688 56296
rect 58716 56176 58768 56228
rect 93308 56176 93360 56228
rect 219164 56176 219216 56228
rect 266360 56176 266412 56228
rect 379704 56176 379756 56228
rect 426440 56176 426492 56228
rect 56232 56108 56284 56160
rect 88708 56108 88760 56160
rect 219348 56108 219400 56160
rect 253388 56108 253440 56160
rect 379888 56108 379940 56160
rect 414572 56108 414624 56160
rect 54944 56040 54996 56092
rect 86500 56040 86552 56092
rect 218336 56040 218388 56092
rect 251180 56040 251232 56092
rect 379336 56040 379388 56092
rect 412640 56040 412692 56092
rect 52000 55972 52052 56024
rect 80428 55972 80480 56024
rect 216128 55972 216180 56024
rect 248604 55972 248656 56024
rect 378600 55972 378652 56024
rect 411260 55972 411312 56024
rect 58808 55904 58860 55956
rect 85396 55904 85448 55956
rect 216312 55904 216364 55956
rect 245292 55904 245344 55956
rect 378784 55904 378836 55956
rect 408684 55904 408736 55956
rect 213184 55836 213236 55888
rect 239128 55836 239180 55888
rect 371976 55836 372028 55888
rect 400404 55836 400456 55888
rect 219992 55768 220044 55820
rect 408316 55768 408368 55820
rect 213000 55700 213052 55752
rect 275100 55700 275152 55752
rect 53012 55156 53064 55208
rect 114560 55156 114612 55208
rect 216496 55156 216548 55208
rect 277400 55156 277452 55208
rect 375840 55156 375892 55208
rect 436100 55156 436152 55208
rect 56416 55088 56468 55140
rect 116124 55088 116176 55140
rect 213736 55088 213788 55140
rect 273352 55088 273404 55140
rect 376024 55088 376076 55140
rect 398840 55088 398892 55140
rect 53472 55020 53524 55072
rect 110420 55020 110472 55072
rect 215944 55020 215996 55072
rect 271880 55020 271932 55072
rect 375104 55020 375156 55072
rect 431960 55020 432012 55072
rect 42708 54952 42760 55004
rect 89720 54952 89772 55004
rect 219532 54952 219584 55004
rect 266452 54952 266504 55004
rect 375012 54952 375064 55004
rect 429200 54952 429252 55004
rect 60004 54884 60056 54936
rect 106280 54884 106332 54936
rect 219624 54884 219676 54936
rect 264980 54884 265032 54936
rect 379980 54884 380032 54936
rect 427820 54884 427872 54936
rect 57060 54816 57112 54868
rect 91100 54816 91152 54868
rect 219716 54816 219768 54868
rect 253940 54816 253992 54868
rect 378048 54816 378100 54868
rect 411352 54816 411404 54868
rect 52920 54748 52972 54800
rect 86960 54748 87012 54800
rect 217048 54748 217100 54800
rect 251364 54748 251416 54800
rect 377864 54748 377916 54800
rect 409880 54748 409932 54800
rect 58624 54680 58676 54732
rect 91468 54680 91520 54732
rect 217876 54680 217928 54732
rect 249800 54680 249852 54732
rect 376484 54680 376536 54732
rect 407212 54680 407264 54732
rect 53196 54612 53248 54664
rect 81440 54612 81492 54664
rect 216404 54612 216456 54664
rect 247040 54612 247092 54664
rect 375288 54612 375340 54664
rect 405832 54612 405884 54664
rect 51724 54544 51776 54596
rect 78680 54544 78732 54596
rect 215116 54544 215168 54596
rect 244372 54544 244424 54596
rect 375932 54544 375984 54596
rect 404360 54544 404412 54596
rect 218796 54476 218848 54528
rect 245660 54476 245712 54528
rect 373264 54476 373316 54528
rect 401600 54476 401652 54528
rect 216036 54408 216088 54460
rect 242900 54408 242952 54460
rect 373724 54408 373776 54460
rect 433432 54408 433484 54460
rect 213276 54340 213328 54392
rect 237380 54340 237432 54392
rect 213644 54272 213696 54324
rect 240140 54272 240192 54324
rect 572 3408 624 3460
rect 57244 3408 57296 3460
rect 125876 2796 125928 2848
rect 367100 2796 367152 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 636886 3464 684247
rect 18604 639056 18656 639062
rect 18604 638998 18656 639004
rect 3424 636880 3476 636886
rect 3424 636822 3476 636828
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 568546 3464 579935
rect 3424 568540 3476 568546
rect 3424 568482 3476 568488
rect 3422 547904 3478 547913
rect 3422 547839 3478 547848
rect 3436 514865 3464 547839
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 14464 486464 14516 486470
rect 14464 486406 14516 486412
rect 3424 483676 3476 483682
rect 3424 483618 3476 483624
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3436 19417 3464 483618
rect 3514 482216 3570 482225
rect 3514 482151 3570 482160
rect 3528 58585 3556 482151
rect 3608 480956 3660 480962
rect 3608 480898 3660 480904
rect 3620 462641 3648 480898
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 14476 411262 14504 486406
rect 14464 411256 14516 411262
rect 14464 411198 14516 411204
rect 18616 358766 18644 638998
rect 21364 560312 21416 560318
rect 21364 560254 21416 560260
rect 18604 358760 18656 358766
rect 18604 358702 18656 358708
rect 21376 97986 21404 560254
rect 40052 557530 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 59084 649324 59136 649330
rect 59084 649266 59136 649272
rect 56508 633684 56560 633690
rect 56508 633626 56560 633632
rect 54852 633616 54904 633622
rect 54852 633558 54904 633564
rect 54864 568070 54892 633558
rect 55128 633548 55180 633554
rect 55128 633490 55180 633496
rect 54944 630760 54996 630766
rect 54944 630702 54996 630708
rect 54852 568064 54904 568070
rect 54852 568006 54904 568012
rect 40040 557524 40092 557530
rect 40040 557466 40092 557472
rect 54956 549982 54984 630702
rect 55036 630692 55088 630698
rect 55036 630634 55088 630640
rect 55048 550390 55076 630634
rect 55140 550458 55168 633490
rect 56416 630828 56468 630834
rect 56416 630770 56468 630776
rect 55128 550452 55180 550458
rect 55128 550394 55180 550400
rect 55036 550384 55088 550390
rect 55036 550326 55088 550332
rect 56428 550050 56456 630770
rect 56520 550186 56548 633626
rect 57796 630964 57848 630970
rect 57796 630906 57848 630912
rect 57702 622432 57758 622441
rect 57702 622367 57758 622376
rect 57518 619712 57574 619721
rect 57518 619647 57574 619656
rect 57242 595232 57298 595241
rect 57242 595167 57298 595176
rect 57150 589112 57206 589121
rect 57150 589047 57206 589056
rect 57058 576872 57114 576881
rect 57058 576807 57114 576816
rect 57072 562426 57100 576807
rect 57164 568410 57192 589047
rect 57256 569158 57284 595167
rect 57426 591832 57482 591841
rect 57426 591767 57482 591776
rect 57334 579728 57390 579737
rect 57334 579663 57390 579672
rect 57244 569152 57296 569158
rect 57244 569094 57296 569100
rect 57152 568404 57204 568410
rect 57152 568346 57204 568352
rect 57060 562420 57112 562426
rect 57060 562362 57112 562368
rect 57348 552974 57376 579663
rect 57440 563922 57468 591767
rect 57532 566642 57560 619647
rect 57610 613592 57666 613601
rect 57610 613527 57666 613536
rect 57520 566636 57572 566642
rect 57520 566578 57572 566584
rect 57428 563916 57480 563922
rect 57428 563858 57480 563864
rect 57624 558346 57652 613527
rect 57612 558340 57664 558346
rect 57612 558282 57664 558288
rect 57336 552968 57388 552974
rect 57336 552910 57388 552916
rect 57716 551342 57744 622367
rect 57704 551336 57756 551342
rect 57704 551278 57756 551284
rect 57808 550322 57836 630906
rect 58990 628688 59046 628697
rect 58990 628623 59046 628632
rect 58622 616312 58678 616321
rect 58622 616247 58678 616256
rect 57886 604072 57942 604081
rect 57886 604007 57942 604016
rect 57900 569226 57928 604007
rect 58530 585712 58586 585721
rect 58530 585647 58586 585656
rect 58438 573472 58494 573481
rect 58438 573407 58494 573416
rect 57888 569220 57940 569226
rect 57888 569162 57940 569168
rect 57796 550316 57848 550322
rect 57796 550258 57848 550264
rect 56508 550180 56560 550186
rect 56508 550122 56560 550128
rect 56416 550044 56468 550050
rect 56416 549986 56468 549992
rect 54944 549976 54996 549982
rect 54944 549918 54996 549924
rect 57900 518226 57928 569162
rect 58452 555558 58480 573407
rect 58544 567934 58572 585647
rect 58532 567928 58584 567934
rect 58532 567870 58584 567876
rect 58440 555552 58492 555558
rect 58440 555494 58492 555500
rect 58636 554266 58664 616247
rect 58898 610192 58954 610201
rect 58898 610127 58954 610136
rect 58806 601352 58862 601361
rect 58806 601287 58862 601296
rect 58714 597952 58770 597961
rect 58714 597887 58770 597896
rect 58728 568478 58756 597887
rect 58716 568472 58768 568478
rect 58716 568414 58768 568420
rect 58820 568002 58848 601287
rect 58808 567996 58860 568002
rect 58808 567938 58860 567944
rect 58912 556850 58940 610127
rect 59004 566710 59032 628623
rect 59096 607617 59124 649266
rect 104912 647902 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 137744 683188 137796 683194
rect 137744 683130 137796 683136
rect 104900 647896 104952 647902
rect 104900 647838 104952 647844
rect 114192 634092 114244 634098
rect 114192 634034 114244 634040
rect 121644 634092 121696 634098
rect 121644 634034 121696 634040
rect 131120 634092 131172 634098
rect 131120 634034 131172 634040
rect 112536 633956 112588 633962
rect 112536 633898 112588 633904
rect 69296 633888 69348 633894
rect 69296 633830 69348 633836
rect 59360 631372 59412 631378
rect 59360 631314 59412 631320
rect 59268 630896 59320 630902
rect 59268 630838 59320 630844
rect 59174 625832 59230 625841
rect 59174 625767 59230 625776
rect 59082 607608 59138 607617
rect 59082 607543 59138 607552
rect 59082 582992 59138 583001
rect 59082 582927 59138 582936
rect 58992 566704 59044 566710
rect 58992 566646 59044 566652
rect 59096 566030 59124 582927
rect 59084 566024 59136 566030
rect 59084 565966 59136 565972
rect 59188 561066 59216 625767
rect 59176 561060 59228 561066
rect 59176 561002 59228 561008
rect 58900 556844 58952 556850
rect 58900 556786 58952 556792
rect 58624 554260 58676 554266
rect 58624 554202 58676 554208
rect 59280 550118 59308 630838
rect 59372 552786 59400 631314
rect 69308 630986 69336 633830
rect 106648 633820 106700 633826
rect 106648 633762 106700 633768
rect 77300 633684 77352 633690
rect 77300 633626 77352 633632
rect 104072 633684 104124 633690
rect 104072 633626 104124 633632
rect 69046 630958 69336 630986
rect 77312 630986 77340 633626
rect 88708 633616 88760 633622
rect 88708 633558 88760 633564
rect 100668 633616 100720 633622
rect 100668 633558 100720 633564
rect 88720 630986 88748 633558
rect 91836 633548 91888 633554
rect 91836 633490 91888 633496
rect 95056 633548 95108 633554
rect 95056 633490 95108 633496
rect 91848 630986 91876 633490
rect 95068 630986 95096 633490
rect 97724 631372 97776 631378
rect 97724 631314 97776 631320
rect 77312 630958 77418 630986
rect 80256 630970 80638 630986
rect 80244 630964 80638 630970
rect 80296 630958 80638 630964
rect 88720 630958 89010 630986
rect 91848 630958 92230 630986
rect 94806 630958 95096 630986
rect 97736 630986 97764 631314
rect 100680 630986 100708 633558
rect 104084 630986 104112 633626
rect 106660 630986 106688 633762
rect 109960 633480 110012 633486
rect 109960 633422 110012 633428
rect 109972 630986 110000 633422
rect 112548 630986 112576 633898
rect 114204 633690 114232 634034
rect 115664 634024 115716 634030
rect 115664 633966 115716 633972
rect 114192 633684 114244 633690
rect 114192 633626 114244 633632
rect 115676 630986 115704 633966
rect 121460 633820 121512 633826
rect 121460 633762 121512 633768
rect 118240 633684 118292 633690
rect 118240 633626 118292 633632
rect 118252 630986 118280 633626
rect 120908 633548 120960 633554
rect 120908 633490 120960 633496
rect 97736 630958 98026 630986
rect 100602 630958 100708 630986
rect 103822 630958 104112 630986
rect 106398 630958 106688 630986
rect 109618 630958 110000 630986
rect 112194 630958 112576 630986
rect 115414 630958 115704 630986
rect 117990 630958 118280 630986
rect 80244 630906 80296 630912
rect 65524 630896 65576 630902
rect 65576 630844 65826 630850
rect 65524 630838 65826 630844
rect 65536 630822 65826 630838
rect 71240 630834 71622 630850
rect 71228 630828 71622 630834
rect 71280 630822 71622 630828
rect 71228 630770 71280 630776
rect 74632 630760 74684 630766
rect 62960 630698 63250 630714
rect 86776 630760 86828 630766
rect 74684 630708 74842 630714
rect 74632 630702 74842 630708
rect 62948 630692 63250 630698
rect 63000 630686 63250 630692
rect 74644 630686 74842 630702
rect 83214 630698 83504 630714
rect 86434 630708 86776 630714
rect 86434 630702 86828 630708
rect 83214 630692 83516 630698
rect 83214 630686 83464 630692
rect 62948 630634 63000 630640
rect 86434 630686 86816 630702
rect 83464 630634 83516 630640
rect 59464 630414 60030 630442
rect 120566 630414 120764 630442
rect 59464 563786 59492 630414
rect 59542 570788 59598 570797
rect 59542 570723 59598 570732
rect 59452 563780 59504 563786
rect 59452 563722 59504 563728
rect 59556 552906 59584 570723
rect 59912 569152 59964 569158
rect 59912 569094 59964 569100
rect 59924 557534 59952 569094
rect 60740 568472 60792 568478
rect 60740 568414 60792 568420
rect 60030 568126 60320 568154
rect 60292 565078 60320 568126
rect 60280 565072 60332 565078
rect 60280 565014 60332 565020
rect 60752 557534 60780 568414
rect 61384 568404 61436 568410
rect 61384 568346 61436 568352
rect 59924 557506 60412 557534
rect 60752 557506 60964 557534
rect 59544 552900 59596 552906
rect 59544 552842 59596 552848
rect 59372 552758 60320 552786
rect 59268 550112 59320 550118
rect 59268 550054 59320 550060
rect 60292 547963 60320 552758
rect 60384 550254 60412 557506
rect 60372 550248 60424 550254
rect 60372 550190 60424 550196
rect 60936 547963 60964 557506
rect 61396 549914 61424 568346
rect 106280 568268 106332 568274
rect 106280 568210 106332 568216
rect 99564 568200 99616 568206
rect 62606 568126 62896 568154
rect 62120 566024 62172 566030
rect 62120 565966 62172 565972
rect 62132 557534 62160 565966
rect 62868 565146 62896 568126
rect 64984 568126 65182 568154
rect 68402 568126 68784 568154
rect 70978 568126 71360 568154
rect 64880 567860 64932 567866
rect 64880 567802 64932 567808
rect 62856 565140 62908 565146
rect 62856 565082 62908 565088
rect 62580 565072 62632 565078
rect 62580 565014 62632 565020
rect 62592 559638 62620 565014
rect 63500 563712 63552 563718
rect 63500 563654 63552 563660
rect 62580 559632 62632 559638
rect 62580 559574 62632 559580
rect 62132 557506 62436 557534
rect 61384 549908 61436 549914
rect 61384 549850 61436 549856
rect 61660 549364 61712 549370
rect 61660 549306 61712 549312
rect 61672 547963 61700 549306
rect 62408 547963 62436 557506
rect 63132 555484 63184 555490
rect 63132 555426 63184 555432
rect 63144 547963 63172 555426
rect 63512 552786 63540 563654
rect 63592 562352 63644 562358
rect 63592 562294 63644 562300
rect 63604 557534 63632 562294
rect 63604 557506 64552 557534
rect 63512 552758 63816 552786
rect 63788 547963 63816 552758
rect 64524 547963 64552 557506
rect 64892 549250 64920 567802
rect 64984 549370 65012 568126
rect 67640 567928 67692 567934
rect 67640 567870 67692 567876
rect 65064 559564 65116 559570
rect 65064 559506 65116 559512
rect 65076 557534 65104 559506
rect 66352 558204 66404 558210
rect 66352 558146 66404 558152
rect 66364 557534 66392 558146
rect 65076 557506 66024 557534
rect 66364 557506 66760 557534
rect 64972 549364 65024 549370
rect 64972 549306 65024 549312
rect 64892 549222 65288 549250
rect 65260 547963 65288 549222
rect 65996 547963 66024 557506
rect 66732 547963 66760 557506
rect 67652 552770 67680 567870
rect 67732 566500 67784 566506
rect 67732 566442 67784 566448
rect 67744 557534 67772 566442
rect 68756 565282 68784 568126
rect 69020 566568 69072 566574
rect 69020 566510 69072 566516
rect 68744 565276 68796 565282
rect 68744 565218 68796 565224
rect 67744 557506 68140 557534
rect 67640 552764 67692 552770
rect 67640 552706 67692 552712
rect 67364 550452 67416 550458
rect 67364 550394 67416 550400
rect 67376 547963 67404 550394
rect 68112 547963 68140 557506
rect 69032 552770 69060 566510
rect 71332 565214 71360 568126
rect 73816 568126 74198 568154
rect 76774 568126 77064 568154
rect 71320 565208 71372 565214
rect 71320 565150 71372 565156
rect 72424 565140 72476 565146
rect 72424 565082 72476 565088
rect 71780 564460 71832 564466
rect 71780 564402 71832 564408
rect 70400 560992 70452 560998
rect 70400 560934 70452 560940
rect 69572 554056 69624 554062
rect 69572 553998 69624 554004
rect 68836 552764 68888 552770
rect 68836 552706 68888 552712
rect 69020 552764 69072 552770
rect 69020 552706 69072 552712
rect 68848 547963 68876 552706
rect 69584 547963 69612 553998
rect 70412 552786 70440 560934
rect 70492 558272 70544 558278
rect 70492 558214 70544 558220
rect 70504 552906 70532 558214
rect 70492 552900 70544 552906
rect 70492 552842 70544 552848
rect 71688 552900 71740 552906
rect 71688 552842 71740 552848
rect 70308 552764 70360 552770
rect 70412 552758 70992 552786
rect 70308 552706 70360 552712
rect 70320 547963 70348 552706
rect 70964 547963 70992 552758
rect 71700 547963 71728 552842
rect 71792 552786 71820 564402
rect 72436 554130 72464 565082
rect 73816 564466 73844 568126
rect 74540 565412 74592 565418
rect 74540 565354 74592 565360
rect 73804 564460 73856 564466
rect 73804 564402 73856 564408
rect 74552 557534 74580 565354
rect 77036 565350 77064 568126
rect 78876 568126 79994 568154
rect 82570 568126 82768 568154
rect 85790 568126 86080 568154
rect 88366 568126 88656 568154
rect 78772 568064 78824 568070
rect 78772 568006 78824 568012
rect 78680 567928 78732 567934
rect 78680 567870 78732 567876
rect 77300 566704 77352 566710
rect 77300 566646 77352 566652
rect 77024 565344 77076 565350
rect 77024 565286 77076 565292
rect 75920 565140 75972 565146
rect 75920 565082 75972 565088
rect 74552 557506 75316 557534
rect 74540 554260 74592 554266
rect 74540 554202 74592 554208
rect 73160 554192 73212 554198
rect 73160 554134 73212 554140
rect 72424 554124 72476 554130
rect 72424 554066 72476 554072
rect 71792 552758 72464 552786
rect 72436 547963 72464 552758
rect 73172 547963 73200 554134
rect 73804 550044 73856 550050
rect 73804 549986 73856 549992
rect 73816 547963 73844 549986
rect 74552 547963 74580 554202
rect 75288 547963 75316 557506
rect 75932 552770 75960 565082
rect 76012 563780 76064 563786
rect 76012 563722 76064 563728
rect 75920 552764 75972 552770
rect 75920 552706 75972 552712
rect 76024 547963 76052 563722
rect 77312 557534 77340 566646
rect 77312 557506 77432 557534
rect 76748 552764 76800 552770
rect 76748 552706 76800 552712
rect 76760 547963 76788 552706
rect 77404 547963 77432 557506
rect 78692 552786 78720 567870
rect 78784 552922 78812 568006
rect 78876 556918 78904 568126
rect 82740 565486 82768 568126
rect 84200 566704 84252 566710
rect 84200 566646 84252 566652
rect 82912 566636 82964 566642
rect 82912 566578 82964 566584
rect 82728 565480 82780 565486
rect 82728 565422 82780 565428
rect 80060 563780 80112 563786
rect 80060 563722 80112 563728
rect 78864 556912 78916 556918
rect 78864 556854 78916 556860
rect 78784 552894 78996 552922
rect 78968 552786 78996 552894
rect 80072 552786 80100 563722
rect 80152 562488 80204 562494
rect 80152 562430 80204 562436
rect 80164 557534 80192 562430
rect 82924 557534 82952 566578
rect 84212 557534 84240 566646
rect 86052 565350 86080 568126
rect 87052 566840 87104 566846
rect 87052 566782 87104 566788
rect 86960 566636 87012 566642
rect 86960 566578 87012 566584
rect 84844 565344 84896 565350
rect 84844 565286 84896 565292
rect 86040 565344 86092 565350
rect 86040 565286 86092 565292
rect 80164 557506 81020 557534
rect 82924 557506 83228 557534
rect 84212 557506 84608 557534
rect 78692 552758 78904 552786
rect 78968 552758 79640 552786
rect 80072 552758 80376 552786
rect 78128 550044 78180 550050
rect 78128 549986 78180 549992
rect 78140 547963 78168 549986
rect 78876 547963 78904 552758
rect 79612 547963 79640 552758
rect 80348 547963 80376 552758
rect 80992 547963 81020 557506
rect 81716 552832 81768 552838
rect 81716 552774 81768 552780
rect 81728 547963 81756 552774
rect 82452 552764 82504 552770
rect 82452 552706 82504 552712
rect 82464 547963 82492 552706
rect 83200 547963 83228 557506
rect 83924 550180 83976 550186
rect 83924 550122 83976 550128
rect 83936 547963 83964 550122
rect 84580 547963 84608 557506
rect 84856 550594 84884 565286
rect 85672 563848 85724 563854
rect 85672 563790 85724 563796
rect 85684 557534 85712 563790
rect 85684 557506 86080 557534
rect 84844 550588 84896 550594
rect 84844 550530 84896 550536
rect 85304 550180 85356 550186
rect 85304 550122 85356 550128
rect 85316 547963 85344 550122
rect 86052 547963 86080 557506
rect 86972 552838 87000 566578
rect 87064 557534 87092 566782
rect 87604 563916 87656 563922
rect 87604 563858 87656 563864
rect 87064 557506 87460 557534
rect 86960 552832 87012 552838
rect 86960 552774 87012 552780
rect 86776 550588 86828 550594
rect 86776 550530 86828 550536
rect 86788 547963 86816 550530
rect 87432 547963 87460 557506
rect 87616 550594 87644 563858
rect 88628 561134 88656 568126
rect 91204 568126 91586 568154
rect 94162 568126 94544 568154
rect 91100 567996 91152 568002
rect 91100 567938 91152 567944
rect 89812 565480 89864 565486
rect 89812 565422 89864 565428
rect 88616 561128 88668 561134
rect 88616 561070 88668 561076
rect 88432 559768 88484 559774
rect 88432 559710 88484 559716
rect 88444 552838 88472 559710
rect 89824 557534 89852 565422
rect 89824 557506 90404 557534
rect 88156 552832 88208 552838
rect 88156 552774 88208 552780
rect 88432 552832 88484 552838
rect 88432 552774 88484 552780
rect 89628 552832 89680 552838
rect 89628 552774 89680 552780
rect 87604 550588 87656 550594
rect 87604 550530 87656 550536
rect 88168 547963 88196 552774
rect 88892 550384 88944 550390
rect 88892 550326 88944 550332
rect 88904 547963 88932 550326
rect 89640 547963 89668 552774
rect 89720 551336 89772 551342
rect 89720 551278 89772 551284
rect 89732 550390 89760 551278
rect 89720 550384 89772 550390
rect 89720 550326 89772 550332
rect 90376 547963 90404 557506
rect 91008 550588 91060 550594
rect 91008 550530 91060 550536
rect 91020 547963 91048 550530
rect 91112 550338 91140 567938
rect 91204 550458 91232 568126
rect 93860 568064 93912 568070
rect 93860 568006 93912 568012
rect 92572 561060 92624 561066
rect 92572 561002 92624 561008
rect 91192 550452 91244 550458
rect 91192 550394 91244 550400
rect 91112 550310 91784 550338
rect 91756 547963 91784 550310
rect 92584 548162 92612 561002
rect 93872 557534 93900 568006
rect 94516 564942 94544 568126
rect 96712 568132 96764 568138
rect 96712 568074 96764 568080
rect 97000 568126 97382 568154
rect 99564 568142 99616 568148
rect 94504 564936 94556 564942
rect 94504 564878 94556 564884
rect 96724 557534 96752 568074
rect 97000 565418 97028 568126
rect 98092 567996 98144 568002
rect 98092 567938 98144 567944
rect 96988 565412 97040 565418
rect 96988 565354 97040 565360
rect 98104 557534 98132 567938
rect 99576 557534 99604 568142
rect 99958 568126 100248 568154
rect 100220 565418 100248 568126
rect 102888 568126 103178 568154
rect 104912 568126 105754 568154
rect 100208 565412 100260 565418
rect 100208 565354 100260 565360
rect 102784 564936 102836 564942
rect 102784 564878 102836 564884
rect 100760 564460 100812 564466
rect 100760 564402 100812 564408
rect 100772 557534 100800 564402
rect 93872 557506 93992 557534
rect 96724 557506 97488 557534
rect 98104 557506 98224 557534
rect 99576 557506 100432 557534
rect 100772 557506 101812 557534
rect 93216 550316 93268 550322
rect 93216 550258 93268 550264
rect 92508 548134 92612 548162
rect 92508 547944 92536 548134
rect 93228 547963 93256 550258
rect 93964 547963 93992 557506
rect 94596 555620 94648 555626
rect 94596 555562 94648 555568
rect 94608 547963 94636 555562
rect 96804 550452 96856 550458
rect 96804 550394 96856 550400
rect 96068 550316 96120 550322
rect 96068 550258 96120 550264
rect 95332 550248 95384 550254
rect 95332 550190 95384 550196
rect 95344 547963 95372 550190
rect 96080 547963 96108 550258
rect 96816 547963 96844 550394
rect 97460 547963 97488 557506
rect 98092 552832 98144 552838
rect 98092 552774 98144 552780
rect 98104 550322 98132 552774
rect 98092 550316 98144 550322
rect 98092 550258 98144 550264
rect 98196 547963 98224 557506
rect 98920 550112 98972 550118
rect 98920 550054 98972 550060
rect 98932 547963 98960 550054
rect 99656 549976 99708 549982
rect 99656 549918 99708 549924
rect 99668 547963 99696 549918
rect 100404 547963 100432 557506
rect 101036 552696 101088 552702
rect 101036 552638 101088 552644
rect 101048 547963 101076 552638
rect 101784 547963 101812 557506
rect 102508 556844 102560 556850
rect 102508 556786 102560 556792
rect 102520 547963 102548 556786
rect 102796 549370 102824 564878
rect 102888 564466 102916 568126
rect 102876 564460 102928 564466
rect 102876 564402 102928 564408
rect 103520 561128 103572 561134
rect 103520 561070 103572 561076
rect 103532 557534 103560 561070
rect 104912 559774 104940 568126
rect 105544 565276 105596 565282
rect 105544 565218 105596 565224
rect 104900 559768 104952 559774
rect 104900 559710 104952 559716
rect 104992 559632 105044 559638
rect 104992 559574 105044 559580
rect 105004 557534 105032 559574
rect 103532 557506 104664 557534
rect 105004 557506 105400 557534
rect 103244 555552 103296 555558
rect 103244 555494 103296 555500
rect 102784 549364 102836 549370
rect 102784 549306 102836 549312
rect 103256 547963 103284 555494
rect 103980 549976 104032 549982
rect 103980 549918 104032 549924
rect 103992 547963 104020 549918
rect 104636 547963 104664 557506
rect 105372 547963 105400 557506
rect 105556 550526 105584 565218
rect 106292 552702 106320 568210
rect 108592 568126 108974 568154
rect 110616 568126 111550 568154
rect 114572 568126 114770 568154
rect 117346 568126 117452 568154
rect 108304 565344 108356 565350
rect 108304 565286 108356 565292
rect 106924 564460 106976 564466
rect 106924 564402 106976 564408
rect 106936 554198 106964 564402
rect 107752 558340 107804 558346
rect 107752 558282 107804 558288
rect 107764 557534 107792 558282
rect 107764 557506 108252 557534
rect 106924 554192 106976 554198
rect 106924 554134 106976 554140
rect 106280 552696 106332 552702
rect 106280 552638 106332 552644
rect 107568 552696 107620 552702
rect 107568 552638 107620 552644
rect 105544 550520 105596 550526
rect 105544 550462 105596 550468
rect 106832 550112 106884 550118
rect 106832 550054 106884 550060
rect 106096 549364 106148 549370
rect 106096 549306 106148 549312
rect 106108 547963 106136 549306
rect 106844 547963 106872 550054
rect 107580 547963 107608 552638
rect 108224 547963 108252 557506
rect 108316 550594 108344 565286
rect 108396 565208 108448 565214
rect 108396 565150 108448 565156
rect 108304 550588 108356 550594
rect 108304 550530 108356 550536
rect 108408 549370 108436 565150
rect 108592 564466 108620 568126
rect 110420 565208 110472 565214
rect 110420 565150 110472 565156
rect 108580 564460 108632 564466
rect 108580 564402 108632 564408
rect 109684 554124 109736 554130
rect 109684 554066 109736 554072
rect 108948 550520 109000 550526
rect 108948 550462 109000 550468
rect 108396 549364 108448 549370
rect 108396 549306 108448 549312
rect 108960 547963 108988 550462
rect 109696 547963 109724 554066
rect 110432 547963 110460 565150
rect 110512 562420 110564 562426
rect 110512 562362 110564 562368
rect 110524 552786 110552 562362
rect 110616 555490 110644 568126
rect 111892 566772 111944 566778
rect 111892 566714 111944 566720
rect 111904 557534 111932 566714
rect 113180 564528 113232 564534
rect 113180 564470 113232 564476
rect 113192 557534 113220 564470
rect 111904 557506 112576 557534
rect 113192 557506 113312 557534
rect 110604 555484 110656 555490
rect 110604 555426 110656 555432
rect 110524 552758 111104 552786
rect 111076 547963 111104 552758
rect 111800 550588 111852 550594
rect 111800 550530 111852 550536
rect 111812 547963 111840 550530
rect 112548 547963 112576 557506
rect 113284 547963 113312 557506
rect 114572 554062 114600 568126
rect 115204 565412 115256 565418
rect 115204 565354 115256 565360
rect 114560 554056 114612 554062
rect 114560 553998 114612 554004
rect 115216 550594 115244 565354
rect 117424 565146 117452 568126
rect 120184 568126 120566 568154
rect 118700 565276 118752 565282
rect 118700 565218 118752 565224
rect 117412 565140 117464 565146
rect 117412 565082 117464 565088
rect 116584 564460 116636 564466
rect 116584 564402 116636 564408
rect 115388 556912 115440 556918
rect 115388 556854 115440 556860
rect 115204 550588 115256 550594
rect 115204 550530 115256 550536
rect 114008 550248 114060 550254
rect 114008 550190 114060 550196
rect 114020 547963 114048 550190
rect 114652 549364 114704 549370
rect 114652 549306 114704 549312
rect 114664 547963 114692 549306
rect 115400 547963 115428 556854
rect 116596 552770 116624 564402
rect 118712 557534 118740 565218
rect 120184 564466 120212 568126
rect 120736 565214 120764 630414
rect 120814 608968 120870 608977
rect 120814 608903 120870 608912
rect 120724 565208 120776 565214
rect 120724 565150 120776 565156
rect 120172 564460 120224 564466
rect 120172 564402 120224 564408
rect 120172 562556 120224 562562
rect 120172 562498 120224 562504
rect 120184 557534 120212 562498
rect 120828 560998 120856 608903
rect 120816 560992 120868 560998
rect 120816 560934 120868 560940
rect 118712 557506 119752 557534
rect 120184 557506 120856 557534
rect 116584 552764 116636 552770
rect 116584 552706 116636 552712
rect 116124 550588 116176 550594
rect 116124 550530 116176 550536
rect 116136 547963 116164 550530
rect 117596 550384 117648 550390
rect 117596 550326 117648 550332
rect 116860 549908 116912 549914
rect 116860 549850 116912 549856
rect 116872 547963 116900 549850
rect 117608 547963 117636 550326
rect 118976 550316 119028 550322
rect 118976 550258 119028 550264
rect 118240 549364 118292 549370
rect 118240 549306 118292 549312
rect 118252 547963 118280 549306
rect 118988 547963 119016 550258
rect 119724 547963 119752 557506
rect 120448 551336 120500 551342
rect 120448 551278 120500 551284
rect 120460 547963 120488 551278
rect 120828 550066 120856 557506
rect 120920 550186 120948 633490
rect 121000 633480 121052 633486
rect 121000 633422 121052 633428
rect 121012 568002 121040 633422
rect 121090 591220 121146 591229
rect 121090 591155 121146 591164
rect 121000 567996 121052 568002
rect 121000 567938 121052 567944
rect 121104 562494 121132 591155
rect 121182 572860 121238 572869
rect 121182 572795 121238 572804
rect 121196 564534 121224 572795
rect 121472 566846 121500 633762
rect 121550 625288 121606 625297
rect 121550 625223 121606 625232
rect 121460 566840 121512 566846
rect 121460 566782 121512 566788
rect 121564 566778 121592 625223
rect 121552 566772 121604 566778
rect 121552 566714 121604 566720
rect 121184 564528 121236 564534
rect 121184 564470 121236 564476
rect 121092 562488 121144 562494
rect 121092 562430 121144 562436
rect 120908 550180 120960 550186
rect 120908 550122 120960 550128
rect 120828 550038 121132 550066
rect 121656 550050 121684 634034
rect 124588 634024 124640 634030
rect 124588 633966 124640 633972
rect 123024 633956 123076 633962
rect 123024 633898 123076 633904
rect 122840 633752 122892 633758
rect 122840 633694 122892 633700
rect 121826 621208 121882 621217
rect 121826 621143 121882 621152
rect 121734 615632 121790 615641
rect 121734 615567 121790 615576
rect 121748 558278 121776 615567
rect 121840 563854 121868 621143
rect 121918 618488 121974 618497
rect 121918 618423 121974 618432
rect 121932 566506 121960 618423
rect 122010 600400 122066 600409
rect 122010 600335 122066 600344
rect 121920 566500 121972 566506
rect 121920 566442 121972 566448
rect 121828 563848 121880 563854
rect 121828 563790 121880 563796
rect 121736 558272 121788 558278
rect 121736 558214 121788 558220
rect 122024 555626 122052 600335
rect 122102 588024 122158 588033
rect 122102 587959 122158 587968
rect 122116 566710 122144 587959
rect 122194 581768 122250 581777
rect 122194 581703 122250 581712
rect 122208 568206 122236 581703
rect 122286 578368 122342 578377
rect 122286 578303 122342 578312
rect 122196 568200 122248 568206
rect 122196 568142 122248 568148
rect 122196 567996 122248 568002
rect 122196 567938 122248 567944
rect 122104 566704 122156 566710
rect 122104 566646 122156 566652
rect 122208 557534 122236 567938
rect 122300 567934 122328 578303
rect 122852 568070 122880 633694
rect 122930 628008 122986 628017
rect 122930 627943 122986 627952
rect 122840 568064 122892 568070
rect 122840 568006 122892 568012
rect 122288 567928 122340 567934
rect 122288 567870 122340 567876
rect 122840 563848 122892 563854
rect 122840 563790 122892 563796
rect 122208 557506 122604 557534
rect 122012 555620 122064 555626
rect 122012 555562 122064 555568
rect 121828 555484 121880 555490
rect 121828 555426 121880 555432
rect 121104 547963 121132 550038
rect 121644 550044 121696 550050
rect 121644 549986 121696 549992
rect 121840 547963 121868 555426
rect 122576 547963 122604 557506
rect 122852 552786 122880 563790
rect 122944 562358 122972 627943
rect 123036 568138 123064 633898
rect 124312 633684 124364 633690
rect 124312 633626 124364 633632
rect 124220 633616 124272 633622
rect 124220 633558 124272 633564
rect 123114 612776 123170 612785
rect 123114 612711 123170 612720
rect 123024 568132 123076 568138
rect 123024 568074 123076 568080
rect 122932 562352 122984 562358
rect 122932 562294 122984 562300
rect 122932 559632 122984 559638
rect 122932 559574 122984 559580
rect 122944 552906 122972 559574
rect 123128 559570 123156 612711
rect 123298 606248 123354 606257
rect 123298 606183 123354 606192
rect 123206 603120 123262 603129
rect 123206 603055 123262 603064
rect 123116 559564 123168 559570
rect 123116 559506 123168 559512
rect 123220 552974 123248 603055
rect 123312 563786 123340 606183
rect 124126 596728 124182 596737
rect 124126 596663 124182 596672
rect 124140 596222 124168 596663
rect 124128 596216 124180 596222
rect 124128 596158 124180 596164
rect 123390 594008 123446 594017
rect 123390 593943 123446 593952
rect 123404 567866 123432 593943
rect 123482 584488 123538 584497
rect 123482 584423 123538 584432
rect 123392 567860 123444 567866
rect 123392 567802 123444 567808
rect 123496 566574 123524 584423
rect 123666 575648 123722 575657
rect 123666 575583 123722 575592
rect 123574 570072 123630 570081
rect 123574 570007 123630 570016
rect 123484 566568 123536 566574
rect 123484 566510 123536 566516
rect 123300 563780 123352 563786
rect 123300 563722 123352 563728
rect 123588 558210 123616 570007
rect 123680 563718 123708 575583
rect 123668 563712 123720 563718
rect 123668 563654 123720 563660
rect 123576 558204 123628 558210
rect 123576 558146 123628 558152
rect 124232 556510 124260 633558
rect 124324 566642 124352 633626
rect 124496 630760 124548 630766
rect 124496 630702 124548 630708
rect 124404 630692 124456 630698
rect 124404 630634 124456 630640
rect 124312 566636 124364 566642
rect 124312 566578 124364 566584
rect 124312 558272 124364 558278
rect 124312 558214 124364 558220
rect 124220 556504 124272 556510
rect 124220 556446 124272 556452
rect 123208 552968 123260 552974
rect 123208 552910 123260 552916
rect 122932 552900 122984 552906
rect 122932 552842 122984 552848
rect 124036 552900 124088 552906
rect 124036 552842 124088 552848
rect 122852 552758 123340 552786
rect 123312 547963 123340 552758
rect 124048 547963 124076 552842
rect 124324 549794 124352 558214
rect 124416 550118 124444 630634
rect 124404 550112 124456 550118
rect 124404 550054 124456 550060
rect 124508 549982 124536 630702
rect 124600 568274 124628 633966
rect 127072 633888 127124 633894
rect 127072 633830 127124 633836
rect 124864 631032 124916 631038
rect 124864 630974 124916 630980
rect 124588 568268 124640 568274
rect 124588 568210 124640 568216
rect 124496 549976 124548 549982
rect 124496 549918 124548 549924
rect 124324 549766 124720 549794
rect 124692 547963 124720 549766
rect 124876 549370 124904 630974
rect 126244 597576 126296 597582
rect 126244 597518 126296 597524
rect 125600 585200 125652 585206
rect 125600 585142 125652 585148
rect 125416 556504 125468 556510
rect 125416 556446 125468 556452
rect 124864 549364 124916 549370
rect 124864 549306 124916 549312
rect 125428 547963 125456 556446
rect 125612 552770 125640 585142
rect 125692 566772 125744 566778
rect 125692 566714 125744 566720
rect 125704 557534 125732 566714
rect 125704 557506 126192 557534
rect 125600 552764 125652 552770
rect 125600 552706 125652 552712
rect 126164 547963 126192 557506
rect 126256 550322 126284 597518
rect 126980 562488 127032 562494
rect 126980 562430 127032 562436
rect 126992 556374 127020 562430
rect 126980 556368 127032 556374
rect 126980 556310 127032 556316
rect 126888 552764 126940 552770
rect 126888 552706 126940 552712
rect 126244 550316 126296 550322
rect 126244 550258 126296 550264
rect 126900 547963 126928 552706
rect 127084 550254 127112 633830
rect 129004 582412 129056 582418
rect 129004 582354 129056 582360
rect 128360 563916 128412 563922
rect 128360 563858 128412 563864
rect 128268 556368 128320 556374
rect 128268 556310 128320 556316
rect 127624 552696 127676 552702
rect 127624 552638 127676 552644
rect 127072 550248 127124 550254
rect 127072 550190 127124 550196
rect 127636 547963 127664 552638
rect 128280 547963 128308 556310
rect 128372 552786 128400 563858
rect 129016 557534 129044 582354
rect 129740 565344 129792 565350
rect 129740 565286 129792 565292
rect 129016 557506 129136 557534
rect 128372 552758 129044 552786
rect 129016 547963 129044 552758
rect 129108 551342 129136 557506
rect 129752 552770 129780 565286
rect 129832 559700 129884 559706
rect 129832 559642 129884 559648
rect 129740 552764 129792 552770
rect 129740 552706 129792 552712
rect 129096 551336 129148 551342
rect 129096 551278 129148 551284
rect 129844 548162 129872 559642
rect 131132 557534 131160 634034
rect 135260 634024 135312 634030
rect 135260 633966 135312 633972
rect 135168 633956 135220 633962
rect 135168 633898 135220 633904
rect 134892 633684 134944 633690
rect 134892 633626 134944 633632
rect 133880 633480 133932 633486
rect 133880 633422 133932 633428
rect 132500 615936 132552 615942
rect 132500 615878 132552 615884
rect 131132 557506 131896 557534
rect 130476 552764 130528 552770
rect 130476 552706 130528 552712
rect 129768 548134 129872 548162
rect 129768 547944 129796 548134
rect 130488 547963 130516 552706
rect 131212 549364 131264 549370
rect 131212 549306 131264 549312
rect 131224 547963 131252 549306
rect 131868 547963 131896 557506
rect 132512 552786 132540 615878
rect 132592 565140 132644 565146
rect 132592 565082 132644 565088
rect 132604 557534 132632 565082
rect 132604 557506 133368 557534
rect 132512 552758 132632 552786
rect 132604 547963 132632 552758
rect 133340 547963 133368 557506
rect 133892 557002 133920 633422
rect 134524 596216 134576 596222
rect 134524 596158 134576 596164
rect 134536 568478 134564 596158
rect 134524 568472 134576 568478
rect 134524 568414 134576 568420
rect 134904 568070 134932 633626
rect 134984 631100 135036 631106
rect 134984 631042 135036 631048
rect 134892 568064 134944 568070
rect 134892 568006 134944 568012
rect 133972 565208 134024 565214
rect 133972 565150 134024 565156
rect 133984 557534 134012 565150
rect 134524 558340 134576 558346
rect 134524 558282 134576 558288
rect 133984 557506 134196 557534
rect 133892 556974 134104 557002
rect 134076 547963 134104 556974
rect 134168 549250 134196 557506
rect 134536 549370 134564 558282
rect 134996 550526 135024 631042
rect 135076 630896 135128 630902
rect 135076 630838 135128 630844
rect 134984 550520 135036 550526
rect 134984 550462 135036 550468
rect 135088 550322 135116 630838
rect 135180 550390 135208 633898
rect 135272 557534 135300 633966
rect 136548 633888 136600 633894
rect 136548 633830 136600 633836
rect 136456 630964 136508 630970
rect 136456 630906 136508 630912
rect 135272 557506 136220 557534
rect 135444 550588 135496 550594
rect 135444 550530 135496 550536
rect 135168 550384 135220 550390
rect 135168 550326 135220 550332
rect 135076 550316 135128 550322
rect 135076 550258 135128 550264
rect 134524 549364 134576 549370
rect 134524 549306 134576 549312
rect 134168 549222 134748 549250
rect 134720 547963 134748 549222
rect 135456 547963 135484 550530
rect 136192 547963 136220 557506
rect 136468 550050 136496 630906
rect 136560 550118 136588 633830
rect 137652 633548 137704 633554
rect 137652 633490 137704 633496
rect 136640 630828 136692 630834
rect 136640 630770 136692 630776
rect 136652 557534 136680 630770
rect 137282 628688 137338 628697
rect 137282 628623 137338 628632
rect 136730 616312 136786 616321
rect 136730 616247 136786 616256
rect 136744 615942 136772 616247
rect 136732 615936 136784 615942
rect 136732 615878 136784 615884
rect 136730 597952 136786 597961
rect 136730 597887 136786 597896
rect 136744 597582 136772 597887
rect 136732 597576 136784 597582
rect 136732 597518 136784 597524
rect 136730 585712 136786 585721
rect 136730 585647 136786 585656
rect 136744 585206 136772 585647
rect 136732 585200 136784 585206
rect 136732 585142 136784 585148
rect 136730 582992 136786 583001
rect 136730 582927 136786 582936
rect 136744 582418 136772 582927
rect 136732 582412 136784 582418
rect 136732 582354 136784 582360
rect 137190 573472 137246 573481
rect 137190 573407 137246 573416
rect 137204 566506 137232 573407
rect 137192 566500 137244 566506
rect 137192 566442 137244 566448
rect 136652 557506 137140 557534
rect 136916 554124 136968 554130
rect 136916 554066 136968 554072
rect 136548 550112 136600 550118
rect 136548 550054 136600 550060
rect 136456 550044 136508 550050
rect 136456 549986 136508 549992
rect 136928 547963 136956 554066
rect 137112 550474 137140 557506
rect 137296 550594 137324 628623
rect 137558 619712 137614 619721
rect 137558 619647 137614 619656
rect 137374 595232 137430 595241
rect 137374 595167 137430 595176
rect 137388 569906 137416 595167
rect 137466 579728 137522 579737
rect 137466 579663 137522 579672
rect 137376 569900 137428 569906
rect 137376 569842 137428 569848
rect 137480 552922 137508 579663
rect 137572 566302 137600 619647
rect 137664 568206 137692 633490
rect 137756 607617 137784 683130
rect 169772 645182 169800 702406
rect 235184 700330 235212 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 299492 646542 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 304264 700324 304316 700330
rect 304264 700266 304316 700272
rect 299480 646536 299532 646542
rect 299480 646478 299532 646484
rect 169760 645176 169812 645182
rect 169760 645118 169812 645124
rect 284944 643136 284996 643142
rect 284944 643078 284996 643084
rect 280986 640384 281042 640393
rect 280986 640319 281042 640328
rect 280712 639668 280764 639674
rect 280712 639610 280764 639616
rect 219164 639124 219216 639130
rect 219164 639066 219216 639072
rect 218704 638988 218756 638994
rect 218704 638930 218756 638936
rect 151268 634092 151320 634098
rect 151268 634034 151320 634040
rect 210424 634092 210476 634098
rect 210424 634034 210476 634040
rect 139124 633820 139176 633826
rect 139124 633762 139176 633768
rect 137836 630760 137888 630766
rect 137836 630702 137888 630708
rect 137742 607608 137798 607617
rect 137742 607543 137798 607552
rect 137742 591832 137798 591841
rect 137742 591767 137798 591776
rect 137652 568200 137704 568206
rect 137652 568142 137704 568148
rect 137560 566296 137612 566302
rect 137560 566238 137612 566244
rect 137756 554418 137784 591767
rect 137848 557534 137876 630702
rect 137928 630692 137980 630698
rect 137928 630634 137980 630640
rect 137940 604081 137968 630634
rect 139030 625832 139086 625841
rect 139030 625767 139086 625776
rect 138938 613592 138994 613601
rect 138938 613527 138994 613536
rect 138846 610192 138902 610201
rect 138846 610127 138902 610136
rect 137926 604072 137982 604081
rect 137926 604007 137982 604016
rect 137940 603106 137968 604007
rect 137940 603078 138060 603106
rect 137926 601352 137982 601361
rect 137926 601287 137982 601296
rect 137940 558210 137968 601287
rect 138032 569226 138060 603078
rect 138754 589112 138810 589121
rect 138754 589047 138810 589056
rect 138662 576872 138718 576881
rect 138662 576807 138718 576816
rect 138572 572348 138624 572354
rect 138572 572290 138624 572296
rect 138020 569220 138072 569226
rect 138020 569162 138072 569168
rect 138584 567866 138612 572290
rect 138572 567860 138624 567866
rect 138572 567802 138624 567808
rect 138676 559570 138704 576807
rect 138768 562426 138796 589047
rect 138860 563718 138888 610127
rect 138848 563712 138900 563718
rect 138848 563654 138900 563660
rect 138756 562420 138808 562426
rect 138756 562362 138808 562368
rect 138952 560998 138980 613527
rect 139044 568138 139072 625767
rect 139136 572354 139164 633762
rect 139216 633752 139268 633758
rect 139216 633694 139268 633700
rect 139124 572348 139176 572354
rect 139124 572290 139176 572296
rect 139228 572234 139256 633694
rect 140136 633548 140188 633554
rect 140136 633490 140188 633496
rect 139676 633480 139728 633486
rect 139676 633422 139728 633428
rect 139688 630850 139716 633422
rect 139688 630822 140070 630850
rect 140148 630426 140176 633490
rect 142988 631100 143040 631106
rect 142988 631042 143040 631048
rect 143000 630986 143028 631042
rect 151280 630986 151308 634034
rect 183560 634024 183612 634030
rect 183560 633966 183612 633972
rect 160284 633956 160336 633962
rect 160284 633898 160336 633904
rect 157524 633548 157576 633554
rect 157524 633490 157576 633496
rect 157536 630986 157564 633490
rect 143000 630958 143290 630986
rect 149086 630970 149192 630986
rect 149086 630964 149204 630970
rect 149086 630958 149152 630964
rect 151280 630958 151662 630986
rect 157458 630958 157564 630986
rect 160296 630986 160324 633898
rect 162860 633888 162912 633894
rect 162860 633830 162912 633836
rect 162872 630986 162900 633830
rect 166172 633820 166224 633826
rect 166172 633762 166224 633768
rect 166184 630986 166212 633762
rect 174452 633752 174504 633758
rect 174452 633694 174504 633700
rect 171876 633616 171928 633622
rect 171876 633558 171928 633564
rect 171888 630986 171916 633558
rect 174464 630986 174492 633694
rect 180340 633684 180392 633690
rect 180340 633626 180392 633632
rect 178132 631032 178184 631038
rect 160296 630958 160678 630986
rect 162872 630958 163254 630986
rect 166184 630958 166474 630986
rect 171888 630958 172270 630986
rect 174464 630958 174846 630986
rect 178066 630980 178132 630986
rect 178066 630974 178184 630980
rect 180352 630986 180380 633626
rect 183572 630986 183600 633966
rect 190000 633684 190052 633690
rect 190000 633626 190052 633632
rect 204444 633684 204496 633690
rect 204444 633626 204496 633632
rect 209780 633684 209832 633690
rect 209780 633626 209832 633632
rect 186504 633480 186556 633486
rect 186504 633422 186556 633428
rect 178066 630958 178172 630974
rect 180352 630958 180642 630986
rect 183572 630958 183862 630986
rect 149152 630906 149204 630912
rect 154580 630896 154632 630902
rect 186516 630850 186544 633422
rect 190012 630986 190040 633626
rect 192576 633548 192628 633554
rect 192576 633490 192628 633496
rect 201684 633548 201736 633554
rect 201684 633490 201736 633496
rect 192588 630986 192616 633490
rect 195704 633480 195756 633486
rect 195704 633422 195756 633428
rect 200856 633480 200908 633486
rect 200856 633422 200908 633428
rect 195716 630986 195744 633422
rect 189658 630958 190040 630986
rect 192234 630958 192616 630986
rect 195454 630958 195744 630986
rect 154632 630844 154882 630850
rect 154580 630838 154882 630844
rect 154592 630822 154882 630838
rect 168760 630834 169050 630850
rect 168748 630828 169050 630834
rect 168800 630822 169050 630828
rect 186438 630822 186544 630850
rect 168748 630770 168800 630776
rect 145564 630760 145616 630766
rect 145616 630708 145866 630714
rect 145564 630702 145866 630708
rect 145576 630686 145866 630702
rect 198030 630426 198320 630442
rect 139860 630420 139912 630426
rect 139860 630362 139912 630368
rect 140136 630420 140188 630426
rect 198030 630420 198332 630426
rect 198030 630414 198280 630420
rect 140136 630362 140188 630368
rect 200606 630414 200712 630442
rect 198280 630362 198332 630368
rect 139306 622432 139362 622441
rect 139306 622367 139362 622376
rect 139136 572206 139256 572234
rect 139032 568132 139084 568138
rect 139032 568074 139084 568080
rect 139136 567662 139164 572206
rect 139214 570752 139270 570761
rect 139214 570687 139270 570696
rect 139228 567934 139256 570687
rect 139216 567928 139268 567934
rect 139216 567870 139268 567876
rect 139124 567656 139176 567662
rect 139124 567598 139176 567604
rect 138940 560992 138992 560998
rect 138940 560934 138992 560940
rect 138664 559564 138716 559570
rect 138664 559506 138716 559512
rect 137928 558204 137980 558210
rect 137928 558146 137980 558152
rect 137848 557506 137968 557534
rect 137756 554390 137876 554418
rect 137480 552894 137784 552922
rect 137756 552022 137784 552894
rect 137744 552016 137796 552022
rect 137744 551958 137796 551964
rect 137848 551410 137876 554390
rect 137836 551404 137888 551410
rect 137836 551346 137888 551352
rect 137284 550588 137336 550594
rect 137284 550530 137336 550536
rect 137112 550446 137692 550474
rect 137664 547963 137692 550446
rect 137940 550186 137968 557506
rect 139032 552832 139084 552838
rect 139032 552774 139084 552780
rect 138296 550248 138348 550254
rect 138296 550190 138348 550196
rect 137928 550180 137980 550186
rect 137928 550122 137980 550128
rect 138308 547963 138336 550190
rect 139044 547963 139072 552774
rect 139320 549914 139348 622367
rect 139768 569900 139820 569906
rect 139768 569842 139820 569848
rect 139400 562352 139452 562358
rect 139400 562294 139452 562300
rect 139412 551342 139440 562294
rect 139780 557534 139808 569842
rect 139872 566098 139900 630362
rect 145024 568262 145222 568290
rect 159836 568262 160034 568290
rect 164332 568268 164384 568274
rect 140070 568126 140176 568154
rect 140148 567194 140176 568126
rect 142356 568126 142646 568154
rect 142160 567656 142212 567662
rect 142160 567598 142212 567604
rect 139964 567166 140176 567194
rect 139860 566092 139912 566098
rect 139860 566034 139912 566040
rect 139964 562358 139992 567166
rect 140780 566296 140832 566302
rect 140780 566238 140832 566244
rect 139952 562352 140004 562358
rect 139952 562294 140004 562300
rect 139780 557506 139900 557534
rect 139768 552016 139820 552022
rect 139768 551958 139820 551964
rect 139400 551336 139452 551342
rect 139400 551278 139452 551284
rect 139308 549908 139360 549914
rect 139308 549850 139360 549856
rect 139780 547963 139808 551958
rect 139872 550458 139900 557506
rect 140504 556844 140556 556850
rect 140504 556786 140556 556792
rect 139860 550452 139912 550458
rect 139860 550394 139912 550400
rect 140516 547963 140544 556786
rect 140792 552786 140820 566238
rect 140872 566092 140924 566098
rect 140872 566034 140924 566040
rect 140884 557534 140912 566034
rect 140884 557506 141924 557534
rect 140792 552758 141280 552786
rect 141252 547963 141280 552758
rect 141896 547963 141924 557506
rect 142172 552770 142200 567598
rect 142252 561060 142304 561066
rect 142252 561002 142304 561008
rect 142264 552786 142292 561002
rect 142356 555626 142384 568126
rect 145024 567194 145052 568262
rect 145288 568200 145340 568206
rect 145288 568142 145340 568148
rect 145024 567166 145144 567194
rect 143540 565548 143592 565554
rect 143540 565490 143592 565496
rect 142344 555620 142396 555626
rect 142344 555562 142396 555568
rect 142160 552764 142212 552770
rect 142264 552758 142660 552786
rect 143552 552770 143580 565490
rect 145116 565282 145144 567166
rect 145104 565276 145156 565282
rect 145104 565218 145156 565224
rect 145300 557534 145328 568142
rect 148442 568126 148824 568154
rect 148796 565622 148824 568126
rect 150624 568132 150676 568138
rect 151018 568126 151400 568154
rect 150624 568074 150676 568080
rect 148784 565616 148836 565622
rect 148784 565558 148836 565564
rect 147772 565480 147824 565486
rect 147772 565422 147824 565428
rect 147680 565276 147732 565282
rect 147680 565218 147732 565224
rect 145300 557506 145512 557534
rect 144092 555552 144144 555558
rect 144092 555494 144144 555500
rect 142160 552706 142212 552712
rect 142632 547963 142660 552758
rect 143356 552764 143408 552770
rect 143356 552706 143408 552712
rect 143540 552764 143592 552770
rect 143540 552706 143592 552712
rect 143368 547963 143396 552706
rect 144104 547963 144132 555494
rect 144736 552764 144788 552770
rect 144736 552706 144788 552712
rect 144748 547963 144776 552706
rect 145484 547963 145512 557506
rect 146944 550520 146996 550526
rect 146944 550462 146996 550468
rect 146208 549976 146260 549982
rect 146208 549918 146260 549924
rect 146220 547963 146248 549918
rect 146956 547963 146984 550462
rect 147692 547963 147720 565218
rect 147784 557534 147812 565422
rect 149152 558204 149204 558210
rect 149152 558146 149204 558152
rect 149164 557534 149192 558146
rect 147784 557506 148364 557534
rect 149164 557506 149836 557534
rect 148336 547963 148364 557506
rect 149060 551404 149112 551410
rect 149060 551346 149112 551352
rect 149072 547963 149100 551346
rect 149808 547963 149836 557506
rect 150636 548162 150664 568074
rect 151372 565690 151400 568126
rect 153856 568126 154238 568154
rect 154580 568132 154632 568138
rect 151820 568064 151872 568070
rect 151820 568006 151872 568012
rect 151360 565684 151412 565690
rect 151360 565626 151412 565632
rect 151832 557534 151860 568006
rect 153856 565350 153884 568126
rect 154580 568074 154632 568080
rect 156432 568126 156814 568154
rect 153844 565344 153896 565350
rect 153844 565286 153896 565292
rect 151832 557506 151952 557534
rect 151268 550384 151320 550390
rect 151268 550326 151320 550332
rect 150560 548134 150664 548162
rect 150560 547944 150588 548134
rect 151280 547963 151308 550326
rect 151924 547963 151952 557506
rect 152648 556912 152700 556918
rect 152648 556854 152700 556860
rect 152660 547963 152688 556854
rect 154592 552770 154620 568074
rect 156052 568064 156104 568070
rect 156052 568006 156104 568012
rect 154672 565412 154724 565418
rect 154672 565354 154724 565360
rect 154684 557534 154712 565354
rect 156064 557534 156092 568006
rect 156432 565554 156460 568126
rect 158720 567928 158772 567934
rect 158720 567870 158772 567876
rect 157984 566840 158036 566846
rect 157984 566782 158036 566788
rect 156420 565548 156472 565554
rect 156420 565490 156472 565496
rect 154684 557506 154896 557534
rect 156064 557506 156276 557534
rect 154580 552764 154632 552770
rect 154580 552706 154632 552712
rect 154120 550588 154172 550594
rect 154120 550530 154172 550536
rect 153384 550452 153436 550458
rect 153384 550394 153436 550400
rect 153396 547963 153424 550394
rect 154132 547963 154160 550530
rect 154868 547963 154896 557506
rect 155500 552764 155552 552770
rect 155500 552706 155552 552712
rect 155512 547963 155540 552706
rect 156248 547963 156276 557506
rect 157248 554192 157300 554198
rect 157248 554134 157300 554140
rect 157260 550594 157288 554134
rect 157248 550588 157300 550594
rect 157248 550530 157300 550536
rect 157708 550316 157760 550322
rect 157708 550258 157760 550264
rect 156972 550180 157024 550186
rect 156972 550122 157024 550128
rect 156984 547963 157012 550122
rect 157720 547963 157748 550258
rect 157996 550254 158024 566782
rect 158732 552786 158760 567870
rect 159836 567194 159864 568262
rect 164332 568210 164384 568216
rect 162320 568126 162610 568154
rect 161664 567860 161716 567866
rect 161664 567802 161716 567808
rect 159836 567166 159956 567194
rect 159364 565616 159416 565622
rect 159364 565558 159416 565564
rect 158812 565344 158864 565350
rect 158812 565286 158864 565292
rect 158824 557534 158852 565286
rect 158824 557506 159220 557534
rect 158732 552758 159128 552786
rect 157984 550248 158036 550254
rect 157984 550190 158036 550196
rect 158352 550180 158404 550186
rect 158352 550122 158404 550128
rect 158364 547963 158392 550122
rect 159100 547963 159128 552758
rect 159192 550202 159220 557506
rect 159376 550390 159404 565558
rect 159928 565554 159956 567166
rect 160100 566500 160152 566506
rect 160100 566442 160152 566448
rect 159916 565548 159968 565554
rect 159916 565490 159968 565496
rect 160112 552770 160140 566442
rect 160744 565684 160796 565690
rect 160744 565626 160796 565632
rect 160192 563712 160244 563718
rect 160192 563654 160244 563660
rect 160204 557534 160232 563654
rect 160204 557506 160600 557534
rect 160100 552764 160152 552770
rect 160100 552706 160152 552712
rect 159364 550384 159416 550390
rect 159364 550326 159416 550332
rect 159192 550174 159864 550202
rect 159836 547963 159864 550174
rect 160572 547963 160600 557506
rect 160756 550254 160784 565626
rect 161676 557534 161704 567802
rect 162320 565486 162348 568126
rect 162308 565480 162360 565486
rect 162308 565422 162360 565428
rect 161676 557506 161980 557534
rect 161296 552764 161348 552770
rect 161296 552706 161348 552712
rect 160744 550248 160796 550254
rect 160744 550190 160796 550196
rect 161308 547963 161336 552706
rect 161952 547963 161980 557506
rect 164344 552770 164372 568210
rect 182364 568200 182416 568206
rect 165632 568126 165830 568154
rect 168406 568126 168512 568154
rect 164884 565548 164936 565554
rect 164884 565490 164936 565496
rect 164332 552764 164384 552770
rect 164332 552706 164384 552712
rect 163412 551336 163464 551342
rect 163412 551278 163464 551284
rect 162676 550520 162728 550526
rect 162676 550462 162728 550468
rect 162688 547963 162716 550462
rect 163424 547963 163452 551278
rect 164896 550458 164924 565490
rect 165528 552764 165580 552770
rect 165528 552706 165580 552712
rect 164884 550452 164936 550458
rect 164884 550394 164936 550400
rect 164148 550316 164200 550322
rect 164148 550258 164200 550264
rect 164160 547963 164188 550258
rect 164884 550112 164936 550118
rect 164884 550054 164936 550060
rect 164896 547963 164924 550054
rect 165540 547963 165568 552706
rect 165632 550594 165660 568126
rect 168484 567194 168512 568126
rect 168392 567166 168512 567194
rect 171336 568126 171626 568154
rect 174004 568126 174202 568154
rect 177040 568126 177422 568154
rect 179524 568126 179998 568154
rect 182364 568142 182416 568148
rect 165712 560992 165764 560998
rect 165712 560934 165764 560940
rect 165724 557534 165752 560934
rect 165724 557506 166304 557534
rect 165620 550588 165672 550594
rect 165620 550530 165672 550536
rect 166276 547963 166304 557506
rect 167736 555620 167788 555626
rect 167736 555562 167788 555568
rect 167000 550384 167052 550390
rect 167000 550326 167052 550332
rect 167012 547963 167040 550326
rect 167748 547963 167776 555562
rect 168392 551562 168420 567166
rect 171336 565418 171364 568126
rect 171324 565412 171376 565418
rect 171324 565354 171376 565360
rect 174004 564466 174032 568126
rect 177040 565146 177068 568126
rect 179420 567860 179472 567866
rect 179420 567802 179472 567808
rect 177028 565140 177080 565146
rect 177028 565082 177080 565088
rect 173164 564460 173216 564466
rect 173164 564402 173216 564408
rect 173992 564460 174044 564466
rect 173992 564402 174044 564408
rect 168472 559564 168524 559570
rect 168472 559506 168524 559512
rect 168484 557534 168512 559506
rect 168484 557506 169156 557534
rect 168392 551534 168512 551562
rect 168380 551404 168432 551410
rect 168380 551346 168432 551352
rect 168392 547963 168420 551346
rect 168484 550526 168512 551534
rect 168472 550520 168524 550526
rect 168472 550462 168524 550468
rect 169128 547963 169156 557506
rect 171324 551472 171376 551478
rect 171324 551414 171376 551420
rect 169852 550588 169904 550594
rect 169852 550530 169904 550536
rect 169864 547963 169892 550530
rect 170588 550112 170640 550118
rect 170588 550054 170640 550060
rect 170600 547963 170628 550054
rect 171336 547963 171364 551414
rect 173176 550322 173204 564402
rect 173900 562352 173952 562358
rect 173900 562294 173952 562300
rect 173912 557534 173940 562294
rect 176660 559768 176712 559774
rect 176660 559710 176712 559716
rect 173912 557506 174952 557534
rect 174176 550588 174228 550594
rect 174176 550530 174228 550536
rect 173440 550452 173492 550458
rect 173440 550394 173492 550400
rect 173164 550316 173216 550322
rect 173164 550258 173216 550264
rect 172704 550248 172756 550254
rect 172704 550190 172756 550196
rect 171968 550044 172020 550050
rect 171968 549986 172020 549992
rect 171980 547963 172008 549986
rect 172716 547963 172744 550190
rect 173452 547963 173480 550394
rect 174188 547963 174216 550530
rect 174924 547963 174952 557506
rect 176672 552786 176700 559710
rect 176752 558408 176804 558414
rect 176752 558350 176804 558356
rect 176764 557534 176792 558350
rect 176764 557506 177804 557534
rect 176672 552758 177068 552786
rect 176292 550044 176344 550050
rect 176292 549986 176344 549992
rect 175556 549908 175608 549914
rect 175556 549850 175608 549856
rect 175568 547963 175596 549850
rect 176304 547963 176332 549986
rect 177040 547963 177068 552758
rect 177776 547963 177804 557506
rect 178500 555620 178552 555626
rect 178500 555562 178552 555568
rect 178512 547963 178540 555562
rect 179144 554056 179196 554062
rect 179144 553998 179196 554004
rect 179156 547963 179184 553998
rect 179432 550474 179460 567802
rect 179524 550594 179552 568126
rect 180892 566568 180944 566574
rect 180892 566510 180944 566516
rect 180800 566500 180852 566506
rect 180800 566442 180852 566448
rect 179604 563712 179656 563718
rect 179604 563654 179656 563660
rect 179616 557534 179644 563654
rect 179616 557506 180656 557534
rect 179512 550588 179564 550594
rect 179512 550530 179564 550536
rect 179432 550446 179920 550474
rect 179892 547963 179920 550446
rect 180628 547963 180656 557506
rect 180812 552770 180840 566442
rect 180904 557534 180932 566510
rect 180904 557506 181392 557534
rect 180800 552764 180852 552770
rect 180800 552706 180852 552712
rect 181364 547963 181392 557506
rect 181996 552764 182048 552770
rect 181996 552706 182048 552712
rect 182008 547963 182036 552706
rect 182376 550066 182404 568142
rect 182928 568126 183218 568154
rect 185504 568126 185794 568154
rect 187896 568126 189014 568154
rect 191208 568126 191590 568154
rect 194810 568126 194916 568154
rect 197386 568126 197492 568154
rect 182824 565412 182876 565418
rect 182824 565354 182876 565360
rect 182836 550186 182864 565354
rect 182928 565350 182956 568126
rect 182916 565344 182968 565350
rect 182916 565286 182968 565292
rect 185504 565282 185532 568126
rect 187792 566636 187844 566642
rect 187792 566578 187844 566584
rect 185492 565276 185544 565282
rect 185492 565218 185544 565224
rect 187700 564936 187752 564942
rect 187700 564878 187752 564884
rect 187712 562562 187740 564878
rect 187700 562556 187752 562562
rect 187700 562498 187752 562504
rect 184940 562420 184992 562426
rect 184940 562362 184992 562368
rect 184952 557534 184980 562362
rect 186320 562352 186372 562358
rect 186320 562294 186372 562300
rect 184952 557506 185624 557534
rect 184940 552900 184992 552906
rect 184940 552842 184992 552848
rect 184204 551336 184256 551342
rect 184204 551278 184256 551284
rect 182824 550180 182876 550186
rect 182824 550122 182876 550128
rect 182376 550038 183508 550066
rect 182732 549908 182784 549914
rect 182732 549850 182784 549856
rect 182744 547963 182772 549850
rect 183480 547963 183508 550038
rect 184216 547963 184244 551278
rect 184952 547963 184980 552842
rect 185596 547963 185624 557506
rect 186332 547963 186360 562294
rect 186412 558204 186464 558210
rect 186412 558146 186464 558152
rect 186424 557534 186452 558146
rect 186424 557506 187096 557534
rect 187068 547963 187096 557506
rect 187804 547963 187832 566578
rect 187896 558346 187924 568126
rect 190644 565276 190696 565282
rect 190644 565218 190696 565224
rect 190552 561196 190604 561202
rect 190552 561138 190604 561144
rect 187884 558340 187936 558346
rect 187884 558282 187936 558288
rect 188528 556980 188580 556986
rect 188528 556922 188580 556928
rect 188540 547963 188568 556922
rect 189908 554260 189960 554266
rect 189908 554202 189960 554208
rect 189172 552764 189224 552770
rect 189172 552706 189224 552712
rect 189184 547963 189212 552706
rect 189920 547963 189948 554202
rect 190564 552786 190592 561138
rect 190656 557534 190684 565218
rect 191208 564942 191236 568126
rect 194600 567928 194652 567934
rect 194600 567870 194652 567876
rect 191840 565140 191892 565146
rect 191840 565082 191892 565088
rect 191196 564936 191248 564942
rect 191196 564878 191248 564884
rect 191852 557534 191880 565082
rect 193220 561128 193272 561134
rect 193220 561070 193272 561076
rect 193232 557534 193260 561070
rect 190656 557506 191420 557534
rect 191852 557506 192800 557534
rect 193232 557506 194272 557534
rect 190564 552758 190684 552786
rect 190656 547963 190684 552758
rect 191392 547963 191420 557506
rect 192116 557048 192168 557054
rect 192116 556990 192168 556996
rect 192128 547963 192156 556990
rect 192772 547963 192800 557506
rect 193496 555688 193548 555694
rect 193496 555630 193548 555636
rect 193508 547963 193536 555630
rect 194244 547963 194272 557506
rect 194612 552514 194640 567870
rect 194888 567194 194916 568126
rect 194704 567166 194916 567194
rect 194704 552702 194732 567166
rect 197464 565214 197492 568126
rect 200224 568126 200606 568154
rect 197452 565208 197504 565214
rect 197452 565150 197504 565156
rect 200224 564466 200252 568126
rect 200304 566704 200356 566710
rect 200304 566646 200356 566652
rect 198004 564460 198056 564466
rect 198004 564402 198056 564408
rect 200212 564460 200264 564466
rect 200212 564402 200264 564408
rect 195980 563780 196032 563786
rect 195980 563722 196032 563728
rect 195992 552786 196020 563722
rect 196072 559564 196124 559570
rect 196072 559506 196124 559512
rect 196084 557534 196112 559506
rect 197360 558340 197412 558346
rect 197360 558282 197412 558288
rect 197372 557534 197400 558282
rect 196084 557506 197124 557534
rect 197372 557506 197860 557534
rect 195992 552758 196388 552786
rect 194692 552696 194744 552702
rect 194692 552638 194744 552644
rect 194612 552486 195008 552514
rect 194980 547963 195008 552486
rect 195612 550180 195664 550186
rect 195612 550122 195664 550128
rect 195624 547963 195652 550122
rect 196360 547963 196388 552758
rect 197096 547963 197124 557506
rect 197832 547963 197860 557506
rect 198016 556850 198044 564402
rect 198740 562556 198792 562562
rect 198740 562498 198792 562504
rect 198752 557534 198780 562498
rect 198752 557506 199240 557534
rect 198004 556844 198056 556850
rect 198004 556786 198056 556792
rect 198556 552696 198608 552702
rect 198556 552638 198608 552644
rect 198568 547963 198596 552638
rect 199212 547963 199240 557506
rect 200316 552786 200344 566646
rect 200684 557534 200712 630414
rect 200762 618488 200818 618497
rect 200762 618423 200818 618432
rect 200776 566778 200804 618423
rect 200868 568274 200896 633422
rect 201592 630420 201644 630426
rect 201592 630362 201644 630368
rect 201038 594620 201094 594629
rect 201038 594555 201094 594564
rect 200948 569900 201000 569906
rect 200948 569842 201000 569848
rect 200856 568268 200908 568274
rect 200856 568210 200908 568216
rect 200764 566772 200816 566778
rect 200764 566714 200816 566720
rect 200684 557506 200804 557534
rect 200316 552758 200712 552786
rect 199936 550316 199988 550322
rect 199936 550258 199988 550264
rect 199948 547963 199976 550258
rect 200684 547963 200712 552758
rect 200776 551410 200804 557506
rect 200764 551404 200816 551410
rect 200764 551346 200816 551352
rect 200960 550118 200988 569842
rect 201052 563854 201080 594555
rect 201498 584488 201554 584497
rect 201498 584423 201554 584432
rect 201130 576260 201186 576269
rect 201130 576195 201186 576204
rect 201040 563848 201092 563854
rect 201040 563790 201092 563796
rect 201144 555490 201172 576195
rect 201222 570140 201278 570149
rect 201222 570075 201278 570084
rect 201236 558278 201264 570075
rect 201512 562494 201540 584423
rect 201500 562488 201552 562494
rect 201500 562430 201552 562436
rect 201500 560992 201552 560998
rect 201500 560934 201552 560940
rect 201224 558272 201276 558278
rect 201224 558214 201276 558220
rect 201132 555484 201184 555490
rect 201132 555426 201184 555432
rect 201408 550588 201460 550594
rect 201408 550530 201460 550536
rect 200948 550112 201000 550118
rect 200948 550054 201000 550060
rect 201420 547963 201448 550530
rect 201512 549794 201540 560934
rect 201604 549982 201632 630362
rect 201696 568138 201724 633490
rect 204260 632732 204312 632738
rect 204260 632674 204312 632680
rect 201774 628008 201830 628017
rect 201774 627943 201830 627952
rect 201684 568132 201736 568138
rect 201684 568074 201736 568080
rect 201788 568002 201816 627943
rect 202970 625288 203026 625297
rect 202970 625223 203026 625232
rect 202234 621208 202290 621217
rect 202234 621143 202290 621152
rect 201866 612776 201922 612785
rect 201866 612711 201922 612720
rect 201776 567996 201828 568002
rect 201776 567938 201828 567944
rect 201880 559638 201908 612711
rect 201958 608968 202014 608977
rect 201958 608903 202014 608912
rect 201972 563922 202000 608903
rect 202050 600400 202106 600409
rect 202050 600335 202106 600344
rect 201960 563916 202012 563922
rect 201960 563858 202012 563864
rect 201868 559632 201920 559638
rect 201868 559574 201920 559580
rect 202064 556918 202092 600335
rect 202142 590744 202198 590753
rect 202142 590679 202198 590688
rect 202052 556912 202104 556918
rect 202052 556854 202104 556860
rect 202156 552906 202184 590679
rect 202248 555558 202276 621143
rect 202878 615632 202934 615641
rect 202878 615567 202934 615576
rect 202326 578368 202382 578377
rect 202326 578303 202382 578312
rect 202236 555552 202288 555558
rect 202236 555494 202288 555500
rect 202340 554130 202368 578303
rect 202892 559706 202920 615567
rect 202984 569906 203012 625223
rect 203154 606384 203210 606393
rect 203154 606319 203210 606328
rect 203062 603120 203118 603129
rect 203062 603055 203118 603064
rect 202972 569900 203024 569906
rect 202972 569842 203024 569848
rect 202880 559700 202932 559706
rect 202880 559642 202932 559648
rect 203076 554198 203104 603055
rect 203168 566846 203196 606319
rect 203246 596728 203302 596737
rect 203246 596663 203248 596672
rect 203300 596663 203302 596672
rect 203248 596634 203300 596640
rect 203246 588024 203302 588033
rect 203246 587959 203302 587968
rect 203156 566840 203208 566846
rect 203156 566782 203208 566788
rect 203260 561066 203288 587959
rect 203338 581768 203394 581777
rect 203338 581703 203394 581712
rect 203352 565350 203380 581703
rect 203430 572792 203486 572801
rect 203430 572727 203486 572736
rect 203340 565344 203392 565350
rect 203340 565286 203392 565292
rect 203248 561060 203300 561066
rect 203248 561002 203300 561008
rect 203064 554192 203116 554198
rect 203064 554134 203116 554140
rect 202328 554124 202380 554130
rect 202328 554066 202380 554072
rect 202144 552900 202196 552906
rect 202144 552842 202196 552848
rect 203444 551478 203472 572727
rect 203432 551472 203484 551478
rect 203432 551414 203484 551420
rect 202788 550520 202840 550526
rect 202788 550462 202840 550468
rect 201592 549976 201644 549982
rect 201592 549918 201644 549924
rect 201512 549766 202184 549794
rect 202156 547963 202184 549766
rect 202800 547963 202828 550462
rect 203524 549364 203576 549370
rect 203524 549306 203576 549312
rect 203536 547963 203564 549306
rect 204272 547963 204300 632674
rect 204352 631032 204404 631038
rect 204352 630974 204404 630980
rect 204364 552786 204392 630974
rect 204456 568070 204484 633626
rect 208400 632256 208452 632262
rect 208400 632198 208452 632204
rect 206284 632188 206336 632194
rect 206284 632130 206336 632136
rect 204904 630964 204956 630970
rect 204904 630906 204956 630912
rect 204536 596692 204588 596698
rect 204536 596634 204588 596640
rect 204548 568478 204576 596634
rect 204536 568472 204588 568478
rect 204536 568414 204588 568420
rect 204444 568064 204496 568070
rect 204444 568006 204496 568012
rect 204916 557534 204944 630906
rect 204996 615528 205048 615534
rect 204996 615470 205048 615476
rect 205008 561202 205036 615470
rect 204996 561196 205048 561202
rect 204996 561138 205048 561144
rect 204916 557506 205128 557534
rect 204364 552758 205036 552786
rect 205008 547963 205036 552758
rect 205100 550322 205128 557506
rect 205640 555484 205692 555490
rect 205640 555426 205692 555432
rect 205088 550316 205140 550322
rect 205088 550258 205140 550264
rect 205652 547963 205680 555426
rect 206296 550594 206324 632130
rect 206376 630896 206428 630902
rect 206376 630838 206428 630844
rect 206388 557534 206416 630838
rect 206468 619676 206520 619682
rect 206468 619618 206520 619624
rect 206480 562562 206508 619618
rect 206560 582412 206612 582418
rect 206560 582354 206612 582360
rect 206468 562556 206520 562562
rect 206468 562498 206520 562504
rect 206388 557506 206508 557534
rect 206376 554124 206428 554130
rect 206376 554066 206428 554072
rect 206284 550588 206336 550594
rect 206284 550530 206336 550536
rect 206388 547963 206416 554066
rect 206480 550186 206508 557506
rect 206572 555626 206600 582354
rect 207020 570648 207072 570654
rect 207020 570590 207072 570596
rect 207032 557534 207060 570590
rect 207032 557506 207888 557534
rect 206560 555620 206612 555626
rect 206560 555562 206612 555568
rect 207112 551132 207164 551138
rect 207112 551074 207164 551080
rect 206468 550180 206520 550186
rect 206468 550122 206520 550128
rect 207124 547963 207152 551074
rect 207860 547963 207888 557506
rect 208412 552838 208440 632198
rect 208492 625184 208544 625190
rect 208492 625126 208544 625132
rect 208504 557534 208532 625126
rect 209044 579692 209096 579698
rect 209044 579634 209096 579640
rect 209056 558346 209084 579634
rect 209044 558340 209096 558346
rect 209044 558282 209096 558288
rect 209792 557534 209820 633626
rect 208504 557506 208624 557534
rect 209792 557506 210004 557534
rect 208492 555552 208544 555558
rect 208492 555494 208544 555500
rect 208400 552832 208452 552838
rect 208400 552774 208452 552780
rect 208504 550526 208532 555494
rect 208492 550520 208544 550526
rect 208492 550462 208544 550468
rect 208596 547963 208624 557506
rect 209228 552832 209280 552838
rect 209228 552774 209280 552780
rect 209240 547963 209268 552774
rect 209976 547963 210004 557506
rect 210436 557054 210464 634034
rect 213920 634024 213972 634030
rect 213920 633966 213972 633972
rect 212540 633956 212592 633962
rect 212540 633898 212592 633904
rect 211804 630760 211856 630766
rect 211804 630702 211856 630708
rect 211160 594856 211212 594862
rect 211160 594798 211212 594804
rect 210516 590708 210568 590714
rect 210516 590650 210568 590656
rect 210424 557048 210476 557054
rect 210424 556990 210476 556996
rect 210528 551138 210556 590650
rect 211172 557534 211200 594798
rect 211172 557506 211476 557534
rect 210700 552900 210752 552906
rect 210700 552842 210752 552848
rect 210516 551132 210568 551138
rect 210516 551074 210568 551080
rect 210712 547963 210740 552842
rect 211448 547963 211476 557506
rect 211816 549370 211844 630702
rect 212552 552838 212580 633898
rect 213184 630828 213236 630834
rect 213184 630770 213236 630776
rect 212632 565344 212684 565350
rect 212632 565286 212684 565292
rect 212644 557534 212672 565286
rect 212644 557506 212856 557534
rect 212540 552832 212592 552838
rect 212540 552774 212592 552780
rect 212172 550112 212224 550118
rect 212172 550054 212224 550060
rect 211804 549364 211856 549370
rect 211804 549306 211856 549312
rect 212184 547963 212212 550054
rect 212828 547963 212856 557506
rect 213196 550050 213224 630770
rect 213276 597576 213328 597582
rect 213276 597518 213328 597524
rect 213288 559774 213316 597518
rect 213276 559768 213328 559774
rect 213276 559710 213328 559716
rect 213932 552838 213960 633966
rect 217876 633888 217928 633894
rect 217876 633830 217928 633836
rect 214012 633616 214064 633622
rect 214012 633558 214064 633564
rect 214024 557534 214052 633558
rect 217324 633480 217376 633486
rect 217324 633422 217376 633428
rect 215300 632324 215352 632330
rect 215300 632266 215352 632272
rect 214024 557506 214328 557534
rect 213552 552832 213604 552838
rect 213552 552774 213604 552780
rect 213920 552832 213972 552838
rect 213920 552774 213972 552780
rect 213184 550044 213236 550050
rect 213184 549986 213236 549992
rect 213564 547963 213592 552774
rect 214300 547963 214328 557506
rect 215024 552832 215076 552838
rect 215024 552774 215076 552780
rect 215312 552786 215340 632266
rect 215942 628688 215998 628697
rect 215942 628623 215998 628632
rect 215392 562556 215444 562562
rect 215392 562498 215444 562504
rect 215404 557534 215432 562498
rect 215404 557506 215892 557534
rect 215864 552786 215892 557506
rect 215956 555694 215984 628623
rect 216678 625832 216734 625841
rect 216678 625767 216734 625776
rect 216692 625190 216720 625767
rect 216680 625184 216732 625190
rect 216680 625126 216732 625132
rect 216678 619712 216734 619721
rect 216678 619647 216680 619656
rect 216732 619647 216734 619656
rect 216680 619618 216732 619624
rect 216678 616312 216734 616321
rect 216678 616247 216734 616256
rect 216692 615534 216720 616247
rect 216680 615528 216732 615534
rect 216680 615470 216732 615476
rect 216678 597952 216734 597961
rect 216678 597887 216734 597896
rect 216692 597582 216720 597887
rect 216680 597576 216732 597582
rect 216680 597518 216732 597524
rect 216678 595232 216734 595241
rect 216678 595167 216734 595176
rect 216692 594862 216720 595167
rect 216680 594856 216732 594862
rect 216680 594798 216732 594804
rect 216678 591832 216734 591841
rect 216678 591767 216734 591776
rect 216692 590714 216720 591767
rect 216680 590708 216732 590714
rect 216680 590650 216732 590656
rect 216034 585712 216090 585721
rect 216034 585647 216090 585656
rect 215944 555688 215996 555694
rect 215944 555630 215996 555636
rect 216048 552974 216076 585647
rect 216678 582992 216734 583001
rect 216678 582927 216734 582936
rect 216692 582418 216720 582927
rect 216680 582412 216732 582418
rect 216680 582354 216732 582360
rect 216678 579728 216734 579737
rect 216678 579663 216680 579672
rect 216732 579663 216734 579672
rect 216680 579634 216732 579640
rect 216678 570752 216734 570761
rect 216678 570687 216734 570696
rect 216692 557534 216720 570687
rect 216692 557506 217180 557534
rect 216036 552968 216088 552974
rect 216036 552910 216088 552916
rect 215036 547963 215064 552774
rect 215312 552758 215800 552786
rect 215864 552758 216444 552786
rect 215772 547963 215800 552758
rect 216416 547963 216444 552758
rect 217152 547963 217180 557506
rect 217336 554266 217364 633422
rect 217690 622432 217746 622441
rect 217690 622367 217746 622376
rect 217414 601352 217470 601361
rect 217414 601287 217470 601296
rect 217428 570654 217456 601287
rect 217598 589112 217654 589121
rect 217598 589047 217654 589056
rect 217506 573472 217562 573481
rect 217506 573407 217562 573416
rect 217416 570648 217468 570654
rect 217416 570590 217468 570596
rect 217324 554260 217376 554266
rect 217324 554202 217376 554208
rect 217520 550594 217548 573407
rect 217612 561066 217640 589047
rect 217704 568614 217732 622367
rect 217782 610192 217838 610201
rect 217782 610127 217838 610136
rect 217692 568608 217744 568614
rect 217692 568550 217744 568556
rect 217600 561060 217652 561066
rect 217600 561002 217652 561008
rect 217796 556238 217824 610127
rect 217888 568002 217916 633830
rect 217968 631100 218020 631106
rect 217968 631042 218020 631048
rect 217876 567996 217928 568002
rect 217876 567938 217928 567944
rect 217784 556232 217836 556238
rect 217784 556174 217836 556180
rect 217876 555688 217928 555694
rect 217876 555630 217928 555636
rect 217508 550588 217560 550594
rect 217508 550530 217560 550536
rect 217888 547963 217916 555630
rect 217980 550050 218008 631042
rect 218716 630698 218744 638930
rect 218888 633820 218940 633826
rect 218888 633762 218940 633768
rect 218796 633752 218848 633758
rect 218796 633694 218848 633700
rect 218704 630692 218756 630698
rect 218704 630634 218756 630640
rect 218716 604217 218744 630634
rect 218702 604208 218758 604217
rect 218702 604143 218758 604152
rect 218808 561134 218836 633694
rect 218900 568206 218928 633762
rect 219176 607617 219204 639066
rect 219716 634092 219768 634098
rect 219716 634034 219768 634040
rect 219348 633548 219400 633554
rect 219348 633490 219400 633496
rect 219254 613592 219310 613601
rect 219254 613527 219310 613536
rect 219162 607608 219218 607617
rect 219162 607543 219218 607552
rect 219162 576872 219218 576881
rect 219162 576807 219218 576816
rect 218888 568200 218940 568206
rect 218888 568142 218940 568148
rect 218796 561128 218848 561134
rect 218796 561070 218848 561076
rect 218612 556232 218664 556238
rect 218612 556174 218664 556180
rect 217968 550044 218020 550050
rect 217968 549986 218020 549992
rect 218624 547963 218652 556174
rect 219176 551410 219204 576807
rect 219268 563854 219296 613527
rect 219360 568070 219388 633490
rect 219728 630986 219756 634034
rect 225420 634024 225472 634030
rect 225420 633966 225472 633972
rect 222844 631032 222896 631038
rect 219728 630958 220018 630986
rect 225432 630986 225460 633966
rect 271880 633956 271932 633962
rect 271880 633898 271932 633904
rect 242900 633888 242952 633894
rect 242900 633830 242952 633836
rect 231308 633480 231360 633486
rect 231308 633422 231360 633428
rect 228732 631100 228784 631106
rect 228732 631042 228784 631048
rect 228744 630986 228772 631042
rect 231320 630986 231348 633422
rect 234620 632324 234672 632330
rect 234620 632266 234672 632272
rect 234632 630986 234660 632266
rect 240324 632256 240376 632262
rect 240324 632198 240376 632204
rect 240336 630986 240364 632198
rect 242912 630986 242940 633830
rect 251916 633820 251968 633826
rect 251916 633762 251968 633768
rect 251928 630986 251956 633762
rect 263600 633752 263652 633758
rect 263600 633694 263652 633700
rect 260196 633684 260248 633690
rect 260196 633626 260248 633632
rect 254492 632188 254544 632194
rect 254492 632130 254544 632136
rect 254504 630986 254532 632130
rect 260208 630986 260236 633626
rect 263612 630986 263640 633694
rect 269212 633616 269264 633622
rect 269212 633558 269264 633564
rect 269224 630986 269252 633558
rect 270408 633480 270460 633486
rect 270408 633422 270460 633428
rect 270420 632738 270448 633422
rect 270408 632732 270460 632738
rect 270408 632674 270460 632680
rect 271892 630986 271920 633898
rect 275100 633548 275152 633554
rect 275100 633490 275152 633496
rect 275112 630986 275140 633490
rect 277676 633480 277728 633486
rect 277676 633422 277728 633428
rect 277688 630986 277716 633422
rect 222896 630980 223238 630986
rect 222844 630974 223238 630980
rect 222856 630958 223238 630974
rect 225432 630958 225814 630986
rect 228744 630958 229034 630986
rect 231320 630958 231610 630986
rect 234632 630958 234830 630986
rect 237300 630970 237406 630986
rect 237288 630964 237406 630970
rect 237340 630958 237406 630964
rect 240336 630958 240626 630986
rect 242912 630958 243202 630986
rect 251928 630958 252218 630986
rect 254504 630958 254794 630986
rect 260208 630958 260590 630986
rect 263612 630958 263810 630986
rect 269224 630958 269606 630986
rect 271892 630958 272182 630986
rect 275112 630958 275402 630986
rect 277688 630958 277978 630986
rect 237288 630906 237340 630912
rect 248696 630896 248748 630902
rect 248748 630844 248998 630850
rect 248696 630838 248998 630844
rect 248708 630822 248998 630838
rect 257632 630834 258014 630850
rect 257620 630828 258014 630834
rect 257672 630822 258014 630828
rect 257620 630770 257672 630776
rect 266268 630760 266320 630766
rect 246040 630698 246422 630714
rect 266320 630708 266386 630714
rect 266268 630702 266386 630708
rect 219440 630692 219492 630698
rect 219440 630634 219492 630640
rect 246028 630692 246422 630698
rect 246080 630686 246422 630692
rect 266280 630686 266386 630702
rect 246028 630634 246080 630640
rect 219348 568064 219400 568070
rect 219348 568006 219400 568012
rect 219256 563848 219308 563854
rect 219256 563790 219308 563796
rect 219164 551404 219216 551410
rect 219164 551346 219216 551352
rect 219256 550588 219308 550594
rect 219256 550530 219308 550536
rect 219268 547963 219296 550530
rect 219452 550474 219480 630634
rect 280724 630562 280752 639610
rect 280712 630556 280764 630562
rect 280712 630498 280764 630504
rect 280554 630414 280844 630442
rect 280712 630352 280764 630358
rect 280712 630294 280764 630300
rect 219820 568670 220018 568698
rect 219820 568154 219848 568670
rect 219900 568608 219952 568614
rect 219900 568550 219952 568556
rect 219544 568126 219848 568154
rect 219544 550594 219572 568126
rect 219624 558476 219676 558482
rect 219624 558418 219676 558424
rect 219636 556102 219664 558418
rect 219912 557534 219940 568550
rect 222304 568126 222594 568154
rect 225064 568126 225170 568154
rect 228008 568126 228390 568154
rect 230492 568126 230966 568154
rect 233252 568126 234186 568154
rect 236012 568126 236762 568154
rect 238772 568126 239982 568154
rect 241532 568126 242558 568154
rect 245672 568126 245778 568154
rect 247144 568126 248354 568154
rect 251284 568126 251574 568154
rect 253952 568126 254150 568154
rect 257080 568126 257370 568154
rect 259656 568126 259946 568154
rect 262784 568126 263166 568154
rect 265360 568126 265742 568154
rect 268672 568126 268962 568154
rect 271248 568126 271538 568154
rect 274652 568126 274758 568154
rect 276952 568126 277334 568154
rect 280264 568126 280554 568154
rect 222200 567996 222252 568002
rect 222200 567938 222252 567944
rect 219912 557506 220124 557534
rect 219624 556096 219676 556102
rect 219624 556038 219676 556044
rect 219532 550588 219584 550594
rect 219532 550530 219584 550536
rect 219452 550446 220032 550474
rect 220004 547963 220032 550446
rect 220096 549982 220124 557506
rect 220728 556096 220780 556102
rect 220728 556038 220780 556044
rect 220084 549976 220136 549982
rect 220084 549918 220136 549924
rect 220740 547963 220768 556038
rect 222212 555830 222240 567938
rect 222200 555824 222252 555830
rect 222200 555766 222252 555772
rect 222304 550594 222332 568126
rect 223580 568064 223632 568070
rect 223580 568006 223632 568012
rect 222384 565412 222436 565418
rect 222384 565354 222436 565360
rect 221464 550588 221516 550594
rect 221464 550530 221516 550536
rect 222292 550588 222344 550594
rect 222292 550530 222344 550536
rect 221476 547963 221504 550530
rect 222396 548162 222424 565354
rect 222844 555824 222896 555830
rect 222844 555766 222896 555772
rect 222228 548134 222424 548162
rect 222228 547944 222256 548134
rect 222856 547963 222884 555766
rect 223592 547963 223620 568006
rect 223672 563848 223724 563854
rect 223672 563790 223724 563796
rect 223684 557534 223712 563790
rect 225064 558414 225092 568126
rect 227720 565208 227772 565214
rect 227720 565150 227772 565156
rect 225144 564460 225196 564466
rect 225144 564402 225196 564408
rect 225052 558408 225104 558414
rect 225052 558350 225104 558356
rect 223684 557506 224356 557534
rect 224328 547963 224356 557506
rect 225156 548162 225184 564402
rect 226432 563916 226484 563922
rect 226432 563858 226484 563864
rect 225788 550588 225840 550594
rect 225788 550530 225840 550536
rect 225080 548134 225184 548162
rect 225080 547944 225108 548134
rect 225800 547963 225828 550530
rect 226444 547963 226472 563858
rect 227732 552786 227760 565150
rect 228008 564466 228036 568126
rect 227996 564460 228048 564466
rect 227996 564402 228048 564408
rect 227812 558340 227864 558346
rect 227812 558282 227864 558288
rect 227824 557534 227852 558282
rect 230492 557534 230520 568126
rect 231860 565480 231912 565486
rect 231860 565422 231912 565428
rect 227824 557506 228680 557534
rect 230492 557506 230796 557534
rect 227732 552758 227944 552786
rect 227168 551404 227220 551410
rect 227168 551346 227220 551352
rect 227180 547963 227208 551346
rect 227916 547963 227944 552758
rect 228652 547963 228680 557506
rect 229284 556912 229336 556918
rect 229284 556854 229336 556860
rect 229296 547963 229324 556854
rect 230020 550044 230072 550050
rect 230020 549986 230072 549992
rect 230032 547963 230060 549986
rect 230768 547963 230796 557506
rect 231872 552786 231900 565422
rect 231952 561060 232004 561066
rect 231952 561002 232004 561008
rect 231964 557534 231992 561002
rect 231964 557506 232912 557534
rect 231872 552758 232268 552786
rect 231492 550044 231544 550050
rect 231492 549986 231544 549992
rect 231504 547963 231532 549986
rect 232240 547963 232268 552758
rect 232884 547963 232912 557506
rect 233252 556986 233280 568126
rect 234620 562488 234672 562494
rect 234620 562430 234672 562436
rect 233332 559632 233384 559638
rect 233332 559574 233384 559580
rect 233344 557534 233372 559574
rect 234632 557534 234660 562430
rect 233344 557506 234384 557534
rect 234632 557506 235120 557534
rect 233240 556980 233292 556986
rect 233240 556922 233292 556928
rect 233608 549976 233660 549982
rect 233608 549918 233660 549924
rect 233620 547963 233648 549918
rect 234356 547963 234384 557506
rect 235092 547963 235120 557506
rect 236012 555558 236040 568126
rect 236000 555552 236052 555558
rect 236000 555494 236052 555500
rect 236092 555552 236144 555558
rect 236092 555494 236144 555500
rect 236104 550118 236132 555494
rect 238668 552628 238720 552634
rect 238668 552570 238720 552576
rect 237932 552152 237984 552158
rect 237932 552094 237984 552100
rect 236092 550112 236144 550118
rect 236092 550054 236144 550060
rect 237196 549976 237248 549982
rect 237196 549918 237248 549924
rect 236460 548276 236512 548282
rect 236460 548218 236512 548224
rect 235816 548140 235868 548146
rect 235816 548082 235868 548088
rect 235828 547963 235856 548082
rect 236472 547963 236500 548218
rect 237208 547963 237236 549918
rect 237944 547963 237972 552094
rect 238680 547963 238708 552570
rect 238772 550050 238800 568126
rect 240140 559700 240192 559706
rect 240140 559642 240192 559648
rect 240152 557534 240180 559642
rect 240152 557506 240824 557534
rect 238760 550044 238812 550050
rect 238760 549986 238812 549992
rect 239404 550044 239456 550050
rect 239404 549986 239456 549992
rect 239416 547963 239444 549986
rect 240048 549500 240100 549506
rect 240048 549442 240100 549448
rect 240060 547963 240088 549442
rect 240796 547963 240824 557506
rect 241532 554130 241560 568126
rect 242164 568064 242216 568070
rect 242164 568006 242216 568012
rect 241520 554124 241572 554130
rect 241520 554066 241572 554072
rect 241518 550080 241574 550089
rect 241518 550015 241574 550024
rect 241532 547963 241560 550015
rect 242176 549914 242204 568006
rect 245672 565214 245700 568126
rect 245660 565208 245712 565214
rect 245660 565150 245712 565156
rect 247040 565208 247092 565214
rect 247040 565150 247092 565156
rect 245660 558272 245712 558278
rect 245660 558214 245712 558220
rect 245672 557534 245700 558214
rect 247052 557534 247080 565150
rect 247144 558482 247172 568126
rect 251284 565350 251312 568126
rect 253952 565418 253980 568126
rect 253940 565412 253992 565418
rect 253940 565354 253992 565360
rect 251272 565344 251324 565350
rect 251272 565286 251324 565292
rect 252560 565344 252612 565350
rect 252560 565286 252612 565292
rect 247132 558476 247184 558482
rect 247132 558418 247184 558424
rect 252572 557534 252600 565286
rect 257080 565282 257108 568126
rect 259656 565486 259684 568126
rect 260840 567996 260892 568002
rect 260840 567938 260892 567944
rect 259644 565480 259696 565486
rect 259644 565422 259696 565428
rect 257068 565276 257120 565282
rect 257068 565218 257120 565224
rect 260104 564460 260156 564466
rect 260104 564402 260156 564408
rect 255320 563848 255372 563854
rect 255320 563790 255372 563796
rect 245672 557506 246528 557534
rect 247052 557506 248000 557534
rect 252572 557506 253704 557534
rect 245108 556844 245160 556850
rect 245108 556786 245160 556792
rect 242900 554124 242952 554130
rect 242900 554066 242952 554072
rect 242256 552220 242308 552226
rect 242256 552162 242308 552168
rect 242164 549908 242216 549914
rect 242164 549850 242216 549856
rect 242268 547963 242296 552162
rect 242912 547963 242940 554066
rect 244372 551268 244424 551274
rect 244372 551210 244424 551216
rect 243636 549364 243688 549370
rect 243636 549306 243688 549312
rect 243648 547963 243676 549306
rect 244384 547963 244412 551210
rect 245120 547963 245148 556786
rect 245844 549908 245896 549914
rect 245844 549850 245896 549856
rect 245856 547963 245884 549850
rect 246500 547963 246528 557506
rect 247224 548140 247276 548146
rect 247224 548082 247276 548088
rect 247236 547963 247264 548082
rect 247972 547963 248000 557506
rect 250076 555620 250128 555626
rect 250076 555562 250128 555568
rect 248694 549944 248750 549953
rect 248694 549879 248750 549888
rect 248708 547963 248736 549879
rect 249432 548208 249484 548214
rect 249432 548150 249484 548156
rect 249444 547963 249472 548150
rect 250088 547963 250116 555562
rect 250812 554192 250864 554198
rect 250812 554134 250864 554140
rect 250824 547963 250852 554134
rect 251548 552968 251600 552974
rect 251548 552910 251600 552916
rect 251560 547963 251588 552910
rect 252284 551472 252336 551478
rect 252284 551414 252336 551420
rect 252296 547963 252324 551414
rect 252928 550112 252980 550118
rect 252928 550054 252980 550060
rect 252940 547963 252968 550054
rect 253676 547963 253704 557506
rect 255332 552906 255360 563790
rect 256700 558408 256752 558414
rect 256700 558350 256752 558356
rect 255320 552900 255372 552906
rect 255320 552842 255372 552848
rect 256516 552900 256568 552906
rect 256516 552842 256568 552848
rect 255872 550792 255924 550798
rect 255872 550734 255924 550740
rect 255134 549672 255190 549681
rect 255134 549607 255190 549616
rect 254400 548344 254452 548350
rect 254400 548286 254452 548292
rect 254412 547963 254440 548286
rect 255148 547963 255176 549607
rect 255884 547963 255912 550734
rect 256528 547963 256556 552842
rect 256712 552566 256740 558350
rect 260116 555694 260144 564402
rect 260852 557534 260880 567938
rect 262784 564466 262812 568126
rect 265360 564466 265388 568126
rect 267740 565888 267792 565894
rect 267740 565830 267792 565836
rect 262772 564460 262824 564466
rect 262772 564402 262824 564408
rect 264244 564460 264296 564466
rect 264244 564402 264296 564408
rect 265348 564460 265400 564466
rect 265348 564402 265400 564408
rect 267004 564460 267056 564466
rect 267004 564402 267056 564408
rect 263600 561060 263652 561066
rect 263600 561002 263652 561008
rect 263612 557534 263640 561002
rect 260852 557506 261616 557534
rect 263612 557506 263732 557534
rect 260196 556980 260248 556986
rect 260196 556922 260248 556928
rect 260104 555688 260156 555694
rect 260104 555630 260156 555636
rect 259460 552968 259512 552974
rect 259460 552910 259512 552916
rect 256700 552560 256752 552566
rect 256700 552502 256752 552508
rect 257988 552560 258040 552566
rect 257988 552502 258040 552508
rect 257252 550248 257304 550254
rect 257252 550190 257304 550196
rect 257264 547963 257292 550190
rect 258000 547963 258028 552502
rect 258722 549808 258778 549817
rect 258722 549743 258778 549752
rect 258736 547963 258764 549743
rect 259472 547963 259500 552910
rect 260208 548162 260236 556922
rect 260840 548412 260892 548418
rect 260840 548354 260892 548360
rect 260132 548134 260236 548162
rect 260132 547944 260160 548134
rect 260852 547963 260880 548354
rect 261588 547963 261616 557506
rect 263048 550928 263100 550934
rect 263048 550870 263100 550876
rect 262312 550316 262364 550322
rect 262312 550258 262364 550264
rect 262324 547963 262352 550258
rect 263060 547963 263088 550870
rect 263704 547963 263732 557506
rect 264256 555490 264284 564402
rect 266360 562624 266412 562630
rect 266360 562566 266412 562572
rect 264244 555484 264296 555490
rect 264244 555426 264296 555432
rect 266372 552786 266400 562566
rect 266452 559836 266504 559842
rect 266452 559778 266504 559784
rect 266464 557534 266492 559778
rect 266464 557506 266860 557534
rect 266372 552758 266584 552786
rect 264428 550860 264480 550866
rect 264428 550802 264480 550808
rect 264440 547963 264468 550802
rect 266360 549500 266412 549506
rect 266360 549442 266412 549448
rect 265900 548684 265952 548690
rect 265900 548626 265952 548632
rect 265164 548480 265216 548486
rect 265164 548422 265216 548428
rect 265176 547963 265204 548422
rect 265912 547963 265940 548626
rect 266372 548554 266400 549442
rect 266360 548548 266412 548554
rect 266360 548490 266412 548496
rect 266556 547963 266584 552758
rect 266832 552650 266860 557506
rect 267016 552770 267044 564402
rect 267752 557534 267780 565830
rect 268672 564466 268700 568126
rect 269120 565276 269172 565282
rect 269120 565218 269172 565224
rect 268660 564460 268712 564466
rect 268660 564402 268712 564408
rect 269132 557534 269160 565218
rect 271248 564466 271276 568126
rect 269764 564460 269816 564466
rect 269764 564402 269816 564408
rect 271236 564460 271288 564466
rect 271236 564402 271288 564408
rect 267752 557506 268056 557534
rect 269132 557506 269528 557534
rect 267004 552764 267056 552770
rect 267004 552706 267056 552712
rect 266832 552622 267320 552650
rect 267292 547963 267320 552622
rect 268028 547963 268056 557506
rect 268752 548752 268804 548758
rect 268752 548694 268804 548700
rect 268764 547963 268792 548694
rect 269500 547963 269528 557506
rect 269776 554062 269804 564402
rect 274652 562426 274680 568126
rect 276952 565146 276980 568126
rect 276940 565140 276992 565146
rect 276940 565082 276992 565088
rect 280264 564466 280292 568126
rect 278044 564460 278096 564466
rect 278044 564402 278096 564408
rect 280252 564460 280304 564466
rect 280252 564402 280304 564408
rect 274824 563984 274876 563990
rect 274824 563926 274876 563932
rect 274836 563054 274864 563926
rect 274836 563026 275232 563054
rect 274640 562420 274692 562426
rect 274640 562362 274692 562368
rect 273260 559768 273312 559774
rect 273260 559710 273312 559716
rect 270132 555484 270184 555490
rect 270132 555426 270184 555432
rect 269764 554056 269816 554062
rect 269764 553998 269816 554004
rect 270144 547963 270172 555426
rect 273272 552770 273300 559710
rect 273260 552764 273312 552770
rect 273260 552706 273312 552712
rect 274456 552764 274508 552770
rect 274456 552706 274508 552712
rect 271604 551404 271656 551410
rect 271604 551346 271656 551352
rect 270868 550180 270920 550186
rect 270868 550122 270920 550128
rect 270880 547963 270908 550122
rect 271616 547963 271644 551346
rect 273076 551064 273128 551070
rect 273076 551006 273128 551012
rect 272340 550996 272392 551002
rect 272340 550938 272392 550944
rect 272352 547963 272380 550938
rect 273088 547963 273116 551006
rect 273720 549636 273772 549642
rect 273720 549578 273772 549584
rect 273260 549364 273312 549370
rect 273260 549306 273312 549312
rect 273272 548622 273300 549306
rect 273260 548616 273312 548622
rect 273260 548558 273312 548564
rect 273732 547963 273760 549578
rect 274468 547963 274496 552706
rect 275204 547963 275232 563026
rect 278056 552702 278084 564402
rect 279516 558476 279568 558482
rect 279516 558418 279568 558424
rect 278044 552696 278096 552702
rect 278044 552638 278096 552644
rect 278780 550656 278832 550662
rect 278780 550598 278832 550604
rect 278044 549840 278096 549846
rect 278044 549782 278096 549788
rect 277308 549772 277360 549778
rect 277308 549714 277360 549720
rect 276572 549704 276624 549710
rect 276572 549646 276624 549652
rect 275928 549500 275980 549506
rect 275928 549442 275980 549448
rect 275940 547963 275968 549442
rect 276584 547963 276612 549646
rect 277320 547963 277348 549714
rect 278056 547963 278084 549782
rect 278792 547963 278820 550598
rect 279528 547963 279556 558418
rect 280724 553394 280752 630294
rect 280816 563922 280844 630414
rect 280894 600400 280950 600409
rect 280894 600335 280950 600344
rect 280804 563916 280856 563922
rect 280804 563858 280856 563864
rect 280908 558226 280936 600335
rect 281000 562986 281028 640319
rect 281538 628008 281594 628017
rect 281538 627943 281594 627952
rect 281170 572860 281226 572869
rect 281170 572795 281226 572804
rect 281078 570072 281134 570081
rect 281078 570007 281134 570016
rect 281092 568070 281120 570007
rect 281080 568064 281132 568070
rect 281080 568006 281132 568012
rect 281184 567194 281212 572795
rect 281092 567166 281212 567194
rect 281092 563054 281120 567166
rect 281552 563718 281580 627943
rect 282918 625288 282974 625297
rect 282918 625223 282974 625232
rect 281630 618488 281686 618497
rect 281630 618423 281686 618432
rect 281540 563712 281592 563718
rect 281540 563654 281592 563660
rect 281092 563026 281304 563054
rect 281000 562958 281212 562986
rect 280908 558198 281028 558226
rect 280724 553366 280936 553394
rect 280160 549432 280212 549438
rect 280160 549374 280212 549380
rect 280172 547963 280200 549374
rect 280908 547963 280936 553366
rect 281000 552838 281028 558198
rect 280988 552832 281040 552838
rect 280988 552774 281040 552780
rect 281184 549914 281212 562958
rect 281276 556918 281304 563026
rect 281540 562284 281592 562290
rect 281540 562226 281592 562232
rect 281264 556912 281316 556918
rect 281264 556854 281316 556860
rect 281552 551188 281580 562226
rect 281644 551342 281672 618423
rect 281722 615632 281778 615641
rect 281722 615567 281778 615576
rect 281736 566642 281764 615567
rect 281814 612776 281870 612785
rect 281814 612711 281870 612720
rect 281724 566636 281776 566642
rect 281724 566578 281776 566584
rect 281828 566506 281856 612711
rect 281906 594008 281962 594017
rect 281906 593943 281962 593952
rect 281920 566574 281948 593943
rect 281998 584488 282054 584497
rect 281998 584423 282054 584432
rect 281908 566568 281960 566574
rect 281908 566510 281960 566516
rect 281816 566500 281868 566506
rect 281816 566442 281868 566448
rect 282012 562358 282040 584423
rect 282090 581768 282146 581777
rect 282090 581703 282146 581712
rect 282104 562562 282132 581703
rect 282182 575648 282238 575657
rect 282182 575583 282238 575592
rect 282196 567866 282224 575583
rect 282184 567860 282236 567866
rect 282184 567802 282236 567808
rect 282092 562556 282144 562562
rect 282092 562498 282144 562504
rect 282000 562352 282052 562358
rect 282000 562294 282052 562300
rect 282932 558346 282960 625223
rect 283010 621208 283066 621217
rect 283010 621143 283066 621152
rect 283024 560998 283052 621143
rect 283102 608968 283158 608977
rect 283102 608903 283158 608912
rect 283012 560992 283064 560998
rect 283012 560934 283064 560940
rect 282920 558340 282972 558346
rect 282920 558282 282972 558288
rect 283116 558210 283144 608903
rect 283286 606384 283342 606393
rect 283286 606319 283342 606328
rect 283194 603120 283250 603129
rect 283194 603055 283250 603064
rect 283104 558204 283156 558210
rect 283104 558146 283156 558152
rect 283208 555558 283236 603055
rect 283300 563786 283328 606319
rect 283654 596728 283710 596737
rect 283654 596663 283710 596672
rect 283668 596222 283696 596663
rect 283656 596216 283708 596222
rect 283656 596158 283708 596164
rect 283378 590744 283434 590753
rect 283378 590679 283434 590688
rect 283288 563780 283340 563786
rect 283288 563722 283340 563728
rect 283392 559570 283420 590679
rect 283470 588024 283526 588033
rect 283470 587959 283526 587968
rect 283484 566710 283512 587959
rect 283562 578368 283618 578377
rect 283562 578303 283618 578312
rect 283576 567934 283604 578303
rect 283564 567928 283616 567934
rect 283564 567870 283616 567876
rect 283472 566704 283524 566710
rect 283472 566646 283524 566652
rect 283380 559564 283432 559570
rect 283380 559506 283432 559512
rect 283196 555552 283248 555558
rect 283196 555494 283248 555500
rect 283104 552356 283156 552362
rect 283104 552298 283156 552304
rect 281632 551336 281684 551342
rect 281632 551278 281684 551284
rect 281552 551160 282408 551188
rect 281172 549908 281224 549914
rect 281172 549850 281224 549856
rect 281632 549908 281684 549914
rect 281632 549850 281684 549856
rect 281644 547963 281672 549850
rect 282380 547963 282408 551160
rect 283116 547963 283144 552298
rect 284116 552288 284168 552294
rect 284116 552230 284168 552236
rect 283748 552084 283800 552090
rect 283748 552026 283800 552032
rect 283760 547963 283788 552026
rect 284128 549982 284156 552230
rect 284956 550050 284984 643078
rect 289820 641776 289872 641782
rect 289820 641718 289872 641724
rect 287704 641232 287756 641238
rect 287704 641174 287756 641180
rect 287060 639192 287112 639198
rect 287060 639134 287112 639140
rect 286324 604512 286376 604518
rect 286324 604454 286376 604460
rect 285036 594856 285088 594862
rect 285036 594798 285088 594804
rect 285048 562358 285076 594798
rect 285036 562352 285088 562358
rect 285036 562294 285088 562300
rect 286336 555490 286364 604454
rect 286416 589348 286468 589354
rect 286416 589290 286468 589296
rect 286428 568546 286456 589290
rect 286416 568540 286468 568546
rect 286416 568482 286468 568488
rect 286324 555484 286376 555490
rect 286324 555426 286376 555432
rect 285956 552424 286008 552430
rect 285956 552366 286008 552372
rect 285220 551336 285272 551342
rect 285220 551278 285272 551284
rect 284944 550044 284996 550050
rect 284944 549986 284996 549992
rect 284116 549976 284168 549982
rect 284116 549918 284168 549924
rect 284484 549364 284536 549370
rect 284484 549306 284536 549312
rect 284496 547963 284524 549306
rect 285232 547963 285260 551278
rect 285968 547963 285996 552366
rect 287072 551290 287100 639134
rect 287716 559842 287744 641174
rect 288440 637628 288492 637634
rect 288440 637570 288492 637576
rect 287796 614168 287848 614174
rect 287796 614110 287848 614116
rect 287704 559836 287756 559842
rect 287704 559778 287756 559784
rect 287808 552090 287836 614110
rect 287888 579692 287940 579698
rect 287888 579634 287940 579640
rect 287900 556986 287928 579634
rect 288452 557534 288480 637570
rect 289084 585200 289136 585206
rect 289084 585142 289136 585148
rect 289096 565282 289124 585142
rect 289084 565276 289136 565282
rect 289084 565218 289136 565224
rect 289832 557534 289860 641718
rect 302884 640824 302936 640830
rect 302884 640766 302936 640772
rect 298100 639600 298152 639606
rect 298100 639542 298152 639548
rect 296720 639532 296772 639538
rect 296720 639474 296772 639480
rect 291200 639464 291252 639470
rect 291200 639406 291252 639412
rect 288452 557506 288848 557534
rect 289832 557506 290228 557534
rect 287888 556980 287940 556986
rect 287888 556922 287940 556928
rect 287796 552084 287848 552090
rect 287796 552026 287848 552032
rect 287072 551262 288112 551290
rect 287336 551200 287388 551206
rect 287336 551142 287388 551148
rect 286690 549400 286746 549409
rect 286690 549335 286746 549344
rect 286704 547963 286732 549335
rect 287348 547963 287376 551142
rect 288084 547963 288112 551262
rect 288820 547963 288848 557506
rect 289544 552492 289596 552498
rect 289544 552434 289596 552440
rect 289556 547963 289584 552434
rect 290200 547963 290228 557506
rect 291212 550730 291240 639406
rect 293960 639260 294012 639266
rect 293960 639202 294012 639208
rect 293972 552770 294000 639202
rect 294604 627972 294656 627978
rect 294604 627914 294656 627920
rect 294616 558482 294644 627914
rect 295984 608660 296036 608666
rect 295984 608602 296036 608608
rect 294604 558476 294656 558482
rect 294604 558418 294656 558424
rect 295996 555626 296024 608602
rect 296732 557534 296760 639474
rect 296732 557506 297404 557534
rect 295984 555620 296036 555626
rect 295984 555562 296036 555568
rect 293960 552764 294012 552770
rect 293960 552706 294012 552712
rect 295248 552764 295300 552770
rect 295248 552706 295300 552712
rect 293132 552560 293184 552566
rect 293132 552502 293184 552508
rect 292488 551336 292540 551342
rect 292488 551278 292540 551284
rect 292500 551138 292528 551278
rect 291660 551132 291712 551138
rect 291660 551074 291712 551080
rect 292396 551132 292448 551138
rect 292396 551074 292448 551080
rect 292488 551132 292540 551138
rect 292488 551074 292540 551080
rect 291200 550724 291252 550730
rect 291200 550666 291252 550672
rect 290922 549536 290978 549545
rect 290922 549471 290978 549480
rect 290936 547963 290964 549471
rect 291672 547963 291700 551074
rect 292408 551018 292436 551074
rect 292408 550990 292528 551018
rect 292500 550730 292528 550990
rect 292396 550724 292448 550730
rect 292396 550666 292448 550672
rect 292488 550724 292540 550730
rect 292488 550666 292540 550672
rect 292408 547963 292436 550666
rect 293144 547963 293172 552502
rect 293776 552084 293828 552090
rect 293776 552026 293828 552032
rect 293788 547963 293816 552026
rect 294510 548176 294566 548185
rect 294510 548111 294566 548120
rect 294524 547963 294552 548111
rect 295260 547963 295288 552706
rect 296720 549568 296772 549574
rect 296720 549510 296772 549516
rect 295984 548820 296036 548826
rect 295984 548762 296036 548768
rect 295996 547963 296024 548762
rect 296732 547963 296760 549510
rect 297376 547963 297404 557506
rect 298112 547963 298140 639542
rect 302240 596828 302292 596834
rect 302240 596770 302292 596776
rect 302252 596222 302280 596770
rect 302240 596216 302292 596222
rect 302240 596158 302292 596164
rect 302252 568478 302280 596158
rect 302240 568472 302292 568478
rect 302240 568414 302292 568420
rect 301412 550656 301464 550662
rect 301412 550598 301464 550604
rect 300492 550316 300544 550322
rect 300492 550258 300544 550264
rect 300306 550080 300362 550089
rect 300306 550015 300362 550024
rect 299572 549976 299624 549982
rect 299572 549918 299624 549924
rect 298836 549432 298888 549438
rect 298836 549374 298888 549380
rect 298848 547963 298876 549374
rect 299584 547963 299612 549918
rect 300216 549364 300268 549370
rect 300216 549306 300268 549312
rect 300124 548752 300176 548758
rect 300124 548694 300176 548700
rect 300136 525502 300164 548694
rect 300228 526726 300256 549306
rect 300320 527105 300348 550015
rect 300400 549772 300452 549778
rect 300400 549714 300452 549720
rect 300306 527096 300362 527105
rect 300306 527031 300362 527040
rect 300412 526794 300440 549714
rect 300400 526788 300452 526794
rect 300400 526730 300452 526736
rect 300216 526720 300268 526726
rect 300216 526662 300268 526668
rect 300504 526250 300532 550258
rect 300676 549840 300728 549846
rect 300676 549782 300728 549788
rect 300582 549672 300638 549681
rect 300582 549607 300638 549616
rect 300596 528358 300624 549607
rect 300584 528352 300636 528358
rect 300584 528294 300636 528300
rect 300688 528290 300716 549782
rect 301228 548276 301280 548282
rect 301228 548218 301280 548224
rect 301240 542366 301268 548218
rect 301424 547874 301452 550598
rect 301964 550248 302016 550254
rect 301964 550190 302016 550196
rect 301688 549704 301740 549710
rect 301688 549646 301740 549652
rect 301502 549536 301558 549545
rect 301502 549471 301558 549480
rect 301412 547868 301464 547874
rect 301412 547810 301464 547816
rect 301228 542360 301280 542366
rect 301228 542302 301280 542308
rect 300676 528284 300728 528290
rect 300676 528226 300728 528232
rect 300492 526244 300544 526250
rect 300492 526186 300544 526192
rect 300124 525496 300176 525502
rect 300124 525438 300176 525444
rect 301516 524346 301544 549471
rect 301594 547904 301650 547913
rect 301594 547839 301650 547848
rect 301608 525162 301636 547839
rect 301700 526522 301728 549646
rect 301872 549636 301924 549642
rect 301872 549578 301924 549584
rect 301780 548684 301832 548690
rect 301780 548626 301832 548632
rect 301688 526516 301740 526522
rect 301688 526458 301740 526464
rect 301792 525366 301820 548626
rect 301884 527202 301912 549578
rect 301976 528222 302004 550190
rect 302056 549296 302108 549302
rect 302056 549238 302108 549244
rect 301964 528216 302016 528222
rect 301964 528158 302016 528164
rect 302068 528154 302096 549238
rect 302056 528148 302108 528154
rect 302056 528090 302108 528096
rect 301872 527196 301924 527202
rect 301872 527138 301924 527144
rect 301780 525360 301832 525366
rect 301780 525302 301832 525308
rect 301596 525156 301648 525162
rect 301596 525098 301648 525104
rect 301504 524340 301556 524346
rect 301504 524282 301556 524288
rect 44088 518220 44140 518226
rect 44088 518162 44140 518168
rect 57888 518220 57940 518226
rect 57888 518162 57940 518168
rect 43904 480072 43956 480078
rect 43904 480014 43956 480020
rect 43812 480004 43864 480010
rect 43812 479946 43864 479952
rect 42524 479732 42576 479738
rect 42524 479674 42576 479680
rect 42432 477216 42484 477222
rect 42432 477158 42484 477164
rect 42340 471912 42392 471918
rect 42340 471854 42392 471860
rect 41328 467560 41380 467566
rect 41328 467502 41380 467508
rect 41236 467492 41288 467498
rect 41236 467434 41288 467440
rect 41144 467356 41196 467362
rect 41144 467298 41196 467304
rect 41052 467288 41104 467294
rect 41052 467230 41104 467236
rect 41064 166394 41092 467230
rect 41052 166388 41104 166394
rect 41052 166330 41104 166336
rect 41156 166326 41184 467298
rect 41144 166320 41196 166326
rect 41144 166262 41196 166268
rect 21364 97980 21416 97986
rect 21364 97922 21416 97928
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 41248 57798 41276 467434
rect 41236 57792 41288 57798
rect 41236 57734 41288 57740
rect 41340 56574 41368 467502
rect 42248 467424 42300 467430
rect 42248 467366 42300 467372
rect 42260 268938 42288 467366
rect 42352 271794 42380 471854
rect 42340 271788 42392 271794
rect 42340 271730 42392 271736
rect 42444 271726 42472 477158
rect 42536 272882 42564 479674
rect 42616 477352 42668 477358
rect 42616 477294 42668 477300
rect 42524 272876 42576 272882
rect 42524 272818 42576 272824
rect 42432 271720 42484 271726
rect 42432 271662 42484 271668
rect 42248 268932 42300 268938
rect 42248 268874 42300 268880
rect 42628 251054 42656 477294
rect 43628 477148 43680 477154
rect 43628 477090 43680 477096
rect 43260 476876 43312 476882
rect 43260 476818 43312 476824
rect 42708 467628 42760 467634
rect 42708 467570 42760 467576
rect 42616 251048 42668 251054
rect 42616 250990 42668 250996
rect 41328 56568 41380 56574
rect 41328 56510 41380 56516
rect 42720 55010 42748 467570
rect 43272 391950 43300 476818
rect 43536 474496 43588 474502
rect 43536 474438 43588 474444
rect 43444 466064 43496 466070
rect 43444 466006 43496 466012
rect 43352 465928 43404 465934
rect 43352 465870 43404 465876
rect 43260 391944 43312 391950
rect 43260 391886 43312 391892
rect 43364 378010 43392 465870
rect 43352 378004 43404 378010
rect 43352 377946 43404 377952
rect 43456 377505 43484 466006
rect 43442 377496 43498 377505
rect 43442 377431 43498 377440
rect 43548 271862 43576 474438
rect 43536 271856 43588 271862
rect 43536 271798 43588 271804
rect 43640 268462 43668 477090
rect 43720 477080 43772 477086
rect 43720 477022 43772 477028
rect 43732 268530 43760 477022
rect 43824 268734 43852 479946
rect 43916 268802 43944 480014
rect 43996 477284 44048 477290
rect 43996 477226 44048 477232
rect 43904 268796 43956 268802
rect 43904 268738 43956 268744
rect 43812 268728 43864 268734
rect 43812 268670 43864 268676
rect 43720 268524 43772 268530
rect 43720 268466 43772 268472
rect 43628 268456 43680 268462
rect 43628 268398 43680 268404
rect 44008 251122 44036 477226
rect 44100 389842 44128 518162
rect 57900 517993 57928 518162
rect 57886 517984 57942 517993
rect 57886 517919 57942 517928
rect 302252 510513 302280 568414
rect 302896 562630 302924 640766
rect 302884 562624 302936 562630
rect 302884 562566 302936 562572
rect 302884 551064 302936 551070
rect 302884 551006 302936 551012
rect 302790 540424 302846 540433
rect 302790 540359 302846 540368
rect 302804 539646 302832 540359
rect 302792 539640 302844 539646
rect 302792 539582 302844 539588
rect 302330 525464 302386 525473
rect 302330 525399 302386 525408
rect 302344 523734 302372 525399
rect 302896 525298 302924 551006
rect 303160 549908 303212 549914
rect 303160 549850 303212 549856
rect 303066 549808 303122 549817
rect 303066 549743 303122 549752
rect 302976 548344 303028 548350
rect 302976 548286 303028 548292
rect 302884 525292 302936 525298
rect 302884 525234 302936 525240
rect 302988 525026 303016 548286
rect 303080 526969 303108 549743
rect 303066 526960 303122 526969
rect 303066 526895 303122 526904
rect 303172 526658 303200 549850
rect 304276 527270 304304 700266
rect 364352 643754 364380 702406
rect 401140 646536 401192 646542
rect 401140 646478 401192 646484
rect 364340 643748 364392 643754
rect 364340 643690 364392 643696
rect 317052 643204 317104 643210
rect 317052 643146 317104 643152
rect 311256 641164 311308 641170
rect 311256 641106 311308 641112
rect 309784 640552 309836 640558
rect 309784 640494 309836 640500
rect 307024 618316 307076 618322
rect 307024 618258 307076 618264
rect 307036 558278 307064 618258
rect 309796 558414 309824 640494
rect 311164 637696 311216 637702
rect 311164 637638 311216 637644
rect 309784 558408 309836 558414
rect 309784 558350 309836 558356
rect 307024 558272 307076 558278
rect 307024 558214 307076 558220
rect 311176 552974 311204 637638
rect 311268 561066 311296 641106
rect 312636 641096 312688 641102
rect 312636 641038 312688 641044
rect 312544 623824 312596 623830
rect 312544 623766 312596 623772
rect 311256 561060 311308 561066
rect 311256 561002 311308 561008
rect 311164 552968 311216 552974
rect 311164 552910 311216 552916
rect 309784 550724 309836 550730
rect 309784 550666 309836 550672
rect 304354 549400 304410 549409
rect 304354 549335 304410 549344
rect 304264 527264 304316 527270
rect 304264 527206 304316 527212
rect 303160 526652 303212 526658
rect 303160 526594 303212 526600
rect 302976 525020 303028 525026
rect 302976 524962 303028 524968
rect 304368 524414 304396 549335
rect 305644 548480 305696 548486
rect 305644 548422 305696 548428
rect 304448 548412 304500 548418
rect 304448 548354 304500 548360
rect 304460 524958 304488 548354
rect 305656 525638 305684 548422
rect 309796 526998 309824 550666
rect 311164 539640 311216 539646
rect 311164 539582 311216 539588
rect 309784 526992 309836 526998
rect 309784 526934 309836 526940
rect 305644 525632 305696 525638
rect 305644 525574 305696 525580
rect 304448 524952 304500 524958
rect 304448 524894 304500 524900
rect 304356 524408 304408 524414
rect 304356 524350 304408 524356
rect 302332 523728 302384 523734
rect 302332 523670 302384 523676
rect 311176 515438 311204 539582
rect 311164 515432 311216 515438
rect 311164 515374 311216 515380
rect 302238 510504 302294 510513
rect 302238 510439 302294 510448
rect 302238 495544 302294 495553
rect 302238 495479 302240 495488
rect 302292 495479 302294 495488
rect 302240 495450 302292 495456
rect 59372 488022 60214 488050
rect 60598 488022 60688 488050
rect 53748 485784 53800 485790
rect 53748 485726 53800 485732
rect 50896 485512 50948 485518
rect 50896 485454 50948 485460
rect 47860 482928 47912 482934
rect 47860 482870 47912 482876
rect 46664 482792 46716 482798
rect 46664 482734 46716 482740
rect 46572 482724 46624 482730
rect 46572 482666 46624 482672
rect 46388 482588 46440 482594
rect 46388 482530 46440 482536
rect 46296 482520 46348 482526
rect 46296 482462 46348 482468
rect 45928 482384 45980 482390
rect 45928 482326 45980 482332
rect 45468 480140 45520 480146
rect 45468 480082 45520 480088
rect 45100 474564 45152 474570
rect 45100 474506 45152 474512
rect 45008 472796 45060 472802
rect 45008 472738 45060 472744
rect 44824 468512 44876 468518
rect 44824 468454 44876 468460
rect 44732 465996 44784 466002
rect 44732 465938 44784 465944
rect 44640 416832 44692 416838
rect 44640 416774 44692 416780
rect 44088 389836 44140 389842
rect 44088 389778 44140 389784
rect 44100 281518 44128 389778
rect 44652 377330 44680 416774
rect 44744 377942 44772 465938
rect 44732 377936 44784 377942
rect 44732 377878 44784 377884
rect 44640 377324 44692 377330
rect 44640 377266 44692 377272
rect 44088 281512 44140 281518
rect 44088 281454 44140 281460
rect 44836 273494 44864 468454
rect 44916 467152 44968 467158
rect 44916 467094 44968 467100
rect 44824 273488 44876 273494
rect 44824 273430 44876 273436
rect 44928 268326 44956 467094
rect 45020 273290 45048 472738
rect 45112 273358 45140 474506
rect 45192 474088 45244 474094
rect 45192 474030 45244 474036
rect 45204 273426 45232 474030
rect 45284 472728 45336 472734
rect 45284 472670 45336 472676
rect 45192 273420 45244 273426
rect 45192 273362 45244 273368
rect 45100 273352 45152 273358
rect 45100 273294 45152 273300
rect 45008 273284 45060 273290
rect 45008 273226 45060 273232
rect 45296 272542 45324 472670
rect 45376 472660 45428 472666
rect 45376 472602 45428 472608
rect 45284 272536 45336 272542
rect 45284 272478 45336 272484
rect 45388 269006 45416 472602
rect 45376 269000 45428 269006
rect 45376 268942 45428 268948
rect 45480 268394 45508 480082
rect 45940 271289 45968 482326
rect 46112 479528 46164 479534
rect 46112 479470 46164 479476
rect 46020 469056 46072 469062
rect 46020 468998 46072 469004
rect 46032 383654 46060 468998
rect 46124 389162 46152 479470
rect 46204 471164 46256 471170
rect 46204 471106 46256 471112
rect 46112 389156 46164 389162
rect 46112 389098 46164 389104
rect 46032 383626 46152 383654
rect 46124 379409 46152 383626
rect 46110 379400 46166 379409
rect 46110 379335 46166 379344
rect 45926 271280 45982 271289
rect 45926 271215 45982 271224
rect 46124 271046 46152 379335
rect 46216 378622 46244 471106
rect 46204 378616 46256 378622
rect 46204 378558 46256 378564
rect 46308 303618 46336 482462
rect 46296 303612 46348 303618
rect 46296 303554 46348 303560
rect 46400 300830 46428 482530
rect 46480 479460 46532 479466
rect 46480 479402 46532 479408
rect 46388 300824 46440 300830
rect 46388 300766 46440 300772
rect 46492 271658 46520 479402
rect 46584 272406 46612 482666
rect 46676 272474 46704 482734
rect 46848 482452 46900 482458
rect 46848 482394 46900 482400
rect 46664 272468 46716 272474
rect 46664 272410 46716 272416
rect 46572 272400 46624 272406
rect 46572 272342 46624 272348
rect 46756 272196 46808 272202
rect 46756 272138 46808 272144
rect 46480 271652 46532 271658
rect 46480 271594 46532 271600
rect 46112 271040 46164 271046
rect 46112 270982 46164 270988
rect 45468 268388 45520 268394
rect 45468 268330 45520 268336
rect 44916 268320 44968 268326
rect 44916 268262 44968 268268
rect 46124 267734 46152 270982
rect 46664 269816 46716 269822
rect 46664 269758 46716 269764
rect 46480 268524 46532 268530
rect 46480 268466 46532 268472
rect 46124 267706 46428 267734
rect 43996 251116 44048 251122
rect 43996 251058 44048 251064
rect 46400 145858 46428 267706
rect 46492 164150 46520 268466
rect 46570 268424 46626 268433
rect 46570 268359 46626 268368
rect 46584 164218 46612 268359
rect 46572 164212 46624 164218
rect 46572 164154 46624 164160
rect 46480 164144 46532 164150
rect 46480 164086 46532 164092
rect 46676 148714 46704 269758
rect 46664 148708 46716 148714
rect 46664 148650 46716 148656
rect 46768 148646 46796 272138
rect 46860 268666 46888 482394
rect 47768 479596 47820 479602
rect 47768 479538 47820 479544
rect 47676 476944 47728 476950
rect 47676 476886 47728 476892
rect 47584 474632 47636 474638
rect 47584 474574 47636 474580
rect 47492 471096 47544 471102
rect 47492 471038 47544 471044
rect 47400 466540 47452 466546
rect 47400 466482 47452 466488
rect 47412 418130 47440 466482
rect 47400 418124 47452 418130
rect 47400 418066 47452 418072
rect 47400 411324 47452 411330
rect 47400 411266 47452 411272
rect 46940 378616 46992 378622
rect 46940 378558 46992 378564
rect 46952 378214 46980 378558
rect 46940 378208 46992 378214
rect 46940 378150 46992 378156
rect 46952 272202 46980 378150
rect 47412 377058 47440 411266
rect 47504 379273 47532 471038
rect 47490 379264 47546 379273
rect 47490 379199 47546 379208
rect 47400 377052 47452 377058
rect 47400 376994 47452 377000
rect 47504 373994 47532 379199
rect 47596 378554 47624 474574
rect 47688 379098 47716 476886
rect 47780 379438 47808 479538
rect 47768 379432 47820 379438
rect 47768 379374 47820 379380
rect 47676 379092 47728 379098
rect 47676 379034 47728 379040
rect 47584 378548 47636 378554
rect 47584 378490 47636 378496
rect 47504 373966 47808 373994
rect 47492 272468 47544 272474
rect 47492 272410 47544 272416
rect 46940 272196 46992 272202
rect 46940 272138 46992 272144
rect 46952 271561 46980 272138
rect 46938 271552 46994 271561
rect 46938 271487 46994 271496
rect 46848 268660 46900 268666
rect 46848 268602 46900 268608
rect 46756 148640 46808 148646
rect 46756 148582 46808 148588
rect 46388 145852 46440 145858
rect 46388 145794 46440 145800
rect 47504 145382 47532 272410
rect 47676 272400 47728 272406
rect 47676 272342 47728 272348
rect 47688 271998 47716 272342
rect 47676 271992 47728 271998
rect 47676 271934 47728 271940
rect 47688 145450 47716 271934
rect 47780 270978 47808 373966
rect 47872 272746 47900 482870
rect 49240 482860 49292 482866
rect 49240 482802 49292 482808
rect 48134 482624 48190 482633
rect 48134 482559 48190 482568
rect 48042 482488 48098 482497
rect 48042 482423 48098 482432
rect 47952 479392 48004 479398
rect 47952 479334 48004 479340
rect 47860 272740 47912 272746
rect 47860 272682 47912 272688
rect 47768 270972 47820 270978
rect 47768 270914 47820 270920
rect 47780 146266 47808 270914
rect 47964 269074 47992 479334
rect 48056 271386 48084 482423
rect 48148 271454 48176 482559
rect 49056 479664 49108 479670
rect 49056 479606 49108 479612
rect 48964 477012 49016 477018
rect 48964 476954 49016 476960
rect 48228 469192 48280 469198
rect 48228 469134 48280 469140
rect 48240 467945 48268 469134
rect 48226 467936 48282 467945
rect 48226 467871 48282 467880
rect 48228 465724 48280 465730
rect 48228 465666 48280 465672
rect 48136 271448 48188 271454
rect 48136 271390 48188 271396
rect 48044 271380 48096 271386
rect 48044 271322 48096 271328
rect 47952 269068 48004 269074
rect 47952 269010 48004 269016
rect 47860 268456 47912 268462
rect 47860 268398 47912 268404
rect 47872 163742 47900 268398
rect 47860 163736 47912 163742
rect 47860 163678 47912 163684
rect 47768 146260 47820 146266
rect 47768 146202 47820 146208
rect 47676 145444 47728 145450
rect 47676 145386 47728 145392
rect 47492 145376 47544 145382
rect 47492 145318 47544 145324
rect 48240 59430 48268 465666
rect 48872 414044 48924 414050
rect 48872 413986 48924 413992
rect 48780 412820 48832 412826
rect 48780 412762 48832 412768
rect 48792 380662 48820 412762
rect 48884 380798 48912 413986
rect 48872 380792 48924 380798
rect 48872 380734 48924 380740
rect 48780 380656 48832 380662
rect 48780 380598 48832 380604
rect 48976 380322 49004 476954
rect 48964 380316 49016 380322
rect 48964 380258 49016 380264
rect 49068 378690 49096 479606
rect 49148 477488 49200 477494
rect 49148 477430 49200 477436
rect 49056 378684 49108 378690
rect 49056 378626 49108 378632
rect 49056 378548 49108 378554
rect 49056 378490 49108 378496
rect 49068 378282 49096 378490
rect 49056 378276 49108 378282
rect 49056 378218 49108 378224
rect 49068 271833 49096 378218
rect 49054 271824 49110 271833
rect 49054 271759 49110 271768
rect 49160 268870 49188 477430
rect 49252 272678 49280 482802
rect 49332 482656 49384 482662
rect 49332 482598 49384 482604
rect 49240 272672 49292 272678
rect 49240 272614 49292 272620
rect 49344 272066 49372 482598
rect 50160 482316 50212 482322
rect 50160 482258 50212 482264
rect 49608 471844 49660 471850
rect 49608 471786 49660 471792
rect 49516 471504 49568 471510
rect 49516 471446 49568 471452
rect 49424 468580 49476 468586
rect 49424 468522 49476 468528
rect 49332 272060 49384 272066
rect 49332 272002 49384 272008
rect 49238 271824 49294 271833
rect 49238 271759 49294 271768
rect 49148 268864 49200 268870
rect 49148 268806 49200 268812
rect 49160 162858 49188 268806
rect 49148 162852 49200 162858
rect 49148 162794 49200 162800
rect 49252 148578 49280 271759
rect 49240 148572 49292 148578
rect 49240 148514 49292 148520
rect 49344 145722 49372 272002
rect 49436 164801 49464 468522
rect 49528 166258 49556 471446
rect 49516 166252 49568 166258
rect 49516 166194 49568 166200
rect 49620 164898 49648 471786
rect 50068 471708 50120 471714
rect 50068 471650 50120 471656
rect 50080 465798 50108 471650
rect 50068 465792 50120 465798
rect 50068 465734 50120 465740
rect 50172 378894 50200 482258
rect 50436 482248 50488 482254
rect 50436 482190 50488 482196
rect 50344 479324 50396 479330
rect 50344 479266 50396 479272
rect 50252 474292 50304 474298
rect 50252 474234 50304 474240
rect 50160 378888 50212 378894
rect 50160 378830 50212 378836
rect 50264 271182 50292 474234
rect 50252 271176 50304 271182
rect 50252 271118 50304 271124
rect 50356 270502 50384 479266
rect 50448 272814 50476 482190
rect 50526 479496 50582 479505
rect 50526 479431 50582 479440
rect 50436 272808 50488 272814
rect 50436 272750 50488 272756
rect 50344 270496 50396 270502
rect 50344 270438 50396 270444
rect 50436 268592 50488 268598
rect 50436 268534 50488 268540
rect 50448 268394 50476 268534
rect 50436 268388 50488 268394
rect 50436 268330 50488 268336
rect 49608 164892 49660 164898
rect 49608 164834 49660 164840
rect 49422 164792 49478 164801
rect 49422 164727 49478 164736
rect 49332 145716 49384 145722
rect 49332 145658 49384 145664
rect 50448 144634 50476 268330
rect 50540 251190 50568 479431
rect 50804 471572 50856 471578
rect 50804 471514 50856 471520
rect 50712 469124 50764 469130
rect 50712 469066 50764 469072
rect 50620 468648 50672 468654
rect 50620 468590 50672 468596
rect 50528 251184 50580 251190
rect 50528 251126 50580 251132
rect 50540 165578 50568 251126
rect 50528 165572 50580 165578
rect 50528 165514 50580 165520
rect 50632 165481 50660 468590
rect 50724 467945 50752 469066
rect 50710 467936 50766 467945
rect 50710 467871 50766 467880
rect 50712 465792 50764 465798
rect 50712 465734 50764 465740
rect 50724 166190 50752 465734
rect 50816 166870 50844 471514
rect 50908 166938 50936 485454
rect 51632 485104 51684 485110
rect 51632 485046 51684 485052
rect 53470 485072 53526 485081
rect 50988 484424 51040 484430
rect 50988 484366 51040 484372
rect 50896 166932 50948 166938
rect 50896 166874 50948 166880
rect 50804 166864 50856 166870
rect 50804 166806 50856 166812
rect 50712 166184 50764 166190
rect 50712 166126 50764 166132
rect 50618 165472 50674 165481
rect 50618 165407 50674 165416
rect 50436 144628 50488 144634
rect 50436 144570 50488 144576
rect 48228 59424 48280 59430
rect 48228 59366 48280 59372
rect 51000 58750 51028 484366
rect 51540 466132 51592 466138
rect 51540 466074 51592 466080
rect 50988 58744 51040 58750
rect 50988 58686 51040 58692
rect 51552 57458 51580 466074
rect 51644 410854 51672 485046
rect 53470 485007 53526 485016
rect 51908 482996 51960 483002
rect 51908 482938 51960 482944
rect 51816 474360 51868 474366
rect 51816 474302 51868 474308
rect 51724 474224 51776 474230
rect 51724 474166 51776 474172
rect 51632 410848 51684 410854
rect 51632 410790 51684 410796
rect 51632 409896 51684 409902
rect 51632 409838 51684 409844
rect 51644 380594 51672 409838
rect 51632 380588 51684 380594
rect 51632 380530 51684 380536
rect 51630 378992 51686 379001
rect 51630 378927 51686 378936
rect 51644 282198 51672 378927
rect 51632 282192 51684 282198
rect 51632 282134 51684 282140
rect 51736 271250 51764 474166
rect 51828 271318 51856 474302
rect 51920 272610 51948 482938
rect 52276 471980 52328 471986
rect 52276 471922 52328 471928
rect 52184 471776 52236 471782
rect 52184 471718 52236 471724
rect 52092 471232 52144 471238
rect 52092 471174 52144 471180
rect 52000 465792 52052 465798
rect 52000 465734 52052 465740
rect 51908 272604 51960 272610
rect 51908 272546 51960 272552
rect 51908 271448 51960 271454
rect 51906 271416 51908 271425
rect 51960 271416 51962 271425
rect 51906 271351 51962 271360
rect 51816 271312 51868 271318
rect 51816 271254 51868 271260
rect 51724 271244 51776 271250
rect 51724 271186 51776 271192
rect 51816 270496 51868 270502
rect 51816 270438 51868 270444
rect 51828 270094 51856 270438
rect 51906 270328 51962 270337
rect 51906 270263 51962 270272
rect 51816 270088 51868 270094
rect 51816 270030 51868 270036
rect 51632 165572 51684 165578
rect 51632 165514 51684 165520
rect 51644 164286 51672 165514
rect 51632 164280 51684 164286
rect 51632 164222 51684 164228
rect 51644 58886 51672 164222
rect 51724 146260 51776 146266
rect 51724 146202 51776 146208
rect 51736 145790 51764 146202
rect 51724 145784 51776 145790
rect 51724 145726 51776 145732
rect 51632 58880 51684 58886
rect 51632 58822 51684 58828
rect 51540 57452 51592 57458
rect 51540 57394 51592 57400
rect 42708 55004 42760 55010
rect 42708 54946 42760 54952
rect 51736 54602 51764 145726
rect 51828 144838 51856 270030
rect 51816 144832 51868 144838
rect 51816 144774 51868 144780
rect 51920 144770 51948 270263
rect 52012 167006 52040 465734
rect 52000 167000 52052 167006
rect 52000 166942 52052 166948
rect 52104 164830 52132 471174
rect 52196 164966 52224 471718
rect 52288 465798 52316 471922
rect 52920 471640 52972 471646
rect 52920 471582 52972 471588
rect 52932 467974 52960 471582
rect 53104 471300 53156 471306
rect 53104 471242 53156 471248
rect 52920 467968 52972 467974
rect 52920 467910 52972 467916
rect 52368 466336 52420 466342
rect 52368 466278 52420 466284
rect 52276 465792 52328 465798
rect 52276 465734 52328 465740
rect 52380 465225 52408 466278
rect 53012 465792 53064 465798
rect 53012 465734 53064 465740
rect 52366 465216 52422 465225
rect 52366 465151 52422 465160
rect 52920 464704 52972 464710
rect 52920 464646 52972 464652
rect 52276 464364 52328 464370
rect 52276 464306 52328 464312
rect 52288 380390 52316 464306
rect 52368 408536 52420 408542
rect 52368 408478 52420 408484
rect 52380 380905 52408 408478
rect 52366 380896 52422 380905
rect 52366 380831 52422 380840
rect 52276 380384 52328 380390
rect 52276 380326 52328 380332
rect 52274 379536 52330 379545
rect 52274 379471 52330 379480
rect 52184 164960 52236 164966
rect 52184 164902 52236 164908
rect 52092 164824 52144 164830
rect 52092 164766 52144 164772
rect 52184 164144 52236 164150
rect 52184 164086 52236 164092
rect 52196 163606 52224 164086
rect 52184 163600 52236 163606
rect 52184 163542 52236 163548
rect 52000 148640 52052 148646
rect 52000 148582 52052 148588
rect 51908 144764 51960 144770
rect 51908 144706 51960 144712
rect 52012 56030 52040 148582
rect 52196 56506 52224 163542
rect 52288 57866 52316 379471
rect 52932 271522 52960 464646
rect 52920 271516 52972 271522
rect 52920 271458 52972 271464
rect 52366 271416 52422 271425
rect 53024 271386 53052 465734
rect 53116 271454 53144 471242
rect 53286 471200 53342 471209
rect 53286 471135 53342 471144
rect 53196 468784 53248 468790
rect 53196 468726 53248 468732
rect 53104 271448 53156 271454
rect 53104 271390 53156 271396
rect 52366 271351 52422 271360
rect 52460 271380 52512 271386
rect 52380 163470 52408 271351
rect 52460 271322 52512 271328
rect 53012 271380 53064 271386
rect 53012 271322 53064 271328
rect 52472 271153 52500 271322
rect 52458 271144 52514 271153
rect 52458 271079 52514 271088
rect 52826 271144 52882 271153
rect 52826 271079 52882 271088
rect 52840 163946 52868 271079
rect 53104 268388 53156 268394
rect 53104 268330 53156 268336
rect 53116 267753 53144 268330
rect 53102 267744 53158 267753
rect 53102 267679 53158 267688
rect 52920 252000 52972 252006
rect 52920 251942 52972 251948
rect 52932 251054 52960 251942
rect 52920 251048 52972 251054
rect 52920 250990 52972 250996
rect 52828 163940 52880 163946
rect 52828 163882 52880 163888
rect 52932 163878 52960 250990
rect 52920 163872 52972 163878
rect 52920 163814 52972 163820
rect 52368 163464 52420 163470
rect 52368 163406 52420 163412
rect 53012 148368 53064 148374
rect 53012 148310 53064 148316
rect 52920 146124 52972 146130
rect 52920 146066 52972 146072
rect 52368 145852 52420 145858
rect 52368 145794 52420 145800
rect 52276 57860 52328 57866
rect 52276 57802 52328 57808
rect 52380 57322 52408 145794
rect 52368 57316 52420 57322
rect 52368 57258 52420 57264
rect 52184 56500 52236 56506
rect 52184 56442 52236 56448
rect 52000 56024 52052 56030
rect 52000 55966 52052 55972
rect 52932 54806 52960 146066
rect 53024 55214 53052 148310
rect 53116 144702 53144 267679
rect 53208 165170 53236 468726
rect 53300 165374 53328 471135
rect 53380 467968 53432 467974
rect 53380 467910 53432 467916
rect 53288 165368 53340 165374
rect 53288 165310 53340 165316
rect 53196 165164 53248 165170
rect 53196 165106 53248 165112
rect 53288 164212 53340 164218
rect 53288 164154 53340 164160
rect 53300 163538 53328 164154
rect 53392 164150 53420 467910
rect 53484 165345 53512 485007
rect 53564 479868 53616 479874
rect 53564 479810 53616 479816
rect 53576 379030 53604 479810
rect 53656 466404 53708 466410
rect 53656 466346 53708 466352
rect 53668 466041 53696 466346
rect 53654 466032 53710 466041
rect 53654 465967 53710 465976
rect 53656 465860 53708 465866
rect 53656 465802 53708 465808
rect 53564 379024 53616 379030
rect 53564 378966 53616 378972
rect 53562 378856 53618 378865
rect 53562 378791 53618 378800
rect 53470 165336 53526 165345
rect 53470 165271 53526 165280
rect 53380 164144 53432 164150
rect 53380 164086 53432 164092
rect 53380 163736 53432 163742
rect 53380 163678 53432 163684
rect 53288 163532 53340 163538
rect 53288 163474 53340 163480
rect 53196 148572 53248 148578
rect 53196 148514 53248 148520
rect 53104 144696 53156 144702
rect 53104 144638 53156 144644
rect 53012 55208 53064 55214
rect 53012 55150 53064 55156
rect 52920 54800 52972 54806
rect 52920 54742 52972 54748
rect 53208 54670 53236 148514
rect 53300 57662 53328 163474
rect 53288 57656 53340 57662
rect 53288 57598 53340 57604
rect 53392 56370 53420 163678
rect 53472 162852 53524 162858
rect 53472 162794 53524 162800
rect 53484 162178 53512 162794
rect 53472 162172 53524 162178
rect 53472 162114 53524 162120
rect 53380 56364 53432 56370
rect 53380 56306 53432 56312
rect 53484 55078 53512 162114
rect 53576 58682 53604 378791
rect 53668 58818 53696 465802
rect 53656 58812 53708 58818
rect 53656 58754 53708 58760
rect 53564 58676 53616 58682
rect 53564 58618 53616 58624
rect 53760 57730 53788 485726
rect 56508 485716 56560 485722
rect 56508 485658 56560 485664
rect 56324 485580 56376 485586
rect 56324 485522 56376 485528
rect 56232 485444 56284 485450
rect 56232 485386 56284 485392
rect 55956 485240 56008 485246
rect 55956 485182 56008 485188
rect 54760 483744 54812 483750
rect 54760 483686 54812 483692
rect 54668 482180 54720 482186
rect 54668 482122 54720 482128
rect 54206 471472 54262 471481
rect 54206 471407 54262 471416
rect 53840 273148 53892 273154
rect 53840 273090 53892 273096
rect 53852 271726 53880 273090
rect 53932 272128 53984 272134
rect 53932 272070 53984 272076
rect 53840 271720 53892 271726
rect 53840 271662 53892 271668
rect 53944 271658 53972 272070
rect 53932 271652 53984 271658
rect 53932 271594 53984 271600
rect 53944 270450 53972 271594
rect 53944 270422 54064 270450
rect 53932 270292 53984 270298
rect 53932 270234 53984 270240
rect 53840 270224 53892 270230
rect 53840 270166 53892 270172
rect 53852 269074 53880 270166
rect 53840 269068 53892 269074
rect 53840 269010 53892 269016
rect 53944 268666 53972 270234
rect 53932 268660 53984 268666
rect 53932 268602 53984 268608
rect 54036 258074 54064 270422
rect 53852 258046 54064 258074
rect 53852 146130 53880 258046
rect 54220 165578 54248 471407
rect 54576 471368 54628 471374
rect 54576 471310 54628 471316
rect 54484 466200 54536 466206
rect 54484 466142 54536 466148
rect 54392 464432 54444 464438
rect 54392 464374 54444 464380
rect 54300 412752 54352 412758
rect 54300 412694 54352 412700
rect 54312 380866 54340 412694
rect 54300 380860 54352 380866
rect 54300 380802 54352 380808
rect 54404 380186 54432 464374
rect 54392 380180 54444 380186
rect 54392 380122 54444 380128
rect 54496 377874 54524 466142
rect 54484 377868 54536 377874
rect 54484 377810 54536 377816
rect 54392 271720 54444 271726
rect 54392 271662 54444 271668
rect 54208 165572 54260 165578
rect 54208 165514 54260 165520
rect 54404 164014 54432 271662
rect 54588 271590 54616 471310
rect 54576 271584 54628 271590
rect 54576 271526 54628 271532
rect 54680 271114 54708 482122
rect 54668 271108 54720 271114
rect 54668 271050 54720 271056
rect 54772 269278 54800 483686
rect 55034 471608 55090 471617
rect 55034 471543 55090 471552
rect 54852 468988 54904 468994
rect 54852 468930 54904 468936
rect 54760 269272 54812 269278
rect 54760 269214 54812 269220
rect 54576 269068 54628 269074
rect 54576 269010 54628 269016
rect 54484 268660 54536 268666
rect 54484 268602 54536 268608
rect 54392 164008 54444 164014
rect 54392 163950 54444 163956
rect 53840 146124 53892 146130
rect 53840 146066 53892 146072
rect 54496 144906 54524 268602
rect 54588 161474 54616 269010
rect 54864 165034 54892 468930
rect 54944 468852 54996 468858
rect 54944 468794 54996 468800
rect 54956 165238 54984 468794
rect 55048 165510 55076 471543
rect 55864 464636 55916 464642
rect 55864 464578 55916 464584
rect 55772 464568 55824 464574
rect 55772 464510 55824 464516
rect 55680 413976 55732 413982
rect 55680 413918 55732 413924
rect 55692 379982 55720 413918
rect 55680 379976 55732 379982
rect 55680 379918 55732 379924
rect 55784 379302 55812 464510
rect 55876 412758 55904 464578
rect 55864 412752 55916 412758
rect 55864 412694 55916 412700
rect 55864 410848 55916 410854
rect 55864 410790 55916 410796
rect 55772 379296 55824 379302
rect 55772 379238 55824 379244
rect 55128 303952 55180 303958
rect 55128 303894 55180 303900
rect 55140 282266 55168 303894
rect 55128 282260 55180 282266
rect 55128 282202 55180 282208
rect 55876 273562 55904 410790
rect 55968 381002 55996 485182
rect 56138 471336 56194 471345
rect 56138 471271 56194 471280
rect 56048 468920 56100 468926
rect 56048 468862 56100 468868
rect 55956 380996 56008 381002
rect 55956 380938 56008 380944
rect 55956 358760 56008 358766
rect 55956 358702 56008 358708
rect 55864 273556 55916 273562
rect 55864 273498 55916 273504
rect 55968 271658 55996 358702
rect 55956 271652 56008 271658
rect 55956 271594 56008 271600
rect 55956 270020 56008 270026
rect 55956 269962 56008 269968
rect 55968 269278 55996 269962
rect 55956 269272 56008 269278
rect 55956 269214 56008 269220
rect 55864 252204 55916 252210
rect 55864 252146 55916 252152
rect 55036 165504 55088 165510
rect 55036 165446 55088 165452
rect 54944 165232 54996 165238
rect 54944 165174 54996 165180
rect 54852 165028 54904 165034
rect 54852 164970 54904 164976
rect 55876 164082 55904 252146
rect 55864 164076 55916 164082
rect 55864 164018 55916 164024
rect 55036 164008 55088 164014
rect 55036 163950 55088 163956
rect 54588 161446 54984 161474
rect 54760 146260 54812 146266
rect 54760 146202 54812 146208
rect 54576 145716 54628 145722
rect 54576 145658 54628 145664
rect 54484 144900 54536 144906
rect 54484 144842 54536 144848
rect 54588 59566 54616 145658
rect 54668 145444 54720 145450
rect 54668 145386 54720 145392
rect 54680 59702 54708 145386
rect 54668 59696 54720 59702
rect 54668 59638 54720 59644
rect 54576 59560 54628 59566
rect 54576 59502 54628 59508
rect 54772 59498 54800 146202
rect 54956 145926 54984 161446
rect 54944 145920 54996 145926
rect 54944 145862 54996 145868
rect 54852 145376 54904 145382
rect 54852 145318 54904 145324
rect 54760 59492 54812 59498
rect 54760 59434 54812 59440
rect 53748 57724 53800 57730
rect 53748 57666 53800 57672
rect 54864 57254 54892 145318
rect 54852 57248 54904 57254
rect 54852 57190 54904 57196
rect 54956 56098 54984 145862
rect 55048 59634 55076 163950
rect 55128 163872 55180 163878
rect 55128 163814 55180 163820
rect 55036 59628 55088 59634
rect 55036 59570 55088 59576
rect 55140 57526 55168 163814
rect 55968 161474 55996 269214
rect 56060 165102 56088 468862
rect 56152 165209 56180 471271
rect 56244 166734 56272 485386
rect 56232 166728 56284 166734
rect 56232 166670 56284 166676
rect 56336 165306 56364 485522
rect 56416 485036 56468 485042
rect 56416 484978 56468 484984
rect 56324 165300 56376 165306
rect 56324 165242 56376 165248
rect 56138 165200 56194 165209
rect 56138 165135 56194 165144
rect 56048 165096 56100 165102
rect 56048 165038 56100 165044
rect 56428 164762 56456 484978
rect 56520 165442 56548 485658
rect 58532 484900 58584 484906
rect 58532 484842 58584 484848
rect 56876 481024 56928 481030
rect 56876 480966 56928 480972
rect 56600 477420 56652 477426
rect 56600 477362 56652 477368
rect 56612 402974 56640 477362
rect 56612 402946 56824 402974
rect 56796 388822 56824 402946
rect 56784 388816 56836 388822
rect 56784 388758 56836 388764
rect 56690 388648 56746 388657
rect 56690 388583 56746 388592
rect 56600 380860 56652 380866
rect 56600 380802 56652 380808
rect 56612 303958 56640 380802
rect 56600 303952 56652 303958
rect 56600 303894 56652 303900
rect 56704 252521 56732 388583
rect 56888 309913 56916 480966
rect 57336 479800 57388 479806
rect 57336 479742 57388 479748
rect 57060 476740 57112 476746
rect 57060 476682 57112 476688
rect 57072 413982 57100 476682
rect 57152 464500 57204 464506
rect 57152 464442 57204 464448
rect 57060 413976 57112 413982
rect 57060 413918 57112 413924
rect 56966 410408 57022 410417
rect 56966 410343 57022 410352
rect 56980 409902 57008 410343
rect 56968 409896 57020 409902
rect 56968 409838 57020 409844
rect 57164 378962 57192 464442
rect 57242 417344 57298 417353
rect 57242 417279 57298 417288
rect 57256 416838 57284 417279
rect 57244 416832 57296 416838
rect 57244 416774 57296 416780
rect 57348 393314 57376 479742
rect 58440 476672 58492 476678
rect 58440 476614 58492 476620
rect 57428 474428 57480 474434
rect 57428 474370 57480 474376
rect 57256 393286 57376 393314
rect 57256 387802 57284 393286
rect 57440 390386 57468 474370
rect 57796 474156 57848 474162
rect 57796 474098 57848 474104
rect 57704 471436 57756 471442
rect 57704 471378 57756 471384
rect 57612 469872 57664 469878
rect 57612 469814 57664 469820
rect 57520 467220 57572 467226
rect 57520 467162 57572 467168
rect 57428 390380 57480 390386
rect 57428 390322 57480 390328
rect 57532 390266 57560 467162
rect 57348 390238 57560 390266
rect 57348 388414 57376 390238
rect 57428 390108 57480 390114
rect 57428 390050 57480 390056
rect 57336 388408 57388 388414
rect 57336 388350 57388 388356
rect 57244 387796 57296 387802
rect 57244 387738 57296 387744
rect 57440 381954 57468 390050
rect 57624 389994 57652 469814
rect 57532 389966 57652 389994
rect 57532 388498 57560 389966
rect 57612 389836 57664 389842
rect 57612 389778 57664 389784
rect 57624 389745 57652 389778
rect 57610 389736 57666 389745
rect 57610 389671 57666 389680
rect 57612 389156 57664 389162
rect 57612 389098 57664 389104
rect 57624 389065 57652 389098
rect 57610 389056 57666 389065
rect 57610 388991 57666 389000
rect 57532 388470 57652 388498
rect 57520 388408 57572 388414
rect 57520 388350 57572 388356
rect 57428 381948 57480 381954
rect 57428 381890 57480 381896
rect 57152 378956 57204 378962
rect 57152 378898 57204 378904
rect 57152 357876 57204 357882
rect 57152 357818 57204 357824
rect 56874 309904 56930 309913
rect 56874 309839 56930 309848
rect 56888 296714 56916 309839
rect 56968 300824 57020 300830
rect 56968 300766 57020 300772
rect 56796 296686 56916 296714
rect 56690 252512 56746 252521
rect 56690 252447 56746 252456
rect 56796 209774 56824 296686
rect 56876 251116 56928 251122
rect 56876 251058 56928 251064
rect 56612 209746 56824 209774
rect 56612 203017 56640 209746
rect 56598 203008 56654 203017
rect 56598 202943 56654 202952
rect 56508 165436 56560 165442
rect 56508 165378 56560 165384
rect 56416 164756 56468 164762
rect 56416 164698 56468 164704
rect 56508 163940 56560 163946
rect 56508 163882 56560 163888
rect 55968 161446 56272 161474
rect 56244 151814 56272 161446
rect 56152 151786 56272 151814
rect 56046 146296 56102 146305
rect 56046 146231 56102 146240
rect 55864 144900 55916 144906
rect 55864 144842 55916 144848
rect 55876 59362 55904 144842
rect 56060 142154 56088 146231
rect 56152 145994 56180 151786
rect 56232 148504 56284 148510
rect 56232 148446 56284 148452
rect 56140 145988 56192 145994
rect 56140 145930 56192 145936
rect 56152 144514 56180 145930
rect 56244 144650 56272 148446
rect 56324 148436 56376 148442
rect 56324 148378 56376 148384
rect 56336 144786 56364 148378
rect 56416 145648 56468 145654
rect 56416 145590 56468 145596
rect 56428 144906 56456 145590
rect 56416 144900 56468 144906
rect 56416 144842 56468 144848
rect 56336 144758 56456 144786
rect 56244 144622 56364 144650
rect 56152 144486 56272 144514
rect 56060 142126 56180 142154
rect 55864 59356 55916 59362
rect 55864 59298 55916 59304
rect 56152 59022 56180 142126
rect 56140 59016 56192 59022
rect 56140 58958 56192 58964
rect 55128 57520 55180 57526
rect 55128 57462 55180 57468
rect 56244 56166 56272 144486
rect 56336 56438 56364 144622
rect 56324 56432 56376 56438
rect 56324 56374 56376 56380
rect 56232 56160 56284 56166
rect 56232 56102 56284 56108
rect 54944 56092 54996 56098
rect 54944 56034 54996 56040
rect 56428 55146 56456 144758
rect 56520 59090 56548 163882
rect 56612 96529 56640 202943
rect 56782 201376 56838 201385
rect 56782 201311 56838 201320
rect 56598 96520 56654 96529
rect 56598 96455 56654 96464
rect 56796 93809 56824 201311
rect 56888 164121 56916 251058
rect 56980 195265 57008 300766
rect 57164 271726 57192 357818
rect 57532 311137 57560 388350
rect 57518 311128 57574 311137
rect 57518 311063 57574 311072
rect 57336 303612 57388 303618
rect 57336 303554 57388 303560
rect 57348 296714 57376 303554
rect 57426 301608 57482 301617
rect 57426 301543 57482 301552
rect 57440 300830 57468 301543
rect 57428 300824 57480 300830
rect 57428 300766 57480 300772
rect 57348 296686 57468 296714
rect 57244 281512 57296 281518
rect 57244 281454 57296 281460
rect 57152 271720 57204 271726
rect 57152 271662 57204 271668
rect 57060 269884 57112 269890
rect 57060 269826 57112 269832
rect 57072 268734 57100 269826
rect 57060 268728 57112 268734
rect 57060 268670 57112 268676
rect 56966 195256 57022 195265
rect 56966 195191 57022 195200
rect 56874 164112 56930 164121
rect 56874 164047 56930 164056
rect 57072 162858 57100 268670
rect 57150 204232 57206 204241
rect 57150 204167 57206 204176
rect 57060 162852 57112 162858
rect 57060 162794 57112 162800
rect 57060 146192 57112 146198
rect 57060 146134 57112 146140
rect 56782 93800 56838 93809
rect 56782 93735 56838 93744
rect 56508 59084 56560 59090
rect 56508 59026 56560 59032
rect 56416 55140 56468 55146
rect 56416 55082 56468 55088
rect 53472 55072 53524 55078
rect 53472 55014 53524 55020
rect 57072 54874 57100 146134
rect 57164 97481 57192 204167
rect 57256 175409 57284 281454
rect 57334 198792 57390 198801
rect 57334 198727 57390 198736
rect 57242 175400 57298 175409
rect 57242 175335 57298 175344
rect 57244 163464 57296 163470
rect 57244 163406 57296 163412
rect 57150 97472 57206 97481
rect 57150 97407 57206 97416
rect 57256 59158 57284 163406
rect 57348 93401 57376 198727
rect 57440 196353 57468 296686
rect 57532 287054 57560 311063
rect 57624 305017 57652 388470
rect 57716 306785 57744 471378
rect 57808 307873 57836 474098
rect 57888 418124 57940 418130
rect 57888 418066 57940 418072
rect 57900 417217 57928 418066
rect 57886 417208 57942 417217
rect 57886 417143 57942 417152
rect 57886 414216 57942 414225
rect 57886 414151 57942 414160
rect 57900 414050 57928 414151
rect 57888 414044 57940 414050
rect 57888 413986 57940 413992
rect 57886 413264 57942 413273
rect 57886 413199 57942 413208
rect 57900 412826 57928 413199
rect 57888 412820 57940 412826
rect 57888 412762 57940 412768
rect 57886 411496 57942 411505
rect 57886 411431 57942 411440
rect 57900 411330 57928 411431
rect 57888 411324 57940 411330
rect 57888 411266 57940 411272
rect 57886 408640 57942 408649
rect 57886 408575 57942 408584
rect 57900 408542 57928 408575
rect 57888 408536 57940 408542
rect 57888 408478 57940 408484
rect 57888 391944 57940 391950
rect 57888 391886 57940 391892
rect 57900 391513 57928 391886
rect 57886 391504 57942 391513
rect 57886 391439 57942 391448
rect 58452 388482 58480 476614
rect 58544 388521 58572 484842
rect 58808 482112 58860 482118
rect 58808 482054 58860 482060
rect 58624 479936 58676 479942
rect 58624 479878 58676 479884
rect 58530 388512 58586 388521
rect 57888 388476 57940 388482
rect 57888 388418 57940 388424
rect 58440 388476 58492 388482
rect 58530 388447 58586 388456
rect 58440 388418 58492 388424
rect 57900 380934 57928 388418
rect 58532 387796 58584 387802
rect 58532 387738 58584 387744
rect 57888 380928 57940 380934
rect 57888 380870 57940 380876
rect 58544 380254 58572 387738
rect 58636 380526 58664 479878
rect 58716 472864 58768 472870
rect 58716 472806 58768 472812
rect 58624 380520 58676 380526
rect 58624 380462 58676 380468
rect 58532 380248 58584 380254
rect 58532 380190 58584 380196
rect 58624 357400 58676 357406
rect 58624 357342 58676 357348
rect 57794 307864 57850 307873
rect 57794 307799 57850 307808
rect 57702 306776 57758 306785
rect 57702 306711 57758 306720
rect 57610 305008 57666 305017
rect 57610 304943 57666 304952
rect 57610 303648 57666 303657
rect 57610 303583 57612 303592
rect 57664 303583 57666 303592
rect 57612 303554 57664 303560
rect 57532 287026 57652 287054
rect 57518 282296 57574 282305
rect 57518 282231 57574 282240
rect 57532 281518 57560 282231
rect 57520 281512 57572 281518
rect 57520 281454 57572 281460
rect 57624 277394 57652 287026
rect 57532 277366 57652 277394
rect 57532 204241 57560 277366
rect 57612 251864 57664 251870
rect 57612 251806 57664 251812
rect 57624 251122 57652 251806
rect 57612 251116 57664 251122
rect 57612 251058 57664 251064
rect 57518 204232 57574 204241
rect 57518 204167 57574 204176
rect 57716 199889 57744 306711
rect 57808 306374 57836 307799
rect 57808 306346 57928 306374
rect 57794 305008 57850 305017
rect 57794 304943 57850 304952
rect 57702 199880 57758 199889
rect 57702 199815 57758 199824
rect 57716 198801 57744 199815
rect 57702 198792 57758 198801
rect 57702 198727 57758 198736
rect 57808 198121 57836 304943
rect 57900 201385 57928 306346
rect 58532 282192 58584 282198
rect 58532 282134 58584 282140
rect 58544 272474 58572 282134
rect 58636 272950 58664 357342
rect 58728 284209 58756 472806
rect 58714 284200 58770 284209
rect 58714 284135 58770 284144
rect 58716 282260 58768 282266
rect 58716 282202 58768 282208
rect 58728 277394 58756 282202
rect 58820 282033 58848 482054
rect 59082 479904 59138 479913
rect 59082 479839 59138 479848
rect 58992 464840 59044 464846
rect 58992 464782 59044 464788
rect 58900 464772 58952 464778
rect 58900 464714 58952 464720
rect 58806 282024 58862 282033
rect 58806 281959 58862 281968
rect 58728 277366 58848 277394
rect 58820 273193 58848 277366
rect 58806 273184 58862 273193
rect 58806 273119 58862 273128
rect 58624 272944 58676 272950
rect 58624 272886 58676 272892
rect 58532 272468 58584 272474
rect 58532 272410 58584 272416
rect 57980 269952 58032 269958
rect 57980 269894 58032 269900
rect 57992 268802 58020 269894
rect 57980 268796 58032 268802
rect 57980 268738 58032 268744
rect 57886 201376 57942 201385
rect 57886 201311 57942 201320
rect 57794 198112 57850 198121
rect 57794 198047 57850 198056
rect 57426 196344 57482 196353
rect 57426 196279 57482 196288
rect 57334 93392 57390 93401
rect 57334 93327 57390 93336
rect 57440 90545 57468 196279
rect 57808 196194 57836 198047
rect 57716 196166 57836 196194
rect 57716 180794 57744 196166
rect 57794 195256 57850 195265
rect 57794 195191 57850 195200
rect 57624 180766 57744 180794
rect 57520 164076 57572 164082
rect 57520 164018 57572 164024
rect 57532 163985 57560 164018
rect 57518 163976 57574 163985
rect 57518 163911 57574 163920
rect 57532 163402 57560 163911
rect 57520 163396 57572 163402
rect 57520 163338 57572 163344
rect 57624 91089 57652 180766
rect 57702 164112 57758 164121
rect 57702 164047 57704 164056
rect 57756 164047 57758 164056
rect 57704 164018 57756 164024
rect 57610 91080 57666 91089
rect 57610 91015 57666 91024
rect 57426 90536 57482 90545
rect 57426 90471 57482 90480
rect 57808 88233 57836 195191
rect 57886 175400 57942 175409
rect 57886 175335 57942 175344
rect 57794 88224 57850 88233
rect 57794 88159 57850 88168
rect 57900 68921 57928 175335
rect 57992 146198 58020 268738
rect 58716 252544 58768 252550
rect 58716 252486 58768 252492
rect 58624 251932 58676 251938
rect 58624 251874 58676 251880
rect 58636 251161 58664 251874
rect 58622 251152 58678 251161
rect 58622 251087 58678 251096
rect 58636 164218 58664 251087
rect 58624 164212 58676 164218
rect 58624 164154 58676 164160
rect 57980 146192 58032 146198
rect 58728 146180 58756 252486
rect 58820 146305 58848 273119
rect 58912 166462 58940 464714
rect 59004 166802 59032 464782
rect 59096 177585 59124 479839
rect 59372 474026 59400 488022
rect 60004 485648 60056 485654
rect 60004 485590 60056 485596
rect 59728 480208 59780 480214
rect 59728 480150 59780 480156
rect 59360 474020 59412 474026
rect 59360 473962 59412 473968
rect 59174 471744 59230 471753
rect 59174 471679 59230 471688
rect 59082 177576 59138 177585
rect 59082 177511 59138 177520
rect 58992 166796 59044 166802
rect 58992 166738 59044 166744
rect 59188 166598 59216 471679
rect 59268 466268 59320 466274
rect 59268 466210 59320 466216
rect 59176 166592 59228 166598
rect 59176 166534 59228 166540
rect 58900 166456 58952 166462
rect 58900 166398 58952 166404
rect 59176 162852 59228 162858
rect 59176 162794 59228 162800
rect 59188 162246 59216 162794
rect 59176 162240 59228 162246
rect 59176 162182 59228 162188
rect 58806 146296 58862 146305
rect 58806 146231 58862 146240
rect 59082 146296 59138 146305
rect 59082 146231 59138 146240
rect 59096 146180 59124 146231
rect 58728 146152 59124 146180
rect 57980 146134 58032 146140
rect 57992 146062 58020 146134
rect 57980 146056 58032 146062
rect 57980 145998 58032 146004
rect 58714 145752 58770 145761
rect 58714 145687 58770 145696
rect 58624 145580 58676 145586
rect 58624 145522 58676 145528
rect 58636 144770 58664 145522
rect 58624 144764 58676 144770
rect 58624 144706 58676 144712
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57244 59152 57296 59158
rect 57244 59094 57296 59100
rect 57900 57934 57928 68847
rect 57244 57928 57296 57934
rect 57244 57870 57296 57876
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57060 54868 57112 54874
rect 57060 54810 57112 54816
rect 53196 54664 53248 54670
rect 53196 54606 53248 54612
rect 51724 54596 51776 54602
rect 51724 54538 51776 54544
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 57256 3466 57284 57870
rect 58636 54738 58664 144706
rect 58728 144634 58756 145687
rect 58898 145616 58954 145625
rect 58898 145551 58954 145560
rect 58808 145512 58860 145518
rect 58808 145454 58860 145460
rect 58820 144838 58848 145454
rect 58808 144832 58860 144838
rect 58808 144774 58860 144780
rect 58716 144628 58768 144634
rect 58716 144570 58768 144576
rect 58728 56234 58756 144570
rect 58716 56228 58768 56234
rect 58716 56170 58768 56176
rect 58820 55962 58848 144774
rect 58912 144702 58940 145551
rect 58900 144696 58952 144702
rect 58900 144638 58952 144644
rect 58912 58954 58940 144638
rect 58900 58948 58952 58954
rect 58900 58890 58952 58896
rect 59096 57594 59124 146152
rect 59188 59294 59216 162182
rect 59176 59288 59228 59294
rect 59176 59230 59228 59236
rect 59084 57588 59136 57594
rect 59084 57530 59136 57536
rect 59280 57390 59308 466210
rect 59544 388816 59596 388822
rect 59544 388758 59596 388764
rect 59360 381948 59412 381954
rect 59360 381890 59412 381896
rect 59372 357882 59400 381890
rect 59452 380996 59504 381002
rect 59452 380938 59504 380944
rect 59464 358766 59492 380938
rect 59556 380458 59584 388758
rect 59544 380452 59596 380458
rect 59544 380394 59596 380400
rect 59636 379976 59688 379982
rect 59636 379918 59688 379924
rect 59452 358760 59504 358766
rect 59452 358702 59504 358708
rect 59360 357876 59412 357882
rect 59360 357818 59412 357824
rect 59648 272882 59676 379918
rect 59740 379166 59768 480150
rect 59818 479632 59874 479641
rect 59818 479567 59874 479576
rect 59728 379160 59780 379166
rect 59728 379102 59780 379108
rect 59636 272876 59688 272882
rect 59636 272818 59688 272824
rect 59728 272468 59780 272474
rect 59728 272410 59780 272416
rect 59634 271280 59690 271289
rect 59634 271215 59690 271224
rect 59648 270609 59676 271215
rect 59634 270600 59690 270609
rect 59634 270535 59690 270544
rect 59358 164248 59414 164257
rect 59358 164183 59414 164192
rect 59372 163674 59400 164183
rect 59360 163668 59412 163674
rect 59360 163610 59412 163616
rect 59372 140865 59400 163610
rect 59648 145314 59676 270535
rect 59740 146266 59768 272410
rect 59832 270502 59860 479567
rect 59912 468716 59964 468722
rect 59912 468658 59964 468664
rect 59820 270496 59872 270502
rect 59820 270438 59872 270444
rect 59832 269822 59860 270438
rect 59820 269816 59872 269822
rect 59820 269758 59872 269764
rect 59924 166530 59952 468658
rect 60016 166666 60044 485590
rect 60660 483818 60688 488022
rect 61028 485178 61056 488036
rect 61120 488022 61502 488050
rect 61672 488022 61962 488050
rect 61016 485172 61068 485178
rect 61016 485114 61068 485120
rect 61120 484106 61148 488022
rect 60752 484078 61148 484106
rect 60648 483812 60700 483818
rect 60648 483754 60700 483760
rect 60752 466070 60780 484078
rect 61672 470594 61700 488022
rect 62120 484220 62172 484226
rect 62120 484162 62172 484168
rect 60844 470566 61700 470594
rect 60740 466064 60792 466070
rect 60740 466006 60792 466012
rect 60844 465934 60872 470566
rect 62132 466002 62160 484162
rect 62212 484152 62264 484158
rect 62212 484094 62264 484100
rect 62224 476814 62252 484094
rect 62316 478174 62344 488036
rect 62408 488022 62790 488050
rect 62960 488022 63250 488050
rect 63512 488022 63710 488050
rect 62408 484158 62436 488022
rect 62960 484226 62988 488022
rect 62948 484220 63000 484226
rect 62948 484162 63000 484168
rect 62396 484152 62448 484158
rect 62396 484094 62448 484100
rect 62304 478168 62356 478174
rect 62304 478110 62356 478116
rect 62212 476808 62264 476814
rect 62212 476750 62264 476756
rect 63512 466206 63540 488022
rect 64156 484974 64184 488036
rect 64248 488022 64538 488050
rect 64892 488022 64998 488050
rect 65076 488022 65458 488050
rect 65536 488022 65918 488050
rect 64144 484968 64196 484974
rect 64144 484910 64196 484916
rect 64248 470594 64276 488022
rect 64892 471102 64920 488022
rect 65076 484140 65104 488022
rect 64984 484112 65104 484140
rect 64984 471170 65012 484112
rect 65536 474638 65564 488022
rect 66364 485353 66392 488036
rect 66456 488022 66746 488050
rect 66824 488022 67206 488050
rect 66350 485344 66406 485353
rect 66350 485279 66406 485288
rect 66456 484140 66484 488022
rect 66272 484112 66484 484140
rect 65524 474632 65576 474638
rect 65524 474574 65576 474580
rect 64972 471164 65024 471170
rect 64972 471106 65024 471112
rect 64880 471096 64932 471102
rect 64880 471038 64932 471044
rect 63604 470566 64276 470594
rect 63604 469062 63632 470566
rect 63592 469056 63644 469062
rect 63592 468998 63644 469004
rect 63500 466200 63552 466206
rect 63500 466142 63552 466148
rect 66272 466138 66300 484112
rect 66824 470594 66852 488022
rect 66364 470566 66852 470594
rect 66364 467634 66392 470566
rect 66352 467628 66404 467634
rect 66352 467570 66404 467576
rect 67652 466274 67680 488036
rect 67836 488022 68126 488050
rect 68204 488022 68494 488050
rect 67732 484152 67784 484158
rect 67732 484094 67784 484100
rect 67744 468353 67772 484094
rect 67836 469849 67864 488022
rect 68204 484158 68232 488022
rect 68466 485752 68522 485761
rect 68466 485687 68522 485696
rect 68284 485308 68336 485314
rect 68284 485250 68336 485256
rect 68192 484152 68244 484158
rect 68192 484094 68244 484100
rect 68296 474570 68324 485250
rect 68376 484764 68428 484770
rect 68376 484706 68428 484712
rect 68284 474564 68336 474570
rect 68284 474506 68336 474512
rect 68388 474502 68416 484706
rect 68480 484430 68508 485687
rect 68940 484945 68968 488036
rect 69124 488022 69414 488050
rect 69584 488022 69874 488050
rect 69952 488022 70334 488050
rect 70596 488022 70702 488050
rect 70872 488022 71162 488050
rect 71240 488022 71622 488050
rect 71792 488022 72082 488050
rect 68926 484936 68982 484945
rect 68926 484871 68982 484880
rect 68468 484424 68520 484430
rect 68468 484366 68520 484372
rect 69020 484152 69072 484158
rect 69020 484094 69072 484100
rect 68376 474496 68428 474502
rect 68376 474438 68428 474444
rect 67822 469840 67878 469849
rect 67822 469775 67878 469784
rect 67730 468344 67786 468353
rect 67730 468279 67786 468288
rect 67640 466268 67692 466274
rect 67640 466210 67692 466216
rect 66260 466132 66312 466138
rect 66260 466074 66312 466080
rect 62120 465996 62172 466002
rect 62120 465938 62172 465944
rect 60832 465928 60884 465934
rect 60832 465870 60884 465876
rect 69032 465730 69060 484094
rect 69020 465724 69072 465730
rect 69020 465666 69072 465672
rect 69124 465633 69152 488022
rect 69584 484158 69612 488022
rect 69572 484152 69624 484158
rect 69572 484094 69624 484100
rect 69952 470594 69980 488022
rect 70400 484152 70452 484158
rect 70400 484094 70452 484100
rect 69216 470566 69980 470594
rect 69216 469169 69244 470566
rect 69202 469160 69258 469169
rect 69202 469095 69258 469104
rect 70412 466041 70440 484094
rect 70492 480412 70544 480418
rect 70492 480354 70544 480360
rect 70504 467566 70532 480354
rect 70596 469033 70624 488022
rect 70872 484158 70900 488022
rect 70860 484152 70912 484158
rect 70860 484094 70912 484100
rect 71240 480418 71268 488022
rect 71228 480412 71280 480418
rect 71228 480354 71280 480360
rect 70582 469024 70638 469033
rect 70582 468959 70638 468968
rect 70492 467560 70544 467566
rect 70492 467502 70544 467508
rect 71792 466449 71820 488022
rect 72424 484968 72476 484974
rect 72424 484910 72476 484916
rect 71872 484152 71924 484158
rect 71872 484094 71924 484100
rect 71884 467498 71912 484094
rect 71872 467492 71924 467498
rect 71872 467434 71924 467440
rect 71778 466440 71834 466449
rect 71778 466375 71834 466384
rect 70398 466032 70454 466041
rect 70398 465967 70454 465976
rect 72436 465730 72464 484910
rect 72528 484809 72556 488036
rect 72620 488022 72910 488050
rect 72514 484800 72570 484809
rect 72514 484735 72570 484744
rect 72620 484158 72648 488022
rect 72608 484152 72660 484158
rect 72608 484094 72660 484100
rect 73356 467129 73384 488036
rect 73816 485625 73844 488036
rect 74276 485790 74304 488036
rect 74264 485784 74316 485790
rect 74264 485726 74316 485732
rect 74356 485784 74408 485790
rect 74356 485726 74408 485732
rect 73802 485616 73858 485625
rect 73802 485551 73858 485560
rect 73894 485344 73950 485353
rect 73894 485279 73950 485288
rect 73804 484968 73856 484974
rect 73804 484910 73856 484916
rect 73816 467430 73844 484910
rect 73804 467424 73856 467430
rect 73804 467366 73856 467372
rect 73908 467362 73936 485279
rect 74368 471918 74396 485726
rect 74540 484152 74592 484158
rect 74540 484094 74592 484100
rect 74356 471912 74408 471918
rect 74356 471854 74408 471860
rect 73896 467356 73948 467362
rect 73896 467298 73948 467304
rect 73342 467120 73398 467129
rect 73342 467055 73398 467064
rect 74552 465905 74580 484094
rect 74644 466177 74672 488036
rect 74736 488022 75118 488050
rect 75288 488022 75578 488050
rect 74736 484158 74764 488022
rect 74724 484152 74776 484158
rect 74724 484094 74776 484100
rect 75288 470594 75316 488022
rect 76024 485489 76052 488036
rect 76208 488022 76498 488050
rect 76576 488022 76866 488050
rect 76010 485480 76066 485489
rect 76010 485415 76066 485424
rect 75920 484152 75972 484158
rect 75920 484094 75972 484100
rect 74736 470566 75316 470594
rect 74630 466168 74686 466177
rect 74630 466103 74686 466112
rect 74538 465896 74594 465905
rect 74736 465866 74764 470566
rect 75932 466342 75960 484094
rect 76208 470594 76236 488022
rect 76576 484158 76604 488022
rect 77312 485761 77340 488036
rect 77404 488022 77786 488050
rect 77864 488022 78246 488050
rect 78722 488022 78904 488050
rect 77298 485752 77354 485761
rect 77298 485687 77354 485696
rect 76654 484528 76710 484537
rect 76654 484463 76710 484472
rect 76564 484152 76616 484158
rect 76564 484094 76616 484100
rect 76668 470594 76696 484463
rect 77404 484106 77432 488022
rect 76024 470566 76236 470594
rect 76576 470566 76696 470594
rect 77312 484078 77432 484106
rect 75920 466336 75972 466342
rect 75920 466278 75972 466284
rect 74538 465831 74594 465840
rect 74724 465860 74776 465866
rect 74724 465802 74776 465808
rect 76024 465769 76052 470566
rect 76576 466313 76604 470566
rect 77312 466410 77340 484078
rect 77864 470594 77892 488022
rect 78036 484968 78088 484974
rect 78220 484968 78272 484974
rect 78088 484916 78220 484922
rect 78036 484910 78272 484916
rect 78048 484894 78260 484910
rect 78680 484220 78732 484226
rect 78680 484162 78732 484168
rect 77404 470566 77892 470594
rect 77404 468625 77432 470566
rect 78692 469130 78720 484162
rect 78772 484152 78824 484158
rect 78772 484094 78824 484100
rect 78680 469124 78732 469130
rect 78680 469066 78732 469072
rect 77390 468616 77446 468625
rect 77390 468551 77446 468560
rect 78784 468489 78812 484094
rect 78876 468897 78904 488022
rect 78968 488022 79074 488050
rect 79152 488022 79534 488050
rect 79704 488022 79994 488050
rect 80256 488022 80454 488050
rect 78968 484158 78996 488022
rect 78956 484152 79008 484158
rect 78956 484094 79008 484100
rect 79152 470594 79180 488022
rect 79324 485512 79376 485518
rect 79324 485454 79376 485460
rect 79232 485376 79284 485382
rect 79232 485318 79284 485324
rect 79244 484770 79272 485318
rect 79336 485042 79364 485454
rect 79324 485036 79376 485042
rect 79324 484978 79376 484984
rect 79232 484764 79284 484770
rect 79232 484706 79284 484712
rect 79704 484226 79732 488022
rect 79692 484220 79744 484226
rect 79692 484162 79744 484168
rect 78968 470566 79180 470594
rect 78862 468888 78918 468897
rect 78862 468823 78918 468832
rect 78968 468761 78996 470566
rect 80256 469198 80284 488022
rect 80808 484537 80836 488036
rect 81268 484838 81296 488036
rect 81728 484906 81756 488036
rect 81820 488022 82202 488050
rect 82280 488022 82662 488050
rect 82924 488022 83030 488050
rect 83200 488022 83490 488050
rect 83568 488022 83950 488050
rect 81716 484900 81768 484906
rect 81716 484842 81768 484848
rect 81256 484832 81308 484838
rect 81256 484774 81308 484780
rect 80794 484528 80850 484537
rect 80794 484463 80850 484472
rect 80704 483812 80756 483818
rect 80704 483754 80756 483760
rect 80244 469192 80296 469198
rect 80244 469134 80296 469140
rect 78954 468752 79010 468761
rect 78954 468687 79010 468696
rect 78770 468480 78826 468489
rect 78770 468415 78826 468424
rect 80716 467838 80744 483754
rect 81820 476114 81848 488022
rect 81544 476086 81848 476114
rect 81544 471238 81572 476086
rect 82280 471850 82308 488022
rect 82820 480888 82872 480894
rect 82820 480830 82872 480836
rect 82832 471986 82860 480830
rect 82820 471980 82872 471986
rect 82820 471922 82872 471928
rect 82268 471844 82320 471850
rect 82268 471786 82320 471792
rect 82924 471714 82952 488022
rect 82912 471708 82964 471714
rect 82912 471650 82964 471656
rect 83200 471510 83228 488022
rect 83568 480894 83596 488022
rect 84396 485042 84424 488036
rect 84488 488022 84870 488050
rect 84948 488022 85238 488050
rect 85714 488022 85804 488050
rect 84384 485036 84436 485042
rect 84384 484978 84436 484984
rect 83556 480888 83608 480894
rect 83556 480830 83608 480836
rect 84488 476114 84516 488022
rect 84304 476086 84516 476114
rect 84304 471782 84332 476086
rect 84292 471776 84344 471782
rect 84292 471718 84344 471724
rect 84948 471578 84976 488022
rect 85776 483014 85804 488022
rect 85684 482986 85804 483014
rect 85868 488022 86158 488050
rect 86328 488022 86618 488050
rect 86972 488022 87078 488050
rect 87156 488022 87446 488050
rect 87524 488022 87906 488050
rect 85580 480888 85632 480894
rect 85580 480830 85632 480836
rect 84936 471572 84988 471578
rect 84936 471514 84988 471520
rect 83188 471504 83240 471510
rect 83188 471446 83240 471452
rect 81532 471232 81584 471238
rect 81532 471174 81584 471180
rect 85592 468790 85620 480830
rect 85684 478394 85712 482986
rect 85684 478366 85804 478394
rect 85672 478236 85724 478242
rect 85672 478178 85724 478184
rect 85684 468994 85712 478178
rect 85776 471646 85804 478366
rect 85868 478242 85896 488022
rect 86328 480894 86356 488022
rect 86316 480888 86368 480894
rect 86316 480830 86368 480836
rect 85856 478236 85908 478242
rect 85856 478178 85908 478184
rect 85764 471640 85816 471646
rect 85764 471582 85816 471588
rect 85672 468988 85724 468994
rect 85672 468930 85724 468936
rect 86972 468926 87000 488022
rect 87156 476114 87184 488022
rect 87064 476086 87184 476114
rect 86960 468920 87012 468926
rect 86960 468862 87012 468868
rect 87064 468858 87092 476086
rect 87524 471209 87552 488022
rect 88352 485586 88380 488036
rect 88536 488022 88826 488050
rect 88340 485580 88392 485586
rect 88340 485522 88392 485528
rect 88432 480616 88484 480622
rect 88432 480558 88484 480564
rect 88444 471481 88472 480558
rect 88536 471617 88564 488022
rect 89180 485722 89208 488036
rect 89272 488022 89654 488050
rect 89824 488022 90114 488050
rect 89168 485716 89220 485722
rect 89168 485658 89220 485664
rect 89272 480622 89300 488022
rect 89260 480616 89312 480622
rect 89260 480558 89312 480564
rect 88522 471608 88578 471617
rect 88522 471543 88578 471552
rect 88430 471472 88486 471481
rect 88430 471407 88486 471416
rect 89824 471345 89852 488022
rect 90560 485450 90588 488036
rect 90744 488022 91034 488050
rect 90548 485444 90600 485450
rect 90548 485386 90600 485392
rect 89810 471336 89866 471345
rect 89810 471271 89866 471280
rect 87510 471200 87566 471209
rect 87510 471135 87566 471144
rect 90744 470594 90772 488022
rect 91388 485217 91416 488036
rect 91848 485654 91876 488036
rect 91940 488022 92322 488050
rect 92676 488022 92782 488050
rect 92952 488022 93242 488050
rect 93320 488022 93610 488050
rect 91836 485648 91888 485654
rect 91836 485590 91888 485596
rect 91374 485208 91430 485217
rect 91374 485143 91430 485152
rect 91940 471753 91968 488022
rect 92572 484220 92624 484226
rect 92572 484162 92624 484168
rect 92480 484152 92532 484158
rect 92480 484094 92532 484100
rect 91926 471744 91982 471753
rect 91926 471679 91982 471688
rect 89916 470566 90772 470594
rect 87052 468852 87104 468858
rect 87052 468794 87104 468800
rect 85580 468784 85632 468790
rect 85580 468726 85632 468732
rect 80704 467832 80756 467838
rect 80704 467774 80756 467780
rect 77300 466404 77352 466410
rect 77300 466346 77352 466352
rect 76562 466304 76618 466313
rect 76562 466239 76618 466248
rect 76010 465760 76066 465769
rect 72424 465724 72476 465730
rect 76010 465695 76066 465704
rect 72424 465666 72476 465672
rect 69110 465624 69166 465633
rect 69110 465559 69166 465568
rect 89916 464846 89944 470566
rect 89904 464840 89956 464846
rect 89904 464782 89956 464788
rect 92492 464778 92520 484094
rect 92584 468654 92612 484162
rect 92676 468722 92704 488022
rect 92952 484158 92980 488022
rect 93320 484226 93348 488022
rect 94056 485081 94084 488036
rect 94240 488022 94530 488050
rect 94608 488022 94990 488050
rect 94042 485072 94098 485081
rect 94042 485007 94098 485016
rect 93308 484220 93360 484226
rect 93308 484162 93360 484168
rect 92940 484152 92992 484158
rect 92940 484094 92992 484100
rect 93860 484152 93912 484158
rect 93860 484094 93912 484100
rect 92664 468716 92716 468722
rect 92664 468658 92716 468664
rect 92572 468648 92624 468654
rect 92572 468590 92624 468596
rect 93872 467294 93900 484094
rect 94240 470594 94268 488022
rect 94608 484158 94636 488022
rect 95344 485353 95372 488036
rect 95528 488022 95818 488050
rect 95330 485344 95386 485353
rect 95330 485279 95386 485288
rect 94596 484152 94648 484158
rect 94596 484094 94648 484100
rect 95528 479913 95556 488022
rect 96264 482118 96292 488036
rect 96724 482186 96752 488036
rect 97184 482254 97212 488036
rect 97552 482934 97580 488036
rect 97540 482928 97592 482934
rect 97540 482870 97592 482876
rect 98012 482866 98040 488036
rect 98472 483002 98500 488036
rect 98656 488022 98946 488050
rect 99422 488022 99512 488050
rect 98460 482996 98512 483002
rect 98460 482938 98512 482944
rect 98000 482860 98052 482866
rect 98000 482802 98052 482808
rect 97172 482248 97224 482254
rect 97172 482190 97224 482196
rect 96712 482180 96764 482186
rect 96712 482122 96764 482128
rect 96252 482112 96304 482118
rect 96252 482054 96304 482060
rect 95514 479904 95570 479913
rect 95514 479839 95570 479848
rect 98656 474298 98684 488022
rect 98644 474292 98696 474298
rect 98644 474234 98696 474240
rect 99484 474230 99512 488022
rect 99576 488022 99774 488050
rect 99576 474366 99604 488022
rect 100220 484974 100248 488036
rect 100680 485110 100708 488036
rect 100864 488022 101154 488050
rect 101232 488022 101522 488050
rect 101600 488022 101982 488050
rect 102336 488022 102442 488050
rect 100668 485104 100720 485110
rect 100668 485046 100720 485052
rect 100208 484968 100260 484974
rect 100208 484910 100260 484916
rect 100760 484152 100812 484158
rect 100760 484094 100812 484100
rect 99564 474360 99616 474366
rect 99564 474302 99616 474308
rect 99472 474224 99524 474230
rect 99472 474166 99524 474172
rect 93964 470566 94268 470594
rect 93964 468586 93992 470566
rect 93952 468580 94004 468586
rect 93952 468522 94004 468528
rect 93860 467288 93912 467294
rect 93860 467230 93912 467236
rect 92480 464772 92532 464778
rect 92480 464714 92532 464720
rect 100772 464710 100800 484094
rect 100864 465798 100892 488022
rect 101232 471306 101260 488022
rect 101600 484158 101628 488022
rect 101588 484152 101640 484158
rect 101588 484094 101640 484100
rect 102336 471374 102364 488022
rect 102888 485790 102916 488036
rect 102876 485784 102928 485790
rect 102876 485726 102928 485732
rect 103348 485246 103376 488036
rect 103624 488022 103730 488050
rect 103336 485240 103388 485246
rect 103336 485182 103388 485188
rect 103624 474434 103652 488022
rect 104176 485382 104204 488036
rect 104360 488022 104650 488050
rect 105004 488022 105110 488050
rect 104164 485376 104216 485382
rect 104164 485318 104216 485324
rect 103612 474428 103664 474434
rect 103612 474370 103664 474376
rect 102324 471368 102376 471374
rect 102324 471310 102376 471316
rect 101220 471300 101272 471306
rect 101220 471242 101272 471248
rect 104360 470594 104388 488022
rect 105004 474094 105032 488022
rect 105556 485314 105584 488036
rect 105648 488022 105938 488050
rect 105544 485308 105596 485314
rect 105544 485250 105596 485256
rect 104992 474088 105044 474094
rect 104992 474030 105044 474036
rect 105648 472802 105676 488022
rect 106280 484152 106332 484158
rect 106280 484094 106332 484100
rect 105636 472796 105688 472802
rect 105636 472738 105688 472744
rect 103716 470566 104388 470594
rect 103716 468518 103744 470566
rect 103704 468512 103756 468518
rect 103704 468454 103756 468460
rect 106292 467158 106320 484094
rect 106384 472734 106412 488036
rect 106476 488022 106858 488050
rect 106936 488022 107318 488050
rect 106372 472728 106424 472734
rect 106372 472670 106424 472676
rect 106476 472666 106504 488022
rect 106936 484158 106964 488022
rect 106924 484152 106976 484158
rect 106924 484094 106976 484100
rect 107660 484152 107712 484158
rect 107660 484094 107712 484100
rect 106464 472660 106516 472666
rect 106464 472602 106516 472608
rect 107672 468518 107700 484094
rect 107764 468654 107792 488036
rect 107856 488022 108146 488050
rect 108224 488022 108606 488050
rect 109082 488022 109172 488050
rect 107752 468648 107804 468654
rect 107752 468590 107804 468596
rect 107856 468586 107884 488022
rect 108224 484158 108252 488022
rect 108212 484152 108264 484158
rect 108212 484094 108264 484100
rect 109040 484152 109092 484158
rect 109040 484094 109092 484100
rect 109052 468722 109080 484094
rect 109144 471306 109172 488022
rect 109236 488022 109526 488050
rect 109604 488022 109894 488050
rect 109236 471374 109264 488022
rect 109604 484158 109632 488022
rect 110340 485110 110368 488036
rect 110616 488022 110814 488050
rect 110328 485104 110380 485110
rect 110328 485046 110380 485052
rect 109592 484152 109644 484158
rect 109592 484094 109644 484100
rect 110616 472870 110644 488022
rect 111260 482798 111288 488036
rect 111248 482792 111300 482798
rect 111248 482734 111300 482740
rect 111720 482730 111748 488036
rect 111708 482724 111760 482730
rect 111708 482666 111760 482672
rect 112088 482594 112116 488036
rect 112076 482588 112128 482594
rect 112076 482530 112128 482536
rect 112548 482526 112576 488036
rect 112640 488022 113022 488050
rect 112536 482520 112588 482526
rect 112536 482462 112588 482468
rect 110604 472864 110656 472870
rect 110604 472806 110656 472812
rect 109224 471368 109276 471374
rect 109224 471310 109276 471316
rect 109132 471300 109184 471306
rect 109132 471242 109184 471248
rect 112640 470594 112668 488022
rect 113272 483404 113324 483410
rect 113272 483346 113324 483352
rect 113284 474162 113312 483346
rect 113468 480298 113496 488036
rect 113560 488022 113942 488050
rect 113560 483410 113588 488022
rect 113548 483404 113600 483410
rect 113548 483346 113600 483352
rect 114296 481030 114324 488036
rect 114284 481024 114336 481030
rect 114284 480966 114336 480972
rect 113376 480270 113496 480298
rect 113272 474156 113324 474162
rect 113272 474098 113324 474104
rect 113376 471442 113404 480270
rect 113364 471436 113416 471442
rect 113364 471378 113416 471384
rect 111996 470566 112668 470594
rect 111996 469878 112024 470566
rect 111984 469872 112036 469878
rect 111984 469814 112036 469820
rect 109040 468716 109092 468722
rect 109040 468658 109092 468664
rect 107844 468580 107896 468586
rect 107844 468522 107896 468528
rect 107660 468512 107712 468518
rect 107660 468454 107712 468460
rect 114756 467226 114784 488036
rect 115216 482662 115244 488036
rect 115204 482656 115256 482662
rect 115204 482598 115256 482604
rect 115676 482458 115704 488036
rect 115952 488022 116058 488050
rect 116136 488022 116518 488050
rect 116688 488022 116978 488050
rect 117332 488022 117438 488050
rect 117516 488022 117898 488050
rect 117976 488022 118266 488050
rect 118742 488022 118832 488050
rect 115664 482452 115716 482458
rect 115664 482394 115716 482400
rect 115952 479330 115980 488022
rect 116032 484152 116084 484158
rect 116032 484094 116084 484100
rect 116044 479466 116072 484094
rect 116032 479460 116084 479466
rect 116032 479402 116084 479408
rect 116136 479398 116164 488022
rect 116584 485172 116636 485178
rect 116584 485114 116636 485120
rect 116124 479392 116176 479398
rect 116124 479334 116176 479340
rect 115940 479324 115992 479330
rect 115940 479266 115992 479272
rect 116596 469878 116624 485114
rect 116688 484158 116716 488022
rect 116676 484152 116728 484158
rect 116676 484094 116728 484100
rect 117332 483750 117360 488022
rect 117516 484106 117544 488022
rect 117424 484078 117544 484106
rect 117320 483744 117372 483750
rect 117320 483686 117372 483692
rect 117424 480010 117452 484078
rect 117976 480078 118004 488022
rect 117964 480072 118016 480078
rect 117964 480014 118016 480020
rect 117412 480004 117464 480010
rect 117412 479946 117464 479952
rect 118804 479777 118832 488022
rect 118896 488022 119186 488050
rect 118896 480146 118924 488022
rect 119632 482390 119660 488036
rect 120092 482633 120120 488036
rect 120078 482624 120134 482633
rect 120078 482559 120134 482568
rect 120460 482497 120488 488036
rect 120552 488022 120934 488050
rect 120446 482488 120502 482497
rect 120446 482423 120502 482432
rect 119620 482384 119672 482390
rect 119620 482326 119672 482332
rect 118884 480140 118936 480146
rect 118884 480082 118936 480088
rect 118790 479768 118846 479777
rect 118790 479703 118846 479712
rect 120552 477358 120580 488022
rect 121380 482769 121408 488036
rect 121564 488022 121854 488050
rect 121932 488022 122222 488050
rect 122392 488022 122682 488050
rect 123036 488022 123142 488050
rect 123312 488022 123602 488050
rect 123680 488022 124062 488050
rect 121366 482760 121422 482769
rect 121366 482695 121422 482704
rect 120540 477352 120592 477358
rect 120540 477294 120592 477300
rect 121564 477222 121592 488022
rect 121932 479505 121960 488022
rect 121918 479496 121974 479505
rect 121918 479431 121974 479440
rect 121552 477216 121604 477222
rect 121552 477158 121604 477164
rect 122392 476114 122420 488022
rect 123036 479738 123064 488022
rect 123024 479732 123076 479738
rect 123024 479674 123076 479680
rect 123312 477290 123340 488022
rect 123300 477284 123352 477290
rect 123300 477226 123352 477232
rect 123680 476921 123708 488022
rect 124416 482361 124444 488036
rect 124508 488022 124890 488050
rect 124968 488022 125350 488050
rect 125612 488022 125810 488050
rect 125888 488022 126270 488050
rect 126348 488022 126638 488050
rect 127114 488022 127204 488050
rect 124402 482352 124458 482361
rect 124402 482287 124458 482296
rect 124508 479641 124536 488022
rect 124494 479632 124550 479641
rect 124494 479567 124550 479576
rect 124968 477154 124996 488022
rect 125612 477494 125640 488022
rect 125600 477488 125652 477494
rect 125600 477430 125652 477436
rect 124956 477148 125008 477154
rect 124956 477090 125008 477096
rect 125888 477086 125916 488022
rect 125876 477080 125928 477086
rect 125876 477022 125928 477028
rect 123666 476912 123722 476921
rect 123666 476847 123722 476856
rect 126348 476785 126376 488022
rect 127176 482118 127204 488022
rect 127268 488022 127558 488050
rect 127728 488022 128018 488050
rect 128494 488022 128584 488050
rect 127164 482112 127216 482118
rect 127164 482054 127216 482060
rect 126980 480888 127032 480894
rect 126980 480830 127032 480836
rect 126334 476776 126390 476785
rect 126334 476711 126390 476720
rect 121472 476086 122420 476114
rect 116584 469872 116636 469878
rect 116584 469814 116636 469820
rect 114744 467220 114796 467226
rect 114744 467162 114796 467168
rect 106280 467152 106332 467158
rect 106280 467094 106332 467100
rect 100852 465792 100904 465798
rect 100852 465734 100904 465740
rect 100760 464704 100812 464710
rect 100760 464646 100812 464652
rect 121472 464642 121500 476086
rect 126992 464642 127020 480830
rect 127268 473354 127296 488022
rect 127348 482112 127400 482118
rect 127348 482054 127400 482060
rect 127360 474201 127388 482054
rect 127728 480894 127756 488022
rect 128360 487076 128412 487082
rect 128360 487018 128412 487024
rect 127716 480888 127768 480894
rect 127716 480830 127768 480836
rect 128372 476678 128400 487018
rect 128556 485774 128584 488022
rect 128648 488022 128846 488050
rect 128924 488022 129306 488050
rect 129782 488022 129964 488050
rect 128648 487082 128676 488022
rect 128636 487076 128688 487082
rect 128636 487018 128688 487024
rect 128556 485746 128676 485774
rect 128648 476746 128676 485746
rect 128924 479534 128952 488022
rect 129936 479602 129964 488022
rect 130028 488022 130226 488050
rect 130304 488022 130594 488050
rect 130672 488022 131054 488050
rect 131132 488022 131514 488050
rect 131592 488022 131974 488050
rect 132052 488022 132434 488050
rect 129924 479596 129976 479602
rect 129924 479538 129976 479544
rect 128912 479528 128964 479534
rect 128912 479470 128964 479476
rect 128636 476740 128688 476746
rect 128636 476682 128688 476688
rect 128360 476672 128412 476678
rect 128360 476614 128412 476620
rect 127346 474192 127402 474201
rect 127346 474127 127402 474136
rect 127084 473326 127296 473354
rect 127084 464710 127112 473326
rect 127072 464704 127124 464710
rect 127072 464646 127124 464652
rect 121460 464636 121512 464642
rect 121460 464578 121512 464584
rect 126980 464636 127032 464642
rect 126980 464578 127032 464584
rect 130028 464574 130056 488022
rect 130304 480214 130332 488022
rect 130292 480208 130344 480214
rect 130292 480150 130344 480156
rect 130672 479670 130700 488022
rect 131132 482322 131160 488022
rect 131120 482316 131172 482322
rect 131120 482258 131172 482264
rect 131592 479874 131620 488022
rect 131580 479868 131632 479874
rect 131580 479810 131632 479816
rect 130660 479664 130712 479670
rect 130660 479606 130712 479612
rect 132052 470594 132080 488022
rect 132788 479942 132816 488036
rect 132880 488022 133262 488050
rect 133432 488022 133722 488050
rect 133892 488022 134182 488050
rect 134260 488022 134642 488050
rect 134720 488022 135010 488050
rect 135272 488022 135470 488050
rect 135946 488022 136312 488050
rect 136406 488022 136588 488050
rect 132776 479936 132828 479942
rect 132776 479878 132828 479884
rect 132880 476950 132908 488022
rect 133432 477018 133460 488022
rect 133420 477012 133472 477018
rect 133420 476954 133472 476960
rect 132868 476944 132920 476950
rect 132868 476886 132920 476892
rect 131316 470566 132080 470594
rect 130016 464568 130068 464574
rect 130016 464510 130068 464516
rect 131316 464506 131344 470566
rect 131304 464500 131356 464506
rect 131304 464442 131356 464448
rect 133892 464370 133920 488022
rect 134260 476114 134288 488022
rect 134720 477426 134748 488022
rect 135272 479806 135300 488022
rect 136284 482322 136312 488022
rect 136560 482390 136588 488022
rect 136652 488022 136758 488050
rect 136548 482384 136600 482390
rect 136548 482326 136600 482332
rect 136272 482316 136324 482322
rect 136272 482258 136324 482264
rect 135260 479800 135312 479806
rect 135260 479742 135312 479748
rect 134708 477420 134760 477426
rect 134708 477362 134760 477368
rect 133984 476086 134288 476114
rect 133984 464438 134012 476086
rect 136652 464438 136680 488022
rect 137204 482526 137232 488036
rect 137296 488022 137678 488050
rect 138154 488022 138520 488050
rect 138614 488022 138888 488050
rect 138982 488022 139256 488050
rect 137192 482520 137244 482526
rect 137192 482462 137244 482468
rect 137296 470594 137324 488022
rect 138492 482594 138520 488022
rect 138480 482588 138532 482594
rect 138480 482530 138532 482536
rect 138860 482458 138888 488022
rect 139228 485178 139256 488022
rect 139216 485172 139268 485178
rect 139216 485114 139268 485120
rect 139412 485042 139440 488036
rect 139504 488022 139886 488050
rect 140056 488022 140346 488050
rect 140822 488022 140912 488050
rect 139400 485036 139452 485042
rect 139400 484978 139452 484984
rect 139400 484152 139452 484158
rect 139400 484094 139452 484100
rect 138848 482452 138900 482458
rect 138848 482394 138900 482400
rect 139412 471646 139440 484094
rect 139504 474094 139532 488022
rect 140056 484158 140084 488022
rect 140884 486538 140912 488022
rect 140976 488022 141174 488050
rect 141344 488022 141634 488050
rect 141712 488022 142094 488050
rect 142356 488022 142554 488050
rect 142632 488022 142922 488050
rect 143000 488022 143382 488050
rect 143644 488022 143842 488050
rect 143920 488022 144302 488050
rect 144778 488022 144868 488050
rect 145146 488022 145512 488050
rect 145606 488022 145696 488050
rect 140872 486532 140924 486538
rect 140872 486474 140924 486480
rect 140780 484220 140832 484226
rect 140780 484162 140832 484168
rect 140044 484152 140096 484158
rect 140044 484094 140096 484100
rect 139492 474088 139544 474094
rect 139492 474030 139544 474036
rect 139400 471640 139452 471646
rect 139400 471582 139452 471588
rect 136744 470566 137324 470594
rect 133972 464432 134024 464438
rect 133972 464374 134024 464380
rect 136640 464432 136692 464438
rect 136640 464374 136692 464380
rect 136744 464370 136772 470566
rect 140792 465798 140820 484162
rect 140872 484152 140924 484158
rect 140872 484094 140924 484100
rect 140884 471510 140912 484094
rect 140976 471578 141004 488022
rect 141344 484158 141372 488022
rect 141712 484226 141740 488022
rect 141700 484220 141752 484226
rect 141700 484162 141752 484168
rect 142252 484220 142304 484226
rect 142252 484162 142304 484168
rect 141332 484152 141384 484158
rect 141332 484094 141384 484100
rect 142160 484152 142212 484158
rect 142160 484094 142212 484100
rect 140964 471572 141016 471578
rect 140964 471514 141016 471520
rect 140872 471504 140924 471510
rect 140872 471446 140924 471452
rect 142172 466002 142200 484094
rect 142160 465996 142212 466002
rect 142160 465938 142212 465944
rect 142264 465934 142292 484162
rect 142356 471442 142384 488022
rect 142632 484158 142660 488022
rect 143000 484226 143028 488022
rect 142988 484220 143040 484226
rect 142988 484162 143040 484168
rect 142620 484152 142672 484158
rect 142620 484094 142672 484100
rect 143540 484152 143592 484158
rect 143540 484094 143592 484100
rect 143552 474065 143580 484094
rect 143644 476882 143672 488022
rect 143920 484158 143948 488022
rect 143908 484152 143960 484158
rect 143908 484094 143960 484100
rect 144840 483721 144868 488022
rect 145484 485081 145512 488022
rect 145668 485353 145696 488022
rect 145760 488022 146050 488050
rect 146312 488022 146510 488050
rect 146986 488022 147260 488050
rect 147354 488022 147628 488050
rect 147814 488022 148088 488050
rect 145654 485344 145710 485353
rect 145654 485279 145710 485288
rect 145470 485072 145526 485081
rect 145470 485007 145526 485016
rect 144826 483712 144882 483721
rect 144826 483647 144882 483656
rect 145760 478417 145788 488022
rect 145746 478408 145802 478417
rect 145746 478343 145802 478352
rect 143632 476876 143684 476882
rect 143632 476818 143684 476824
rect 143538 474056 143594 474065
rect 143538 473991 143594 474000
rect 142344 471436 142396 471442
rect 142344 471378 142396 471384
rect 146312 467158 146340 488022
rect 147232 480865 147260 488022
rect 147600 485217 147628 488022
rect 147586 485208 147642 485217
rect 147586 485143 147642 485152
rect 148060 482361 148088 488022
rect 148244 485489 148272 488036
rect 148336 488022 148718 488050
rect 149194 488022 149468 488050
rect 148230 485480 148286 485489
rect 148230 485415 148286 485424
rect 148046 482352 148102 482361
rect 148046 482287 148102 482296
rect 147218 480856 147274 480865
rect 147218 480791 147274 480800
rect 148336 479505 148364 488022
rect 149440 485450 149468 488022
rect 149532 485654 149560 488036
rect 149624 488022 150006 488050
rect 149520 485648 149572 485654
rect 149520 485590 149572 485596
rect 149428 485444 149480 485450
rect 149428 485386 149480 485392
rect 148322 479496 148378 479505
rect 148322 479431 148378 479440
rect 149624 470594 149652 488022
rect 150452 485722 150480 488036
rect 150544 488022 150926 488050
rect 150440 485716 150492 485722
rect 150440 485658 150492 485664
rect 150544 484106 150572 488022
rect 151280 485586 151308 488036
rect 151372 488022 151754 488050
rect 151268 485580 151320 485586
rect 151268 485522 151320 485528
rect 150452 484078 150572 484106
rect 150452 476882 150480 484078
rect 151372 478281 151400 488022
rect 152200 485790 152228 488036
rect 152292 488022 152674 488050
rect 152752 488022 153134 488050
rect 153212 488022 153502 488050
rect 153978 488022 154344 488050
rect 154438 488022 154528 488050
rect 152188 485784 152240 485790
rect 152188 485726 152240 485732
rect 152292 484106 152320 488022
rect 151832 484078 152320 484106
rect 151358 478272 151414 478281
rect 151358 478207 151414 478216
rect 150440 476876 150492 476882
rect 150440 476818 150492 476824
rect 149072 470566 149652 470594
rect 149072 467226 149100 470566
rect 149060 467220 149112 467226
rect 149060 467162 149112 467168
rect 146300 467152 146352 467158
rect 151832 467129 151860 484078
rect 152752 472569 152780 488022
rect 153212 474337 153240 488022
rect 154316 485246 154344 488022
rect 154304 485240 154356 485246
rect 154304 485182 154356 485188
rect 154500 482497 154528 488022
rect 154684 488022 154882 488050
rect 154580 484152 154632 484158
rect 154580 484094 154632 484100
rect 154486 482488 154542 482497
rect 154486 482423 154542 482432
rect 153198 474328 153254 474337
rect 153198 474263 153254 474272
rect 152738 472560 152794 472569
rect 152738 472495 152794 472504
rect 154592 467265 154620 484094
rect 154684 479641 154712 488022
rect 155328 484838 155356 488036
rect 155420 488022 155710 488050
rect 156186 488022 156552 488050
rect 156646 488022 156736 488050
rect 155316 484832 155368 484838
rect 155316 484774 155368 484780
rect 155420 484158 155448 488022
rect 155408 484152 155460 484158
rect 155408 484094 155460 484100
rect 156524 483857 156552 488022
rect 156708 485314 156736 488022
rect 156800 488022 157090 488050
rect 156696 485308 156748 485314
rect 156696 485250 156748 485256
rect 156510 483848 156566 483857
rect 156510 483783 156566 483792
rect 154670 479632 154726 479641
rect 154670 479567 154726 479576
rect 156800 475561 156828 488022
rect 157444 485382 157472 488036
rect 157536 488022 157918 488050
rect 158394 488022 158668 488050
rect 158854 488022 158944 488050
rect 157432 485376 157484 485382
rect 157432 485318 157484 485324
rect 157536 476785 157564 488022
rect 157708 485512 157760 485518
rect 157708 485454 157760 485460
rect 157720 485314 157748 485454
rect 157708 485308 157760 485314
rect 157708 485250 157760 485256
rect 157800 485308 157852 485314
rect 157800 485250 157852 485256
rect 157812 484838 157840 485250
rect 158640 484974 158668 488022
rect 158628 484968 158680 484974
rect 158628 484910 158680 484916
rect 157800 484832 157852 484838
rect 157800 484774 157852 484780
rect 158720 481024 158772 481030
rect 158720 480966 158772 480972
rect 157522 476776 157578 476785
rect 157522 476711 157578 476720
rect 156786 475552 156842 475561
rect 156786 475487 156842 475496
rect 154578 467256 154634 467265
rect 154578 467191 154634 467200
rect 146300 467094 146352 467100
rect 151818 467120 151874 467129
rect 151818 467055 151874 467064
rect 142252 465928 142304 465934
rect 142252 465870 142304 465876
rect 158732 465866 158760 480966
rect 158812 480888 158864 480894
rect 158812 480830 158864 480836
rect 158824 468858 158852 480830
rect 158916 474230 158944 488022
rect 159008 488022 159298 488050
rect 159376 488022 159666 488050
rect 159008 480894 159036 488022
rect 159376 481030 159404 488022
rect 160128 487778 160156 488036
rect 160388 488022 160586 488050
rect 160664 488022 161046 488050
rect 160128 487750 160324 487778
rect 160296 481030 160324 487750
rect 159364 481024 159416 481030
rect 159364 480966 159416 480972
rect 160284 481024 160336 481030
rect 160284 480966 160336 480972
rect 158996 480888 159048 480894
rect 158996 480830 159048 480836
rect 160100 480888 160152 480894
rect 160100 480830 160152 480836
rect 158904 474224 158956 474230
rect 158904 474166 158956 474172
rect 160112 469849 160140 480830
rect 160388 472666 160416 488022
rect 160664 480894 160692 488022
rect 160652 480888 160704 480894
rect 160652 480830 160704 480836
rect 160376 472660 160428 472666
rect 160376 472602 160428 472608
rect 160098 469840 160154 469849
rect 160098 469775 160154 469784
rect 158812 468852 158864 468858
rect 158812 468794 158864 468800
rect 161492 468790 161520 488036
rect 161572 480888 161624 480894
rect 161572 480830 161624 480836
rect 161584 471345 161612 480830
rect 161664 479800 161716 479806
rect 161664 479742 161716 479748
rect 161676 475697 161704 479742
rect 161860 476114 161888 488036
rect 161952 488022 162334 488050
rect 162504 488022 162794 488050
rect 163056 488022 163254 488050
rect 163332 488022 163622 488050
rect 163792 488022 164082 488050
rect 161952 479806 161980 488022
rect 162504 480894 162532 488022
rect 162492 480888 162544 480894
rect 162492 480830 162544 480836
rect 161940 479800 161992 479806
rect 161940 479742 161992 479748
rect 163056 479534 163084 488022
rect 163044 479528 163096 479534
rect 163044 479470 163096 479476
rect 163332 476114 163360 488022
rect 163792 476921 163820 488022
rect 164528 484265 164556 488036
rect 164620 488022 165002 488050
rect 165080 488022 165462 488050
rect 165632 488022 165830 488050
rect 166092 488022 166290 488050
rect 166368 488022 166750 488050
rect 167012 488022 167210 488050
rect 167288 488022 167670 488050
rect 167748 488022 168038 488050
rect 168392 488022 168498 488050
rect 168576 488022 168958 488050
rect 169036 488022 169418 488050
rect 169772 488022 169878 488050
rect 169956 488022 170246 488050
rect 170416 488022 170706 488050
rect 164514 484256 164570 484265
rect 164514 484191 164570 484200
rect 163778 476912 163834 476921
rect 163778 476847 163834 476856
rect 164620 476114 164648 488022
rect 165080 478242 165108 488022
rect 165068 478236 165120 478242
rect 165068 478178 165120 478184
rect 161768 476086 161888 476114
rect 162872 476086 163360 476114
rect 164252 476086 164648 476114
rect 161662 475688 161718 475697
rect 161662 475623 161718 475632
rect 161570 471336 161626 471345
rect 161570 471271 161626 471280
rect 161768 471209 161796 476086
rect 162872 471481 162900 476086
rect 164252 475386 164280 476086
rect 164240 475380 164292 475386
rect 164240 475322 164292 475328
rect 162858 471472 162914 471481
rect 162858 471407 162914 471416
rect 161754 471200 161810 471209
rect 161754 471135 161810 471144
rect 161480 468784 161532 468790
rect 161480 468726 161532 468732
rect 158720 465860 158772 465866
rect 158720 465802 158772 465808
rect 140780 465792 140832 465798
rect 165632 465769 165660 488022
rect 166092 484770 166120 488022
rect 166080 484764 166132 484770
rect 166080 484706 166132 484712
rect 166368 470594 166396 488022
rect 165816 470566 166396 470594
rect 165816 465905 165844 470566
rect 167012 466041 167040 488022
rect 167092 484152 167144 484158
rect 167092 484094 167144 484100
rect 167104 468625 167132 484094
rect 167288 468897 167316 488022
rect 167748 484158 167776 488022
rect 167736 484152 167788 484158
rect 167736 484094 167788 484100
rect 167274 468888 167330 468897
rect 167274 468823 167330 468832
rect 168392 468761 168420 488022
rect 168576 484140 168604 488022
rect 168484 484112 168604 484140
rect 168484 474162 168512 484112
rect 168472 474156 168524 474162
rect 168472 474098 168524 474104
rect 169036 470594 169064 488022
rect 168576 470566 169064 470594
rect 168378 468752 168434 468761
rect 168378 468687 168434 468696
rect 167090 468616 167146 468625
rect 167090 468551 167146 468560
rect 168576 468489 168604 470566
rect 169772 469033 169800 488022
rect 169852 484152 169904 484158
rect 169852 484094 169904 484100
rect 169864 469985 169892 484094
rect 169956 472734 169984 488022
rect 170416 484158 170444 488022
rect 171152 485625 171180 488036
rect 171244 488022 171626 488050
rect 171704 488022 171994 488050
rect 172072 488022 172454 488050
rect 172624 488022 172914 488050
rect 173390 488022 173480 488050
rect 171138 485616 171194 485625
rect 171138 485551 171194 485560
rect 170404 484152 170456 484158
rect 170404 484094 170456 484100
rect 171140 484152 171192 484158
rect 171140 484094 171192 484100
rect 169944 472728 169996 472734
rect 169944 472670 169996 472676
rect 169850 469976 169906 469985
rect 169850 469911 169906 469920
rect 169758 469024 169814 469033
rect 169758 468959 169814 468968
rect 168562 468480 168618 468489
rect 168562 468415 168618 468424
rect 166998 466032 167054 466041
rect 166998 465967 167054 465976
rect 165802 465896 165858 465905
rect 165802 465831 165858 465840
rect 140780 465734 140832 465740
rect 165618 465760 165674 465769
rect 165618 465695 165674 465704
rect 171152 464409 171180 484094
rect 171244 472705 171272 488022
rect 171704 484158 171732 488022
rect 171692 484152 171744 484158
rect 171692 484094 171744 484100
rect 172072 479777 172100 488022
rect 172520 484152 172572 484158
rect 172520 484094 172572 484100
rect 172058 479768 172114 479777
rect 172058 479703 172114 479712
rect 171230 472696 171286 472705
rect 171230 472631 171286 472640
rect 172532 467362 172560 484094
rect 172624 471617 172652 488022
rect 173452 482662 173480 488022
rect 173544 488022 173834 488050
rect 173912 488022 174202 488050
rect 174280 488022 174662 488050
rect 174832 488022 175122 488050
rect 175384 488022 175582 488050
rect 173544 484158 173572 488022
rect 173532 484152 173584 484158
rect 173532 484094 173584 484100
rect 173440 482656 173492 482662
rect 173440 482598 173492 482604
rect 172610 471608 172666 471617
rect 172610 471543 172666 471552
rect 172520 467356 172572 467362
rect 172520 467298 172572 467304
rect 173912 466138 173940 488022
rect 174280 484106 174308 488022
rect 174004 484078 174308 484106
rect 173900 466132 173952 466138
rect 173900 466074 173952 466080
rect 174004 466070 174032 484078
rect 174832 471850 174860 488022
rect 175280 484152 175332 484158
rect 175280 484094 175332 484100
rect 174820 471844 174872 471850
rect 174820 471786 174872 471792
rect 175292 468926 175320 484094
rect 175384 472802 175412 488022
rect 176028 482730 176056 488036
rect 176120 488022 176410 488050
rect 176886 488022 176976 488050
rect 176120 484158 176148 488022
rect 176108 484152 176160 484158
rect 176108 484094 176160 484100
rect 176948 483750 176976 488022
rect 177040 488022 177330 488050
rect 177408 488022 177790 488050
rect 178174 488022 178264 488050
rect 176936 483744 176988 483750
rect 176936 483686 176988 483692
rect 176016 482724 176068 482730
rect 176016 482666 176068 482672
rect 177040 478310 177068 488022
rect 177028 478304 177080 478310
rect 177028 478246 177080 478252
rect 177408 476114 177436 488022
rect 178040 487076 178092 487082
rect 178040 487018 178092 487024
rect 176672 476086 177436 476114
rect 176672 475454 176700 476086
rect 176660 475448 176712 475454
rect 176660 475390 176712 475396
rect 175372 472796 175424 472802
rect 175372 472738 175424 472744
rect 178052 470014 178080 487018
rect 178236 485774 178264 488022
rect 178328 488022 178618 488050
rect 179094 488022 179368 488050
rect 178328 487082 178356 488022
rect 178316 487076 178368 487082
rect 178316 487018 178368 487024
rect 178236 485746 178356 485774
rect 178328 479602 178356 485746
rect 179340 481001 179368 488022
rect 179326 480992 179382 481001
rect 179326 480927 179382 480936
rect 179420 480888 179472 480894
rect 179420 480830 179472 480836
rect 178316 479596 178368 479602
rect 178316 479538 178368 479544
rect 178040 470008 178092 470014
rect 178040 469950 178092 469956
rect 179432 469946 179460 480830
rect 179524 474298 179552 488036
rect 179616 488022 179998 488050
rect 180382 488022 180564 488050
rect 180842 488022 180932 488050
rect 179616 480894 179644 488022
rect 180064 485104 180116 485110
rect 180064 485046 180116 485052
rect 179604 480888 179656 480894
rect 179604 480830 179656 480836
rect 179512 474292 179564 474298
rect 179512 474234 179564 474240
rect 179420 469940 179472 469946
rect 179420 469882 179472 469888
rect 175280 468920 175332 468926
rect 175280 468862 175332 468868
rect 178040 467832 178092 467838
rect 178040 467774 178092 467780
rect 178052 466614 178080 467774
rect 178040 466608 178092 466614
rect 178038 466576 178040 466585
rect 178092 466576 178094 466585
rect 178038 466511 178094 466520
rect 180076 466177 180104 485046
rect 180536 481098 180564 488022
rect 180904 481166 180932 488022
rect 180996 488022 181286 488050
rect 181456 488022 181746 488050
rect 182222 488022 182404 488050
rect 180892 481160 180944 481166
rect 180892 481102 180944 481108
rect 180524 481092 180576 481098
rect 180524 481034 180576 481040
rect 180996 478122 181024 488022
rect 181076 481160 181128 481166
rect 181076 481102 181128 481108
rect 180812 478094 181024 478122
rect 180156 474020 180208 474026
rect 180156 473962 180208 473968
rect 180168 467294 180196 473962
rect 180156 467288 180208 467294
rect 180156 467230 180208 467236
rect 180168 466993 180196 467230
rect 180154 466984 180210 466993
rect 180154 466919 180210 466928
rect 180062 466168 180118 466177
rect 180062 466103 180118 466112
rect 173992 466064 174044 466070
rect 173992 466006 174044 466012
rect 180812 464574 180840 478094
rect 181088 473354 181116 481102
rect 180904 473326 181116 473354
rect 180904 466206 180932 473326
rect 181456 470594 181484 488022
rect 182376 481370 182404 488022
rect 182468 488022 182574 488050
rect 182744 488022 183034 488050
rect 183112 488022 183494 488050
rect 183756 488022 183954 488050
rect 184032 488022 184322 488050
rect 184400 488022 184782 488050
rect 185044 488022 185242 488050
rect 185718 488022 185808 488050
rect 182364 481364 182416 481370
rect 182364 481306 182416 481312
rect 182364 481160 182416 481166
rect 182364 481102 182416 481108
rect 182272 480888 182324 480894
rect 182272 480830 182324 480836
rect 182180 474836 182232 474842
rect 182180 474778 182232 474784
rect 180996 470566 181484 470594
rect 180996 468994 181024 470566
rect 180984 468988 181036 468994
rect 180984 468930 181036 468936
rect 182192 468382 182220 474778
rect 182284 471986 182312 480830
rect 182272 471980 182324 471986
rect 182272 471922 182324 471928
rect 182376 471782 182404 481102
rect 182468 474842 182496 488022
rect 182456 474836 182508 474842
rect 182456 474778 182508 474784
rect 182744 471889 182772 488022
rect 183112 480894 183140 488022
rect 183100 480888 183152 480894
rect 183100 480830 183152 480836
rect 183652 480888 183704 480894
rect 183652 480830 183704 480836
rect 183560 480820 183612 480826
rect 183560 480762 183612 480768
rect 182730 471880 182786 471889
rect 182730 471815 182786 471824
rect 182364 471776 182416 471782
rect 182364 471718 182416 471724
rect 182180 468376 182232 468382
rect 182180 468318 182232 468324
rect 183572 466342 183600 480762
rect 183664 471753 183692 480830
rect 183650 471744 183706 471753
rect 183756 471714 183784 488022
rect 184032 480894 184060 488022
rect 184020 480888 184072 480894
rect 184020 480830 184072 480836
rect 184400 480826 184428 488022
rect 184940 480888 184992 480894
rect 184940 480830 184992 480836
rect 184388 480820 184440 480826
rect 184388 480762 184440 480768
rect 183650 471679 183706 471688
rect 183744 471708 183796 471714
rect 183744 471650 183796 471656
rect 184952 467430 184980 480830
rect 185044 476950 185072 488022
rect 185584 485036 185636 485042
rect 185584 484978 185636 484984
rect 185032 476944 185084 476950
rect 185032 476886 185084 476892
rect 185596 474026 185624 484978
rect 185780 484945 185808 488022
rect 185872 488022 186162 488050
rect 186424 488022 186530 488050
rect 187006 488022 187096 488050
rect 185766 484936 185822 484945
rect 185766 484871 185822 484880
rect 185872 480894 185900 488022
rect 185860 480888 185912 480894
rect 185860 480830 185912 480836
rect 186424 478378 186452 488022
rect 187068 485761 187096 488022
rect 187160 488022 187450 488050
rect 187804 488022 187910 488050
rect 188080 488022 188370 488050
rect 188448 488022 188738 488050
rect 187054 485752 187110 485761
rect 187054 485687 187110 485696
rect 186412 478372 186464 478378
rect 186412 478314 186464 478320
rect 187160 476114 187188 488022
rect 187700 480888 187752 480894
rect 187700 480830 187752 480836
rect 186332 476086 187188 476114
rect 185584 474020 185636 474026
rect 185584 473962 185636 473968
rect 184940 467424 184992 467430
rect 184940 467366 184992 467372
rect 183560 466336 183612 466342
rect 183560 466278 183612 466284
rect 180892 466200 180944 466206
rect 180892 466142 180944 466148
rect 180800 464568 180852 464574
rect 180800 464510 180852 464516
rect 186332 464506 186360 476086
rect 187712 465594 187740 480830
rect 187804 466410 187832 488022
rect 188080 474366 188108 488022
rect 188344 485376 188396 485382
rect 188344 485318 188396 485324
rect 188356 485178 188384 485318
rect 188344 485172 188396 485178
rect 188344 485114 188396 485120
rect 188448 480894 188476 488022
rect 189200 487778 189228 488036
rect 189460 488022 189658 488050
rect 189736 488022 190118 488050
rect 189200 487750 189396 487778
rect 189264 485308 189316 485314
rect 189264 485250 189316 485256
rect 189276 485042 189304 485250
rect 189264 485036 189316 485042
rect 189264 484978 189316 484984
rect 189368 481166 189396 487750
rect 189356 481160 189408 481166
rect 189356 481102 189408 481108
rect 188436 480888 188488 480894
rect 188436 480830 188488 480836
rect 189460 476114 189488 488022
rect 189092 476086 189488 476114
rect 188068 474360 188120 474366
rect 188068 474302 188120 474308
rect 189092 467498 189120 476086
rect 189736 470594 189764 488022
rect 189184 470566 189764 470594
rect 189184 469062 189212 470566
rect 189172 469056 189224 469062
rect 189172 468998 189224 469004
rect 189080 467492 189132 467498
rect 189080 467434 189132 467440
rect 187792 466404 187844 466410
rect 187792 466346 187844 466352
rect 187700 465588 187752 465594
rect 187700 465530 187752 465536
rect 190472 464778 190500 488036
rect 190656 488022 190946 488050
rect 191024 488022 191406 488050
rect 191882 488022 192156 488050
rect 190552 479732 190604 479738
rect 190552 479674 190604 479680
rect 190564 471170 190592 479674
rect 190656 471918 190684 488022
rect 191024 479738 191052 488022
rect 191196 485444 191248 485450
rect 191196 485386 191248 485392
rect 191208 485178 191236 485386
rect 191196 485172 191248 485178
rect 191196 485114 191248 485120
rect 192128 481234 192156 488022
rect 192220 488022 192326 488050
rect 192404 488022 192694 488050
rect 192864 488022 193154 488050
rect 193416 488022 193614 488050
rect 193784 488022 194074 488050
rect 194152 488022 194534 488050
rect 194918 488022 195192 488050
rect 192116 481228 192168 481234
rect 192116 481170 192168 481176
rect 192220 481114 192248 488022
rect 192300 481228 192352 481234
rect 192300 481170 192352 481176
rect 191852 481086 192248 481114
rect 191012 479732 191064 479738
rect 191012 479674 191064 479680
rect 190644 471912 190696 471918
rect 190644 471854 190696 471860
rect 190552 471164 190604 471170
rect 190552 471106 190604 471112
rect 190918 466576 190974 466585
rect 190918 466511 190974 466520
rect 190932 466478 190960 466511
rect 190920 466472 190972 466478
rect 190920 466414 190972 466420
rect 191852 464846 191880 481086
rect 191932 480888 191984 480894
rect 191932 480830 191984 480836
rect 191944 469130 191972 480830
rect 192024 480820 192076 480826
rect 192024 480762 192076 480768
rect 191932 469124 191984 469130
rect 191932 469066 191984 469072
rect 192036 468450 192064 480762
rect 192312 471238 192340 481170
rect 192404 480894 192432 488022
rect 192392 480888 192444 480894
rect 192392 480830 192444 480836
rect 192864 480826 192892 488022
rect 193312 480888 193364 480894
rect 193312 480830 193364 480836
rect 192852 480820 192904 480826
rect 192852 480762 192904 480768
rect 193220 480820 193272 480826
rect 193220 480762 193272 480768
rect 192300 471232 192352 471238
rect 192300 471174 192352 471180
rect 192024 468444 192076 468450
rect 192024 468386 192076 468392
rect 193232 466274 193260 480762
rect 193220 466268 193272 466274
rect 193220 466210 193272 466216
rect 193324 465526 193352 480830
rect 193416 469198 193444 488022
rect 193784 480894 193812 488022
rect 193864 485104 193916 485110
rect 193864 485046 193916 485052
rect 193772 480888 193824 480894
rect 193772 480830 193824 480836
rect 193876 470694 193904 485046
rect 194152 480826 194180 488022
rect 195164 484430 195192 488022
rect 195348 485110 195376 488036
rect 195440 488022 195822 488050
rect 196298 488022 196664 488050
rect 195336 485104 195388 485110
rect 195336 485046 195388 485052
rect 195152 484424 195204 484430
rect 195152 484366 195204 484372
rect 194140 480820 194192 480826
rect 194140 480762 194192 480768
rect 193864 470688 193916 470694
rect 193864 470630 193916 470636
rect 195440 470594 195468 488022
rect 194612 470566 195468 470594
rect 193404 469192 193456 469198
rect 193404 469134 193456 469140
rect 194612 465662 194640 470566
rect 194600 465656 194652 465662
rect 194600 465598 194652 465604
rect 193312 465520 193364 465526
rect 193312 465462 193364 465468
rect 191840 464840 191892 464846
rect 191840 464782 191892 464788
rect 190460 464772 190512 464778
rect 190460 464714 190512 464720
rect 186320 464500 186372 464506
rect 186320 464442 186372 464448
rect 171138 464400 171194 464409
rect 133880 464364 133932 464370
rect 133880 464306 133932 464312
rect 136732 464364 136784 464370
rect 171138 464335 171194 464344
rect 136732 464306 136784 464312
rect 60740 380928 60792 380934
rect 60740 380870 60792 380876
rect 60752 357406 60780 380870
rect 155960 380656 156012 380662
rect 155960 380598 156012 380604
rect 105820 380520 105872 380526
rect 105820 380462 105872 380468
rect 138480 380520 138532 380526
rect 138480 380462 138532 380468
rect 105832 380361 105860 380462
rect 118332 380452 118384 380458
rect 118332 380394 118384 380400
rect 135904 380452 135956 380458
rect 135904 380394 135956 380400
rect 113548 380384 113600 380390
rect 105818 380352 105874 380361
rect 105818 380287 105874 380296
rect 110970 380352 111026 380361
rect 110970 380287 110972 380296
rect 111024 380287 111026 380296
rect 113546 380352 113548 380361
rect 118344 380361 118372 380394
rect 123576 380384 123628 380390
rect 113600 380352 113602 380361
rect 113546 380287 113602 380296
rect 115938 380352 115994 380361
rect 115938 380287 115994 380296
rect 118330 380352 118386 380361
rect 118330 380287 118386 380296
rect 120906 380352 120962 380361
rect 120906 380287 120962 380296
rect 123574 380352 123576 380361
rect 135916 380361 135944 380394
rect 138492 380361 138520 380462
rect 155972 380361 156000 380598
rect 158536 380588 158588 380594
rect 158536 380530 158588 380536
rect 158548 380361 158576 380530
rect 123628 380352 123630 380361
rect 123574 380287 123630 380296
rect 128358 380352 128414 380361
rect 128358 380287 128414 380296
rect 133510 380352 133566 380361
rect 133510 380287 133566 380296
rect 135902 380352 135958 380361
rect 135902 380287 135958 380296
rect 138478 380352 138534 380361
rect 138478 380287 138534 380296
rect 148598 380352 148654 380361
rect 148598 380287 148600 380296
rect 110972 380258 111024 380264
rect 115952 380186 115980 380287
rect 120920 380254 120948 380287
rect 120908 380248 120960 380254
rect 120908 380190 120960 380196
rect 128372 380186 128400 380287
rect 133524 380254 133552 380287
rect 148652 380287 148654 380296
rect 155958 380352 156014 380361
rect 155958 380287 156014 380296
rect 158534 380352 158590 380361
rect 158534 380287 158590 380296
rect 160926 380352 160982 380361
rect 160926 380287 160982 380296
rect 163502 380352 163558 380361
rect 163502 380287 163558 380296
rect 166078 380352 166134 380361
rect 166078 380287 166134 380296
rect 148600 380258 148652 380264
rect 133512 380248 133564 380254
rect 133512 380190 133564 380196
rect 115940 380180 115992 380186
rect 115940 380122 115992 380128
rect 128360 380180 128412 380186
rect 128360 380122 128412 380128
rect 160940 380118 160968 380287
rect 160928 380112 160980 380118
rect 160928 380054 160980 380060
rect 163516 379982 163544 380287
rect 166092 380050 166120 380287
rect 166080 380044 166132 380050
rect 166080 379986 166132 379992
rect 163504 379976 163556 379982
rect 163504 379918 163556 379924
rect 86592 379500 86644 379506
rect 86592 379442 86644 379448
rect 86604 379409 86632 379442
rect 88340 379432 88392 379438
rect 80334 379400 80390 379409
rect 80334 379335 80390 379344
rect 85486 379400 85542 379409
rect 85486 379335 85542 379344
rect 86590 379400 86646 379409
rect 86590 379335 86646 379344
rect 87694 379400 87750 379409
rect 87694 379335 87750 379344
rect 88338 379400 88340 379409
rect 92388 379432 92440 379438
rect 88392 379400 88394 379409
rect 88338 379335 88394 379344
rect 88798 379400 88854 379409
rect 88798 379335 88800 379344
rect 77206 378992 77262 379001
rect 77206 378927 77262 378936
rect 77220 376718 77248 378927
rect 80348 378729 80376 379335
rect 81438 378856 81494 378865
rect 81438 378791 81494 378800
rect 80334 378720 80390 378729
rect 80334 378655 80390 378664
rect 80348 378214 80376 378655
rect 81452 378282 81480 378791
rect 85500 378622 85528 379335
rect 85488 378616 85540 378622
rect 85488 378558 85540 378564
rect 81440 378276 81492 378282
rect 81440 378218 81492 378224
rect 87708 378214 87736 379335
rect 88852 379335 88854 379344
rect 90638 379400 90694 379409
rect 90638 379335 90694 379344
rect 91374 379400 91430 379409
rect 91374 379335 91430 379344
rect 92386 379400 92388 379409
rect 92440 379400 92442 379409
rect 92386 379335 92442 379344
rect 93582 379400 93638 379409
rect 93582 379335 93638 379344
rect 96066 379400 96122 379409
rect 96066 379335 96122 379344
rect 98182 379400 98238 379409
rect 98182 379335 98238 379344
rect 101034 379400 101090 379409
rect 101034 379335 101090 379344
rect 103518 379400 103574 379409
rect 103518 379335 103574 379344
rect 105358 379400 105414 379409
rect 105358 379335 105414 379344
rect 108210 379400 108266 379409
rect 108210 379335 108266 379344
rect 108854 379400 108910 379409
rect 108854 379335 108910 379344
rect 111246 379400 111302 379409
rect 111246 379335 111302 379344
rect 112350 379400 112406 379409
rect 112350 379335 112406 379344
rect 113454 379400 113510 379409
rect 113454 379335 113510 379344
rect 114466 379400 114522 379409
rect 114466 379335 114522 379344
rect 115846 379400 115902 379409
rect 115846 379335 115902 379344
rect 141054 379400 141110 379409
rect 141054 379335 141110 379344
rect 143630 379400 143686 379409
rect 143630 379335 143686 379344
rect 146022 379400 146078 379409
rect 146022 379335 146078 379344
rect 150990 379400 151046 379409
rect 150990 379335 151046 379344
rect 153566 379400 153622 379409
rect 153566 379335 153622 379344
rect 88800 379306 88852 379312
rect 90652 379302 90680 379335
rect 90640 379296 90692 379302
rect 90732 379296 90784 379302
rect 90640 379238 90692 379244
rect 90730 379264 90732 379273
rect 90784 379264 90786 379273
rect 91388 379234 91416 379335
rect 93490 379264 93546 379273
rect 90730 379199 90786 379208
rect 91376 379228 91428 379234
rect 93490 379199 93546 379208
rect 91376 379170 91428 379176
rect 93504 379166 93532 379199
rect 93596 379166 93624 379335
rect 95974 379264 96030 379273
rect 95974 379199 96030 379208
rect 93492 379160 93544 379166
rect 93492 379102 93544 379108
rect 93584 379160 93636 379166
rect 93584 379102 93636 379108
rect 94686 378584 94742 378593
rect 94686 378519 94742 378528
rect 80336 378208 80388 378214
rect 80336 378150 80388 378156
rect 87696 378208 87748 378214
rect 87696 378150 87748 378156
rect 77208 376712 77260 376718
rect 77208 376654 77260 376660
rect 94700 376174 94728 378519
rect 95988 377913 96016 379199
rect 96080 378690 96108 379335
rect 98196 378894 98224 379335
rect 98366 379264 98422 379273
rect 98366 379199 98422 379208
rect 99470 379264 99526 379273
rect 99470 379199 99526 379208
rect 98184 378888 98236 378894
rect 98184 378830 98236 378836
rect 96068 378684 96120 378690
rect 96068 378626 96120 378632
rect 97722 378584 97778 378593
rect 97722 378519 97778 378528
rect 95974 377904 96030 377913
rect 95974 377839 96030 377848
rect 97736 376514 97764 378519
rect 98380 377641 98408 379199
rect 98366 377632 98422 377641
rect 98366 377567 98422 377576
rect 97724 376508 97776 376514
rect 97724 376450 97776 376456
rect 94688 376168 94740 376174
rect 94688 376110 94740 376116
rect 99484 375902 99512 379199
rect 101048 379030 101076 379335
rect 102966 379264 103022 379273
rect 102966 379199 103022 379208
rect 101036 379024 101088 379030
rect 101036 378966 101088 378972
rect 100758 378448 100814 378457
rect 100758 378383 100814 378392
rect 99472 375896 99524 375902
rect 99472 375838 99524 375844
rect 100772 375698 100800 378383
rect 101954 378312 102010 378321
rect 101954 378247 102010 378256
rect 100760 375692 100812 375698
rect 100760 375634 100812 375640
rect 101968 375358 101996 378247
rect 101956 375352 102008 375358
rect 101956 375294 102008 375300
rect 102980 374746 103008 379199
rect 103532 378962 103560 379335
rect 103520 378956 103572 378962
rect 103520 378898 103572 378904
rect 104070 378448 104126 378457
rect 104070 378383 104126 378392
rect 104084 375766 104112 378383
rect 105372 377777 105400 379335
rect 108224 379098 108252 379335
rect 108212 379092 108264 379098
rect 108212 379034 108264 379040
rect 108868 378826 108896 379335
rect 111260 378894 111288 379335
rect 112364 379098 112392 379335
rect 112352 379092 112404 379098
rect 112352 379034 112404 379040
rect 111248 378888 111300 378894
rect 111248 378830 111300 378836
rect 108856 378820 108908 378826
rect 108856 378762 108908 378768
rect 113468 378350 113496 379335
rect 114480 378554 114508 379335
rect 115860 378690 115888 379335
rect 115848 378684 115900 378690
rect 115848 378626 115900 378632
rect 114468 378548 114520 378554
rect 114468 378490 114520 378496
rect 125966 378448 126022 378457
rect 125966 378383 126022 378392
rect 131026 378448 131082 378457
rect 131026 378383 131082 378392
rect 113456 378344 113508 378350
rect 113456 378286 113508 378292
rect 106462 378176 106518 378185
rect 106462 378111 106518 378120
rect 107566 378176 107622 378185
rect 107566 378111 107622 378120
rect 105358 377768 105414 377777
rect 105358 377703 105414 377712
rect 104072 375760 104124 375766
rect 104072 375702 104124 375708
rect 106476 375086 106504 378111
rect 107580 375222 107608 378111
rect 125980 376582 126008 378383
rect 125968 376576 126020 376582
rect 125968 376518 126020 376524
rect 131040 376310 131068 378383
rect 141068 377262 141096 379335
rect 143644 377534 143672 379335
rect 143632 377528 143684 377534
rect 143632 377470 143684 377476
rect 146036 377398 146064 379335
rect 146024 377392 146076 377398
rect 146024 377334 146076 377340
rect 141056 377256 141108 377262
rect 141056 377198 141108 377204
rect 151004 377126 151032 379335
rect 153580 377194 153608 379335
rect 195980 379160 196032 379166
rect 195980 379102 196032 379108
rect 195992 379030 196020 379102
rect 195980 379024 196032 379030
rect 195980 378966 196032 378972
rect 183466 378448 183522 378457
rect 183466 378383 183522 378392
rect 182270 378176 182326 378185
rect 182270 378111 182326 378120
rect 182822 378176 182878 378185
rect 182822 378111 182878 378120
rect 182284 377874 182312 378111
rect 182272 377868 182324 377874
rect 182272 377810 182324 377816
rect 153568 377188 153620 377194
rect 153568 377130 153620 377136
rect 150992 377120 151044 377126
rect 150992 377062 151044 377068
rect 131028 376304 131080 376310
rect 131028 376246 131080 376252
rect 107568 375216 107620 375222
rect 107568 375158 107620 375164
rect 106464 375080 106516 375086
rect 106464 375022 106516 375028
rect 102968 374740 103020 374746
rect 102968 374682 103020 374688
rect 179696 358896 179748 358902
rect 178590 358864 178646 358873
rect 178590 358799 178592 358808
rect 178644 358799 178646 358808
rect 179694 358864 179696 358873
rect 179748 358864 179750 358873
rect 179694 358799 179750 358808
rect 178592 358770 178644 358776
rect 182836 358086 182864 378111
rect 183480 377942 183508 378383
rect 183468 377936 183520 377942
rect 183468 377878 183520 377884
rect 183480 374678 183508 377878
rect 196636 377602 196664 488022
rect 196728 378146 196756 488036
rect 196820 488022 197110 488050
rect 197372 488022 197570 488050
rect 197648 488022 198030 488050
rect 198108 488022 198490 488050
rect 196716 378140 196768 378146
rect 196716 378082 196768 378088
rect 196820 377670 196848 488022
rect 197084 484424 197136 484430
rect 197084 484366 197136 484372
rect 196992 482588 197044 482594
rect 196992 482530 197044 482536
rect 196900 471640 196952 471646
rect 196900 471582 196952 471588
rect 196912 380322 196940 471582
rect 197004 465050 197032 482530
rect 196992 465044 197044 465050
rect 196992 464986 197044 464992
rect 196992 380928 197044 380934
rect 196992 380870 197044 380876
rect 196900 380316 196952 380322
rect 196900 380258 196952 380264
rect 196808 377664 196860 377670
rect 196808 377606 196860 377612
rect 196624 377596 196676 377602
rect 196624 377538 196676 377544
rect 183468 374672 183520 374678
rect 183468 374614 183520 374620
rect 190920 359508 190972 359514
rect 190920 359450 190972 359456
rect 190932 358873 190960 359450
rect 190918 358864 190974 358873
rect 190918 358799 190974 358808
rect 182824 358080 182876 358086
rect 182824 358022 182876 358028
rect 60740 357400 60792 357406
rect 60740 357342 60792 357348
rect 95974 273864 96030 273873
rect 95974 273799 96030 273808
rect 60832 273012 60884 273018
rect 60832 272954 60884 272960
rect 60740 272876 60792 272882
rect 60740 272818 60792 272824
rect 60752 252210 60780 272818
rect 60844 272785 60872 272954
rect 61108 272944 61160 272950
rect 61108 272886 61160 272892
rect 61476 272944 61528 272950
rect 61476 272886 61528 272892
rect 76010 272912 76066 272921
rect 60830 272776 60886 272785
rect 60830 272711 60886 272720
rect 61014 272776 61070 272785
rect 61014 272711 61070 272720
rect 60832 272196 60884 272202
rect 60832 272138 60884 272144
rect 60844 270609 60872 272138
rect 60830 270600 60886 270609
rect 60830 270535 60886 270544
rect 61028 270314 61056 272711
rect 60844 270286 61056 270314
rect 60844 252550 60872 270286
rect 61120 258074 61148 272886
rect 61488 272513 61516 272886
rect 61752 272876 61804 272882
rect 76010 272847 76066 272856
rect 90730 272912 90786 272921
rect 90730 272847 90786 272856
rect 93674 272912 93730 272921
rect 93674 272847 93730 272856
rect 95882 272912 95938 272921
rect 95882 272847 95938 272856
rect 61752 272818 61804 272824
rect 61764 272649 61792 272818
rect 61750 272640 61806 272649
rect 61750 272575 61806 272584
rect 61474 272504 61530 272513
rect 61474 272439 61530 272448
rect 76024 272406 76052 272847
rect 90744 272814 90772 272847
rect 90732 272808 90784 272814
rect 90732 272750 90784 272756
rect 93688 272746 93716 272847
rect 93676 272740 93728 272746
rect 93676 272682 93728 272688
rect 95896 272678 95924 272847
rect 95884 272672 95936 272678
rect 95884 272614 95936 272620
rect 76012 272400 76064 272406
rect 76012 272342 76064 272348
rect 95988 272338 96016 273799
rect 110970 273592 111026 273601
rect 110970 273527 110972 273536
rect 111024 273527 111026 273536
rect 133418 273592 133474 273601
rect 133418 273527 133474 273536
rect 135902 273592 135958 273601
rect 135902 273527 135958 273536
rect 138478 273592 138534 273601
rect 138478 273527 138534 273536
rect 140870 273592 140926 273601
rect 140870 273527 140926 273536
rect 110972 273498 111024 273504
rect 133432 273494 133460 273527
rect 133420 273488 133472 273494
rect 133420 273430 133472 273436
rect 135916 273426 135944 273527
rect 135904 273420 135956 273426
rect 135904 273362 135956 273368
rect 138492 273358 138520 273527
rect 138480 273352 138532 273358
rect 138480 273294 138532 273300
rect 140884 273290 140912 273527
rect 140872 273284 140924 273290
rect 140872 273226 140924 273232
rect 100758 273184 100814 273193
rect 100758 273119 100760 273128
rect 100812 273119 100814 273128
rect 100760 273090 100812 273096
rect 98458 272912 98514 272921
rect 98458 272847 98514 272856
rect 99378 272912 99434 272921
rect 99378 272847 99434 272856
rect 98472 272610 98500 272847
rect 98460 272604 98512 272610
rect 98460 272546 98512 272552
rect 99392 272474 99420 272847
rect 143538 272640 143594 272649
rect 143538 272575 143594 272584
rect 143552 272542 143580 272575
rect 143540 272536 143592 272542
rect 143540 272478 143592 272484
rect 99380 272468 99432 272474
rect 99380 272410 99432 272416
rect 96986 272368 97042 272377
rect 65340 272332 65392 272338
rect 65340 272274 65392 272280
rect 95976 272332 96028 272338
rect 96986 272303 97042 272312
rect 95976 272274 96028 272280
rect 65352 271425 65380 272274
rect 97000 272270 97028 272303
rect 67364 272264 67416 272270
rect 67364 272206 67416 272212
rect 96988 272264 97040 272270
rect 96988 272206 97040 272212
rect 113546 272232 113602 272241
rect 65338 271416 65394 271425
rect 65338 271351 65394 271360
rect 67376 271153 67404 272206
rect 94228 272196 94280 272202
rect 113546 272167 113602 272176
rect 94228 272138 94280 272144
rect 86960 272128 87012 272134
rect 86960 272070 87012 272076
rect 82820 272060 82872 272066
rect 82820 272002 82872 272008
rect 83464 272060 83516 272066
rect 83464 272002 83516 272008
rect 75920 271992 75972 271998
rect 75920 271934 75972 271940
rect 75932 271833 75960 271934
rect 82832 271833 82860 272002
rect 75918 271824 75974 271833
rect 75918 271759 75974 271768
rect 82818 271824 82874 271833
rect 82818 271759 82874 271768
rect 67362 271144 67418 271153
rect 67362 271079 67418 271088
rect 77298 271144 77354 271153
rect 77298 271079 77354 271088
rect 77312 271046 77340 271079
rect 77300 271040 77352 271046
rect 77300 270982 77352 270988
rect 78678 271008 78734 271017
rect 78678 270943 78680 270952
rect 78732 270943 78734 270952
rect 78680 270914 78732 270920
rect 81440 270428 81492 270434
rect 81440 270370 81492 270376
rect 63500 270360 63552 270366
rect 63500 270302 63552 270308
rect 63512 268598 63540 270302
rect 80060 270156 80112 270162
rect 80060 270098 80112 270104
rect 77852 269816 77904 269822
rect 77852 269758 77904 269764
rect 63500 268592 63552 268598
rect 63500 268534 63552 268540
rect 77864 268433 77892 269758
rect 80072 268530 80100 270098
rect 80060 268524 80112 268530
rect 80060 268466 80112 268472
rect 81452 268462 81480 270370
rect 81440 268456 81492 268462
rect 77850 268424 77906 268433
rect 81440 268398 81492 268404
rect 77850 268359 77906 268368
rect 60936 258046 61148 258074
rect 60832 252544 60884 252550
rect 60832 252486 60884 252492
rect 60936 252385 60964 258046
rect 60922 252376 60978 252385
rect 60922 252311 60978 252320
rect 60740 252204 60792 252210
rect 60740 252146 60792 252152
rect 75828 252068 75880 252074
rect 75828 252010 75880 252016
rect 75840 251190 75868 252010
rect 83476 252006 83504 272002
rect 86972 271833 87000 272070
rect 94240 271833 94268 272138
rect 98000 272060 98052 272066
rect 98000 272002 98052 272008
rect 98012 271833 98040 272002
rect 98644 271924 98696 271930
rect 98644 271866 98696 271872
rect 100760 271924 100812 271930
rect 100760 271866 100812 271872
rect 84198 271824 84254 271833
rect 84198 271759 84254 271768
rect 86958 271824 87014 271833
rect 86958 271759 87014 271768
rect 94226 271824 94282 271833
rect 94226 271759 94282 271768
rect 97998 271824 98054 271833
rect 97998 271759 98054 271768
rect 84212 270298 84240 271759
rect 84658 271688 84714 271697
rect 84658 271623 84714 271632
rect 84200 270292 84252 270298
rect 84200 270234 84252 270240
rect 84672 270094 84700 271623
rect 88338 271144 88394 271153
rect 88338 271079 88340 271088
rect 88392 271079 88394 271088
rect 88340 271050 88392 271056
rect 88338 271008 88394 271017
rect 88338 270943 88394 270952
rect 89718 271008 89774 271017
rect 89718 270943 89774 270952
rect 85578 270872 85634 270881
rect 85578 270807 85634 270816
rect 85592 270230 85620 270807
rect 85580 270224 85632 270230
rect 85580 270166 85632 270172
rect 84660 270088 84712 270094
rect 84660 270030 84712 270036
rect 88352 270026 88380 270943
rect 88340 270020 88392 270026
rect 88340 269962 88392 269968
rect 89732 269890 89760 270943
rect 92478 270872 92534 270881
rect 92478 270807 92534 270816
rect 91098 270600 91154 270609
rect 91098 270535 91154 270544
rect 91112 269958 91140 270535
rect 92492 270366 92520 270807
rect 92480 270360 92532 270366
rect 92480 270302 92532 270308
rect 91100 269952 91152 269958
rect 91100 269894 91152 269900
rect 89720 269884 89772 269890
rect 89720 269826 89772 269832
rect 98656 252074 98684 271866
rect 100772 271833 100800 271866
rect 100758 271824 100814 271833
rect 100758 271759 100814 271768
rect 103518 271688 103574 271697
rect 103518 271623 103574 271632
rect 100758 271416 100814 271425
rect 100758 271351 100814 271360
rect 100772 271182 100800 271351
rect 103532 271250 103560 271623
rect 104898 271416 104954 271425
rect 113560 271386 113588 272167
rect 114468 271924 114520 271930
rect 114468 271866 114520 271872
rect 127624 271924 127676 271930
rect 127624 271866 127676 271872
rect 114480 271833 114508 271866
rect 114466 271824 114522 271833
rect 114466 271759 114522 271768
rect 123206 271824 123262 271833
rect 123206 271759 123208 271768
rect 123260 271759 123262 271768
rect 123208 271730 123260 271736
rect 120078 271688 120134 271697
rect 120078 271623 120134 271632
rect 125598 271688 125654 271697
rect 125598 271623 125600 271632
rect 120092 271590 120120 271623
rect 125652 271623 125654 271632
rect 125600 271594 125652 271600
rect 120080 271584 120132 271590
rect 115938 271552 115994 271561
rect 115938 271487 115994 271496
rect 117318 271552 117374 271561
rect 127636 271561 127664 271866
rect 129740 271856 129792 271862
rect 128358 271824 128414 271833
rect 128358 271759 128414 271768
rect 129738 271824 129740 271833
rect 151360 271856 151412 271862
rect 129792 271824 129794 271833
rect 129738 271759 129794 271768
rect 151358 271824 151360 271833
rect 151412 271824 151414 271833
rect 151358 271759 151414 271768
rect 154486 271824 154542 271833
rect 154486 271759 154542 271768
rect 157246 271824 157302 271833
rect 157246 271759 157248 271768
rect 128372 271726 128400 271759
rect 154500 271726 154528 271759
rect 157300 271759 157302 271768
rect 196622 271824 196678 271833
rect 196622 271759 196678 271768
rect 157248 271730 157300 271736
rect 128360 271720 128412 271726
rect 128360 271662 128412 271668
rect 154488 271720 154540 271726
rect 154488 271662 154540 271668
rect 158626 271688 158682 271697
rect 158626 271623 158628 271632
rect 158680 271623 158682 271632
rect 161294 271688 161350 271697
rect 161294 271623 161350 271632
rect 164146 271688 164202 271697
rect 164146 271623 164202 271632
rect 158628 271594 158680 271600
rect 161308 271590 161336 271623
rect 161296 271584 161348 271590
rect 120080 271526 120132 271532
rect 127622 271552 127678 271561
rect 117318 271487 117320 271496
rect 115952 271454 115980 271487
rect 117372 271487 117374 271496
rect 161296 271526 161348 271532
rect 164160 271522 164188 271623
rect 196636 271561 196664 271759
rect 196622 271552 196678 271561
rect 127622 271487 127678 271496
rect 164148 271516 164200 271522
rect 117320 271458 117372 271464
rect 196622 271487 196678 271496
rect 164148 271458 164200 271464
rect 115940 271448 115992 271454
rect 115940 271390 115992 271396
rect 183466 271416 183522 271425
rect 104898 271351 104954 271360
rect 113548 271380 113600 271386
rect 104912 271318 104940 271351
rect 183466 271351 183522 271360
rect 113548 271322 113600 271328
rect 183480 271318 183508 271351
rect 104900 271312 104952 271318
rect 104900 271254 104952 271260
rect 183468 271312 183520 271318
rect 183468 271254 183520 271260
rect 103520 271244 103572 271250
rect 103520 271186 103572 271192
rect 100760 271176 100812 271182
rect 183468 271176 183520 271182
rect 100760 271118 100812 271124
rect 183466 271144 183468 271153
rect 183520 271144 183522 271153
rect 183466 271079 183522 271088
rect 106370 271008 106426 271017
rect 106370 270943 106426 270952
rect 107658 271008 107714 271017
rect 107658 270943 107714 270952
rect 111798 271008 111854 271017
rect 111798 270943 111854 270952
rect 104898 270872 104954 270881
rect 104898 270807 104954 270816
rect 106278 270872 106334 270881
rect 106278 270807 106334 270816
rect 98644 252068 98696 252074
rect 98644 252010 98696 252016
rect 83464 252000 83516 252006
rect 83464 251942 83516 251948
rect 104912 251870 104940 270807
rect 106292 251938 106320 270807
rect 106384 268394 106412 270943
rect 107672 270502 107700 270943
rect 110418 270736 110474 270745
rect 110418 270671 110474 270680
rect 107750 270600 107806 270609
rect 107750 270535 107806 270544
rect 109038 270600 109094 270609
rect 109038 270535 109094 270544
rect 107660 270496 107712 270502
rect 107660 270438 107712 270444
rect 107764 268938 107792 270535
rect 109052 270434 109080 270535
rect 109040 270428 109092 270434
rect 109040 270370 109092 270376
rect 107752 268932 107804 268938
rect 107752 268874 107804 268880
rect 110432 268870 110460 270671
rect 111812 270162 111840 270943
rect 113178 270600 113234 270609
rect 113178 270535 113234 270544
rect 115846 270600 115902 270609
rect 115846 270535 115902 270544
rect 117226 270600 117282 270609
rect 117226 270535 117282 270544
rect 144918 270600 144974 270609
rect 144918 270535 144974 270544
rect 147678 270600 147734 270609
rect 147678 270535 147734 270544
rect 111800 270156 111852 270162
rect 111800 270098 111852 270104
rect 113192 269822 113220 270535
rect 115860 270502 115888 270535
rect 115848 270496 115900 270502
rect 115848 270438 115900 270444
rect 117240 270434 117268 270535
rect 117228 270428 117280 270434
rect 117228 270370 117280 270376
rect 113180 269816 113232 269822
rect 113180 269758 113232 269764
rect 144932 269006 144960 270535
rect 144920 269000 144972 269006
rect 144920 268942 144972 268948
rect 110420 268864 110472 268870
rect 110420 268806 110472 268812
rect 106372 268388 106424 268394
rect 106372 268330 106424 268336
rect 147692 268326 147720 270535
rect 147680 268320 147732 268326
rect 147680 268262 147732 268268
rect 191748 253904 191800 253910
rect 191748 253846 191800 253852
rect 191760 253745 191788 253846
rect 191746 253736 191802 253745
rect 191746 253671 191802 253680
rect 180524 253292 180576 253298
rect 180524 253234 180576 253240
rect 179328 253224 179380 253230
rect 179326 253192 179328 253201
rect 180536 253201 180564 253234
rect 179380 253192 179382 253201
rect 179326 253127 179382 253136
rect 180522 253192 180578 253201
rect 180522 253127 180578 253136
rect 106280 251932 106332 251938
rect 106280 251874 106332 251880
rect 104900 251864 104952 251870
rect 104900 251806 104952 251812
rect 75828 251184 75880 251190
rect 75828 251126 75880 251132
rect 101036 167000 101088 167006
rect 101036 166942 101088 166948
rect 101048 166841 101076 166942
rect 103520 166932 103572 166938
rect 103520 166874 103572 166880
rect 103532 166841 103560 166874
rect 108304 166864 108356 166870
rect 101034 166832 101090 166841
rect 101034 166767 101090 166776
rect 103518 166832 103574 166841
rect 103518 166767 103574 166776
rect 108302 166832 108304 166841
rect 108356 166832 108358 166841
rect 108302 166767 108358 166776
rect 138478 166832 138534 166841
rect 138478 166767 138534 166776
rect 140870 166832 140926 166841
rect 140870 166767 140872 166776
rect 138492 166734 138520 166767
rect 140924 166767 140926 166776
rect 145930 166832 145986 166841
rect 145930 166767 145986 166776
rect 140872 166738 140924 166744
rect 138480 166728 138532 166734
rect 138480 166670 138532 166676
rect 145944 166666 145972 166767
rect 148506 166696 148562 166705
rect 60004 166660 60056 166666
rect 60004 166602 60056 166608
rect 145932 166660 145984 166666
rect 148506 166631 148562 166640
rect 163318 166696 163374 166705
rect 163318 166631 163374 166640
rect 165894 166696 165950 166705
rect 165894 166631 165950 166640
rect 145932 166602 145984 166608
rect 148520 166598 148548 166631
rect 148508 166592 148560 166598
rect 107658 166560 107714 166569
rect 59912 166524 59964 166530
rect 148508 166534 148560 166540
rect 150898 166560 150954 166569
rect 107658 166495 107714 166504
rect 150898 166495 150900 166504
rect 59912 166466 59964 166472
rect 96066 166288 96122 166297
rect 96066 166223 96122 166232
rect 98458 166288 98514 166297
rect 98458 166223 98460 166232
rect 96080 166190 96108 166223
rect 98512 166223 98514 166232
rect 98460 166194 98512 166200
rect 96068 166184 96120 166190
rect 96068 166126 96120 166132
rect 81438 165608 81494 165617
rect 81438 165543 81494 165552
rect 84290 165608 84346 165617
rect 84290 165543 84346 165552
rect 91190 165608 91246 165617
rect 91190 165543 91246 165552
rect 95238 165608 95294 165617
rect 95238 165543 95294 165552
rect 99378 165608 99434 165617
rect 99378 165543 99434 165552
rect 100850 165608 100906 165617
rect 100850 165543 100906 165552
rect 105174 165608 105230 165617
rect 105174 165543 105230 165552
rect 105726 165608 105782 165617
rect 105726 165543 105782 165552
rect 106370 165608 106426 165617
rect 106370 165543 106426 165552
rect 78678 164928 78734 164937
rect 78678 164863 78734 164872
rect 76010 164384 76066 164393
rect 76010 164319 76066 164328
rect 73804 164280 73856 164286
rect 73804 164222 73856 164228
rect 75918 164248 75974 164257
rect 60004 164212 60056 164218
rect 60004 164154 60056 164160
rect 60096 164212 60148 164218
rect 60096 164154 60148 164160
rect 60016 163810 60044 164154
rect 60004 163804 60056 163810
rect 60004 163746 60056 163752
rect 59912 148708 59964 148714
rect 59912 148650 59964 148656
rect 59728 146260 59780 146266
rect 59728 146202 59780 146208
rect 59636 145308 59688 145314
rect 59636 145250 59688 145256
rect 59648 142154 59676 145250
rect 59648 142126 59860 142154
rect 59358 140856 59414 140865
rect 59358 140791 59414 140800
rect 59832 59226 59860 142126
rect 59820 59220 59872 59226
rect 59820 59162 59872 59168
rect 59268 57384 59320 57390
rect 59268 57326 59320 57332
rect 59924 56302 59952 148650
rect 59912 56296 59964 56302
rect 59912 56238 59964 56244
rect 58808 55956 58860 55962
rect 58808 55898 58860 55904
rect 60016 54942 60044 163746
rect 60108 163402 60136 164154
rect 60096 163396 60148 163402
rect 60096 163338 60148 163344
rect 73816 146033 73844 164222
rect 75918 164183 75974 164192
rect 73802 146024 73858 146033
rect 73802 145959 73858 145968
rect 75932 145382 75960 164183
rect 76024 145450 76052 164319
rect 77298 164248 77354 164257
rect 77298 164183 77354 164192
rect 77312 145858 77340 164183
rect 77300 145852 77352 145858
rect 77300 145794 77352 145800
rect 78692 145790 78720 164863
rect 80058 164248 80114 164257
rect 80058 164183 80114 164192
rect 80072 148646 80100 164183
rect 80060 148640 80112 148646
rect 80060 148582 80112 148588
rect 81452 148578 81480 165543
rect 82818 164248 82874 164257
rect 82818 164183 82874 164192
rect 84198 164248 84254 164257
rect 84198 164183 84254 164192
rect 81440 148572 81492 148578
rect 81440 148514 81492 148520
rect 78680 145784 78732 145790
rect 78680 145726 78732 145732
rect 82832 145722 82860 164183
rect 82820 145716 82872 145722
rect 82820 145658 82872 145664
rect 84212 145654 84240 164183
rect 84200 145648 84252 145654
rect 84200 145590 84252 145596
rect 84304 145518 84332 165543
rect 90270 165064 90326 165073
rect 90270 164999 90326 165008
rect 88338 164928 88394 164937
rect 88338 164863 88394 164872
rect 88352 164762 88380 164863
rect 90284 164830 90312 164999
rect 90272 164824 90324 164830
rect 90272 164766 90324 164772
rect 88340 164756 88392 164762
rect 88340 164698 88392 164704
rect 87604 164280 87656 164286
rect 85578 164248 85634 164257
rect 85578 164183 85634 164192
rect 86958 164248 87014 164257
rect 87604 164222 87656 164228
rect 88430 164248 88486 164257
rect 86958 164183 87014 164192
rect 85592 145926 85620 164183
rect 86972 146130 87000 164183
rect 87616 148714 87644 164222
rect 88430 164183 88486 164192
rect 89902 164248 89958 164257
rect 89902 164183 89958 164192
rect 91098 164248 91154 164257
rect 91098 164183 91154 164192
rect 87604 148708 87656 148714
rect 87604 148650 87656 148656
rect 86960 146124 87012 146130
rect 86960 146066 87012 146072
rect 88444 145994 88472 164183
rect 89916 162246 89944 164183
rect 89904 162240 89956 162246
rect 89904 162182 89956 162188
rect 91112 146062 91140 164183
rect 91100 146056 91152 146062
rect 91100 145998 91152 146004
rect 88432 145988 88484 145994
rect 88432 145930 88484 145936
rect 85580 145920 85632 145926
rect 85580 145862 85632 145868
rect 91204 145586 91232 165543
rect 92478 164928 92534 164937
rect 92478 164863 92480 164872
rect 92532 164863 92534 164872
rect 92480 164834 92532 164840
rect 92570 164248 92626 164257
rect 92570 164183 92626 164192
rect 93858 164248 93914 164257
rect 93858 164183 93914 164192
rect 92584 145761 92612 164183
rect 92570 145752 92626 145761
rect 92570 145687 92626 145696
rect 91192 145580 91244 145586
rect 91192 145522 91244 145528
rect 84292 145512 84344 145518
rect 84292 145454 84344 145460
rect 76012 145444 76064 145450
rect 76012 145386 76064 145392
rect 75920 145376 75972 145382
rect 75920 145318 75972 145324
rect 93872 145314 93900 164183
rect 95252 163470 95280 165543
rect 96618 164248 96674 164257
rect 96618 164183 96674 164192
rect 97998 164248 98054 164257
rect 97998 164183 98054 164192
rect 96632 163946 96660 164183
rect 96620 163940 96672 163946
rect 96620 163882 96672 163888
rect 98012 163878 98040 164183
rect 98000 163872 98052 163878
rect 98000 163814 98052 163820
rect 95240 163464 95292 163470
rect 95240 163406 95292 163412
rect 99392 146266 99420 165543
rect 100758 164248 100814 164257
rect 100758 164183 100814 164192
rect 99380 146260 99432 146266
rect 99380 146202 99432 146208
rect 100772 146033 100800 164183
rect 100864 164014 100892 165543
rect 102138 164248 102194 164257
rect 102138 164183 102194 164192
rect 103518 164248 103574 164257
rect 103518 164183 103574 164192
rect 100852 164008 100904 164014
rect 100852 163950 100904 163956
rect 102152 146169 102180 164183
rect 103532 146305 103560 164183
rect 105188 164082 105216 165543
rect 105740 164966 105768 165543
rect 105728 164960 105780 164966
rect 105728 164902 105780 164908
rect 105176 164076 105228 164082
rect 105176 164018 105228 164024
rect 106384 163810 106412 165543
rect 106372 163804 106424 163810
rect 106372 163746 106424 163752
rect 103518 146296 103574 146305
rect 103518 146231 103574 146240
rect 102138 146160 102194 146169
rect 102138 146095 102194 146104
rect 100758 146024 100814 146033
rect 100758 145959 100814 145968
rect 107672 145625 107700 166495
rect 150952 166495 150954 166504
rect 153290 166560 153346 166569
rect 153290 166495 153346 166504
rect 150900 166466 150952 166472
rect 153304 166462 153332 166495
rect 153292 166456 153344 166462
rect 153292 166398 153344 166404
rect 163332 166394 163360 166631
rect 163320 166388 163372 166394
rect 163320 166330 163372 166336
rect 165908 166326 165936 166631
rect 183282 166560 183338 166569
rect 183282 166495 183338 166504
rect 165896 166320 165948 166326
rect 165896 166262 165948 166268
rect 108302 165608 108358 165617
rect 108302 165543 108358 165552
rect 109682 165608 109738 165617
rect 109682 165543 109738 165552
rect 110970 165608 111026 165617
rect 110970 165543 111026 165552
rect 111890 165608 111946 165617
rect 111890 165543 111946 165552
rect 113546 165608 113602 165617
rect 113546 165543 113602 165552
rect 115938 165608 115994 165617
rect 115938 165543 115994 165552
rect 117870 165608 117926 165617
rect 117870 165543 117926 165552
rect 118330 165608 118386 165617
rect 118330 165543 118386 165552
rect 119066 165608 119122 165617
rect 119066 165543 119122 165552
rect 120906 165608 120962 165617
rect 120906 165543 120962 165552
rect 123482 165608 123538 165617
rect 123482 165543 123538 165552
rect 125874 165608 125930 165617
rect 125874 165543 125930 165552
rect 128358 165608 128414 165617
rect 128358 165543 128414 165552
rect 129738 165608 129794 165617
rect 129738 165543 129794 165552
rect 132498 165608 132554 165617
rect 132498 165543 132500 165552
rect 108316 164286 108344 165543
rect 108304 164280 108356 164286
rect 108304 164222 108356 164228
rect 109696 163742 109724 165543
rect 110984 164150 111012 165543
rect 111154 164656 111210 164665
rect 111154 164591 111210 164600
rect 110972 164144 111024 164150
rect 110972 164086 111024 164092
rect 109684 163736 109736 163742
rect 109684 163678 109736 163684
rect 111168 162178 111196 164591
rect 111904 163606 111932 165543
rect 113178 165064 113234 165073
rect 113560 165034 113588 165543
rect 115952 165170 115980 165543
rect 115940 165164 115992 165170
rect 115940 165106 115992 165112
rect 113178 164999 113234 165008
rect 113548 165028 113600 165034
rect 111892 163600 111944 163606
rect 111892 163542 111944 163548
rect 113192 163538 113220 164999
rect 113548 164970 113600 164976
rect 117320 165028 117372 165034
rect 117320 164970 117372 164976
rect 115940 164960 115992 164966
rect 114466 164928 114522 164937
rect 114522 164898 114600 164914
rect 115940 164902 115992 164908
rect 114522 164892 114612 164898
rect 114522 164886 114560 164892
rect 114466 164863 114522 164872
rect 114560 164834 114612 164840
rect 113180 163532 113232 163538
rect 113180 163474 113232 163480
rect 111156 162172 111208 162178
rect 111156 162114 111208 162120
rect 114572 148510 114600 164834
rect 115952 164529 115980 164902
rect 117332 164529 117360 164970
rect 115938 164520 115994 164529
rect 115938 164455 115994 164464
rect 117318 164520 117374 164529
rect 117318 164455 117374 164464
rect 114560 148504 114612 148510
rect 114560 148446 114612 148452
rect 115952 148374 115980 164455
rect 117332 148442 117360 164455
rect 117884 164218 117912 165543
rect 118344 165102 118372 165543
rect 118332 165096 118384 165102
rect 118332 165038 118384 165044
rect 117872 164212 117924 164218
rect 117872 164154 117924 164160
rect 119080 163674 119108 165543
rect 120920 165238 120948 165543
rect 123496 165374 123524 165543
rect 123484 165368 123536 165374
rect 123484 165310 123536 165316
rect 125888 165306 125916 165543
rect 128372 165510 128400 165543
rect 128360 165504 128412 165510
rect 128360 165446 128412 165452
rect 129752 165442 129780 165543
rect 132552 165543 132554 165552
rect 132500 165514 132552 165520
rect 129740 165436 129792 165442
rect 129740 165378 129792 165384
rect 125876 165300 125928 165306
rect 125876 165242 125928 165248
rect 183296 165238 183324 166495
rect 183374 165608 183430 165617
rect 183374 165543 183430 165552
rect 120908 165232 120960 165238
rect 120908 165174 120960 165180
rect 183284 165232 183336 165238
rect 183284 165174 183336 165180
rect 183388 165102 183416 165543
rect 183376 165096 183428 165102
rect 183376 165038 183428 165044
rect 196636 164898 196664 271487
rect 197004 270502 197032 380870
rect 197096 377466 197124 484366
rect 197268 468308 197320 468314
rect 197268 468250 197320 468256
rect 197176 380996 197228 381002
rect 197176 380938 197228 380944
rect 197084 377460 197136 377466
rect 197084 377402 197136 377408
rect 196992 270496 197044 270502
rect 196992 270438 197044 270444
rect 197004 267734 197032 270438
rect 197188 270434 197216 380938
rect 197280 379030 197308 468250
rect 197268 379024 197320 379030
rect 197268 378966 197320 378972
rect 197372 377738 197400 488022
rect 197452 484968 197504 484974
rect 197450 484936 197452 484945
rect 197504 484936 197506 484945
rect 197450 484871 197506 484880
rect 197648 484106 197676 488022
rect 197464 484078 197676 484106
rect 197464 377806 197492 484078
rect 198108 483970 198136 488022
rect 198740 484152 198792 484158
rect 198740 484094 198792 484100
rect 197556 483942 198136 483970
rect 197556 377874 197584 483942
rect 198096 482520 198148 482526
rect 198096 482462 198148 482468
rect 197636 471368 197688 471374
rect 197636 471310 197688 471316
rect 197544 377868 197596 377874
rect 197544 377810 197596 377816
rect 197452 377800 197504 377806
rect 197452 377742 197504 377748
rect 197360 377732 197412 377738
rect 197360 377674 197412 377680
rect 197360 374672 197412 374678
rect 197360 374614 197412 374620
rect 197372 271318 197400 374614
rect 197452 359576 197504 359582
rect 197452 359518 197504 359524
rect 197464 358834 197492 359518
rect 197452 358828 197504 358834
rect 197452 358770 197504 358776
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 197176 270428 197228 270434
rect 197176 270370 197228 270376
rect 196728 267706 197032 267734
rect 196728 164966 196756 267706
rect 197188 258074 197216 270370
rect 196820 258046 197216 258074
rect 196820 165034 196848 258046
rect 197372 165238 197400 271254
rect 197464 267734 197492 358770
rect 197648 271590 197676 471310
rect 197728 468716 197780 468722
rect 197728 468658 197780 468664
rect 197636 271584 197688 271590
rect 197636 271526 197688 271532
rect 197740 271522 197768 468658
rect 197820 465996 197872 466002
rect 197820 465938 197872 465944
rect 197832 379982 197860 465938
rect 198004 464704 198056 464710
rect 198004 464646 198056 464652
rect 197912 464432 197964 464438
rect 197912 464374 197964 464380
rect 197924 380186 197952 464374
rect 198016 380934 198044 464646
rect 198108 414730 198136 482462
rect 198096 414724 198148 414730
rect 198096 414666 198148 414672
rect 198096 397588 198148 397594
rect 198096 397530 198148 397536
rect 198004 380928 198056 380934
rect 198004 380870 198056 380876
rect 198108 380882 198136 397530
rect 198188 396840 198240 396846
rect 198188 396782 198240 396788
rect 198200 381002 198228 396782
rect 198646 381032 198702 381041
rect 198188 380996 198240 381002
rect 198646 380967 198702 380976
rect 198188 380938 198240 380944
rect 198280 380928 198332 380934
rect 198108 380854 198228 380882
rect 198280 380870 198332 380876
rect 197912 380180 197964 380186
rect 197912 380122 197964 380128
rect 197820 379976 197872 379982
rect 197820 379918 197872 379924
rect 198200 377126 198228 380854
rect 198188 377120 198240 377126
rect 198188 377062 198240 377068
rect 198292 373994 198320 380870
rect 198016 373966 198320 373994
rect 198016 271862 198044 373966
rect 198096 358760 198148 358766
rect 198096 358702 198148 358708
rect 198004 271856 198056 271862
rect 198004 271798 198056 271804
rect 197728 271516 197780 271522
rect 197728 271458 197780 271464
rect 197464 267706 197584 267734
rect 197556 253230 197584 267706
rect 198108 253298 198136 358702
rect 197636 253292 197688 253298
rect 197636 253234 197688 253240
rect 198096 253292 198148 253298
rect 198096 253234 198148 253240
rect 197544 253224 197596 253230
rect 197544 253166 197596 253172
rect 197452 167000 197504 167006
rect 197452 166942 197504 166948
rect 197360 165232 197412 165238
rect 197360 165174 197412 165180
rect 196808 165028 196860 165034
rect 196808 164970 196860 164976
rect 196716 164960 196768 164966
rect 196716 164902 196768 164908
rect 196624 164892 196676 164898
rect 196624 164834 196676 164840
rect 119068 163668 119120 163674
rect 119068 163610 119120 163616
rect 117320 148436 117372 148442
rect 117320 148378 117372 148384
rect 115940 148368 115992 148374
rect 115940 148310 115992 148316
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 107658 145616 107714 145625
rect 107658 145551 107714 145560
rect 93860 145308 93912 145314
rect 93860 145250 93912 145256
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 191288 145580 191340 145586
rect 191288 145522 191340 145528
rect 191300 144945 191328 145522
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 191286 144936 191342 144945
rect 191286 144871 191342 144880
rect 77114 59800 77170 59809
rect 77114 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 94502 59800 94558 59809
rect 94502 59735 94558 59744
rect 99470 59800 99526 59809
rect 99470 59735 99526 59744
rect 102782 59800 102838 59809
rect 102782 59735 102838 59744
rect 105910 59800 105966 59809
rect 105910 59735 105966 59744
rect 77128 59702 77156 59735
rect 77116 59696 77168 59702
rect 77116 59638 77168 59644
rect 83108 59566 83136 59735
rect 83096 59560 83148 59566
rect 83096 59502 83148 59508
rect 89994 59528 90050 59537
rect 89994 59463 90050 59472
rect 84200 59356 84252 59362
rect 84200 59298 84252 59304
rect 84212 58041 84240 59298
rect 90008 59294 90036 59463
rect 89996 59288 90048 59294
rect 89996 59230 90048 59236
rect 94516 59226 94544 59735
rect 95882 59528 95938 59537
rect 95882 59463 95938 59472
rect 96986 59528 97042 59537
rect 99484 59498 99512 59735
rect 100760 59628 100812 59634
rect 100760 59570 100812 59576
rect 100772 59537 100800 59570
rect 100758 59528 100814 59537
rect 96986 59463 97042 59472
rect 99472 59492 99524 59498
rect 94504 59220 94556 59226
rect 94504 59162 94556 59168
rect 95896 59158 95924 59463
rect 95884 59152 95936 59158
rect 95884 59094 95936 59100
rect 97000 59090 97028 59463
rect 100758 59463 100814 59472
rect 101770 59528 101826 59537
rect 101770 59463 101826 59472
rect 99472 59434 99524 59440
rect 96988 59084 97040 59090
rect 96988 59026 97040 59032
rect 101784 58886 101812 59463
rect 102796 59022 102824 59735
rect 105924 59430 105952 59735
rect 107566 59664 107622 59673
rect 107566 59599 107622 59608
rect 105912 59424 105964 59430
rect 105912 59366 105964 59372
rect 102784 59016 102836 59022
rect 102784 58958 102836 58964
rect 107580 58954 107608 59599
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 138386 58984 138442 58993
rect 107568 58948 107620 58954
rect 138386 58919 138442 58928
rect 107568 58890 107620 58896
rect 101772 58880 101824 58886
rect 101772 58822 101824 58828
rect 138400 58818 138428 58919
rect 138388 58812 138440 58818
rect 138388 58754 138440 58760
rect 148520 58750 148548 59191
rect 148508 58744 148560 58750
rect 148508 58686 148560 58692
rect 150912 58682 150940 59191
rect 150900 58676 150952 58682
rect 150900 58618 150952 58624
rect 84198 58032 84254 58041
rect 84198 57967 84254 57976
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 78678 57896 78734 57905
rect 78678 57831 78734 57840
rect 80426 57896 80482 57905
rect 80426 57831 80482 57840
rect 81438 57896 81494 57905
rect 81438 57831 81494 57840
rect 85394 57896 85450 57905
rect 85394 57831 85450 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88338 57896 88394 57905
rect 88338 57831 88394 57840
rect 88706 57896 88762 57905
rect 88706 57831 88762 57840
rect 89718 57896 89774 57905
rect 89718 57831 89774 57840
rect 91098 57896 91154 57905
rect 91098 57831 91154 57840
rect 91466 57896 91522 57905
rect 91466 57831 91522 57840
rect 93306 57896 93362 57905
rect 93306 57831 93362 57840
rect 93674 57896 93730 57905
rect 93674 57831 93730 57840
rect 98090 57896 98146 57905
rect 98090 57831 98146 57840
rect 103794 57896 103850 57905
rect 103794 57831 103850 57840
rect 108578 57896 108634 57905
rect 108578 57831 108634 57840
rect 109498 57896 109554 57905
rect 109498 57831 109554 57840
rect 112074 57896 112130 57905
rect 112074 57831 112130 57840
rect 113178 57896 113234 57905
rect 113178 57831 113234 57840
rect 114098 57896 114154 57905
rect 114098 57831 114154 57840
rect 115938 57896 115994 57905
rect 115938 57831 115994 57840
rect 117870 57896 117926 57905
rect 117870 57831 117926 57840
rect 119066 57896 119122 57905
rect 119066 57831 119122 57840
rect 123482 57896 123538 57905
rect 123482 57831 123538 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 76024 57254 76052 57831
rect 78232 57322 78260 57831
rect 78220 57316 78272 57322
rect 78220 57258 78272 57264
rect 76012 57248 76064 57254
rect 76012 57190 76064 57196
rect 77852 56636 77904 56642
rect 77852 56578 77904 56584
rect 60004 54936 60056 54942
rect 60004 54878 60056 54884
rect 77864 54777 77892 56578
rect 77850 54768 77906 54777
rect 58624 54732 58676 54738
rect 77850 54703 77906 54712
rect 58624 54674 58676 54680
rect 78692 54602 78720 57831
rect 80440 56030 80468 57831
rect 80428 56024 80480 56030
rect 80428 55966 80480 55972
rect 81452 54670 81480 57831
rect 85408 55962 85436 57831
rect 86512 56098 86540 57831
rect 86500 56092 86552 56098
rect 86500 56034 86552 56040
rect 85396 55956 85448 55962
rect 85396 55898 85448 55904
rect 86972 54806 87000 57831
rect 88352 57458 88380 57831
rect 88340 57452 88392 57458
rect 88340 57394 88392 57400
rect 88720 56166 88748 57831
rect 88708 56160 88760 56166
rect 88708 56102 88760 56108
rect 89732 55010 89760 57831
rect 89720 55004 89772 55010
rect 89720 54946 89772 54952
rect 91112 54874 91140 57831
rect 91100 54868 91152 54874
rect 91100 54810 91152 54816
rect 86960 54800 87012 54806
rect 86960 54742 87012 54748
rect 91480 54738 91508 57831
rect 93320 56234 93348 57831
rect 93688 57390 93716 57831
rect 98104 57526 98132 57831
rect 103808 57594 103836 57831
rect 103796 57588 103848 57594
rect 103796 57530 103848 57536
rect 98092 57520 98144 57526
rect 98092 57462 98144 57468
rect 106278 57488 106334 57497
rect 106278 57423 106334 57432
rect 93676 57384 93728 57390
rect 93676 57326 93728 57332
rect 93308 56228 93360 56234
rect 93308 56170 93360 56176
rect 106292 54942 106320 57423
rect 108592 56302 108620 57831
rect 109512 56370 109540 57831
rect 110418 57488 110474 57497
rect 110418 57423 110474 57432
rect 109500 56364 109552 56370
rect 109500 56306 109552 56312
rect 108580 56296 108632 56302
rect 108580 56238 108632 56244
rect 110432 55078 110460 57423
rect 112088 56506 112116 57831
rect 113192 57662 113220 57831
rect 113180 57656 113232 57662
rect 113180 57598 113232 57604
rect 112076 56500 112128 56506
rect 112076 56442 112128 56448
rect 114112 56438 114140 57831
rect 114558 57488 114614 57497
rect 114558 57423 114614 57432
rect 114100 56432 114152 56438
rect 114100 56374 114152 56380
rect 114572 55214 114600 57423
rect 115952 56574 115980 57831
rect 116122 57488 116178 57497
rect 116122 57423 116178 57432
rect 115940 56568 115992 56574
rect 115940 56510 115992 56516
rect 114560 55208 114612 55214
rect 114560 55150 114612 55156
rect 116136 55146 116164 57423
rect 117884 56642 117912 57831
rect 117872 56636 117924 56642
rect 117872 56578 117924 56584
rect 119080 56137 119108 57831
rect 123496 57798 123524 57831
rect 123484 57792 123536 57798
rect 123484 57734 123536 57740
rect 130856 57730 130884 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 183466 57896 183522 57905
rect 183466 57831 183468 57840
rect 145564 57802 145616 57808
rect 130844 57724 130896 57730
rect 130844 57666 130896 57672
rect 153304 56409 153332 57831
rect 183520 57831 183522 57840
rect 183468 57802 183520 57808
rect 197372 57798 197400 165174
rect 197464 165102 197492 166942
rect 197452 165096 197504 165102
rect 197452 165038 197504 165044
rect 197464 57866 197492 165038
rect 197556 146266 197584 253166
rect 197544 146260 197596 146266
rect 197544 146202 197596 146208
rect 197648 146198 197676 253234
rect 197636 146192 197688 146198
rect 197636 146134 197688 146140
rect 198660 58750 198688 380967
rect 198752 378049 198780 484094
rect 198738 378040 198794 378049
rect 198738 377975 198794 377984
rect 198844 377942 198872 488036
rect 198936 488022 199318 488050
rect 199794 488022 199976 488050
rect 200254 488022 200436 488050
rect 200714 488022 200988 488050
rect 198936 484158 198964 488022
rect 199016 486532 199068 486538
rect 199016 486474 199068 486480
rect 198924 484152 198976 484158
rect 198924 484094 198976 484100
rect 198924 465724 198976 465730
rect 198924 465666 198976 465672
rect 198936 465118 198964 465666
rect 198924 465112 198976 465118
rect 198924 465054 198976 465060
rect 198936 460193 198964 465054
rect 198922 460184 198978 460193
rect 198922 460119 198978 460128
rect 198832 377936 198884 377942
rect 198832 377878 198884 377884
rect 198936 354674 198964 460119
rect 199028 397594 199056 486474
rect 199948 485110 199976 488022
rect 200408 485314 200436 488022
rect 200304 485308 200356 485314
rect 200304 485250 200356 485256
rect 200396 485308 200448 485314
rect 200396 485250 200448 485256
rect 199936 485104 199988 485110
rect 199936 485046 199988 485052
rect 200316 484537 200344 485250
rect 200488 485240 200540 485246
rect 200488 485182 200540 485188
rect 200500 484809 200528 485182
rect 200486 484800 200542 484809
rect 200486 484735 200542 484744
rect 200302 484528 200358 484537
rect 200302 484463 200358 484472
rect 200212 484152 200264 484158
rect 200212 484094 200264 484100
rect 199292 478168 199344 478174
rect 199292 478110 199344 478116
rect 199108 468648 199160 468654
rect 199108 468590 199160 468596
rect 199016 397588 199068 397594
rect 199016 397530 199068 397536
rect 199014 397488 199070 397497
rect 199014 397423 199070 397432
rect 199028 379522 199056 397423
rect 199120 380934 199148 468590
rect 199200 464364 199252 464370
rect 199200 464306 199252 464312
rect 199108 380928 199160 380934
rect 199108 380870 199160 380876
rect 199212 380254 199240 464306
rect 199304 396001 199332 478110
rect 199384 476808 199436 476814
rect 199384 476750 199436 476756
rect 199290 395992 199346 396001
rect 199290 395927 199346 395936
rect 199396 394641 199424 476750
rect 199476 469872 199528 469878
rect 199476 469814 199528 469820
rect 199488 400353 199516 469814
rect 199568 464636 199620 464642
rect 199568 464578 199620 464584
rect 199474 400344 199530 400353
rect 199474 400279 199530 400288
rect 199580 396846 199608 464578
rect 199842 400344 199898 400353
rect 199842 400279 199898 400288
rect 199568 396840 199620 396846
rect 199568 396782 199620 396788
rect 199658 396808 199714 396817
rect 199658 396743 199714 396752
rect 199382 394632 199438 394641
rect 199382 394567 199438 394576
rect 199200 380248 199252 380254
rect 199200 380190 199252 380196
rect 199028 379494 199516 379522
rect 199014 379400 199070 379409
rect 199014 379335 199070 379344
rect 199028 378894 199056 379335
rect 199016 378888 199068 378894
rect 199016 378830 199068 378836
rect 199028 378486 199056 378830
rect 199016 378480 199068 378486
rect 199016 378422 199068 378428
rect 199488 377505 199516 379494
rect 199672 378010 199700 396743
rect 199750 394632 199806 394641
rect 199750 394567 199806 394576
rect 199660 378004 199712 378010
rect 199660 377946 199712 377952
rect 199474 377496 199530 377505
rect 199474 377431 199530 377440
rect 199384 371884 199436 371890
rect 199384 371826 199436 371832
rect 198844 354646 198964 354674
rect 198844 353161 198872 354646
rect 198830 353152 198886 353161
rect 198830 353087 198886 353096
rect 198738 291680 198794 291689
rect 198738 291615 198794 291624
rect 198752 184929 198780 291615
rect 198844 246265 198872 353087
rect 199396 296714 199424 371826
rect 199488 370530 199516 377431
rect 199672 373994 199700 377946
rect 199580 373966 199700 373994
rect 199476 370524 199528 370530
rect 199476 370466 199528 370472
rect 198936 296686 199424 296714
rect 198936 288833 198964 296686
rect 199198 292768 199254 292777
rect 199198 292703 199254 292712
rect 199106 291000 199162 291009
rect 199106 290935 199162 290944
rect 198922 288824 198978 288833
rect 198922 288759 198978 288768
rect 198830 246256 198886 246265
rect 198830 246191 198886 246200
rect 198738 184920 198794 184929
rect 198738 184855 198794 184864
rect 198738 182064 198794 182073
rect 198738 181999 198794 182008
rect 198752 74905 198780 181999
rect 198844 139233 198872 246191
rect 198936 182073 198964 288759
rect 199014 288416 199070 288425
rect 199014 288351 199070 288360
rect 199028 287609 199056 288351
rect 199014 287600 199070 287609
rect 199014 287535 199070 287544
rect 198922 182064 198978 182073
rect 198922 181999 198978 182008
rect 199028 180713 199056 287535
rect 199120 183433 199148 290935
rect 199212 209774 199240 292703
rect 199488 291689 199516 370466
rect 199580 366382 199608 373966
rect 199660 369164 199712 369170
rect 199660 369106 199712 369112
rect 199568 366376 199620 366382
rect 199568 366318 199620 366324
rect 199474 291680 199530 291689
rect 199474 291615 199530 291624
rect 199580 291009 199608 366318
rect 199672 292777 199700 369106
rect 199764 362234 199792 394567
rect 199856 369170 199884 400279
rect 199934 395992 199990 396001
rect 199934 395927 199990 395936
rect 199948 371890 199976 395927
rect 200224 380254 200252 484094
rect 200396 482452 200448 482458
rect 200396 482394 200448 482400
rect 200304 468580 200356 468586
rect 200304 468522 200356 468528
rect 200212 380248 200264 380254
rect 200212 380190 200264 380196
rect 199936 371884 199988 371890
rect 199936 371826 199988 371832
rect 199844 369164 199896 369170
rect 199844 369106 199896 369112
rect 199752 362228 199804 362234
rect 199752 362170 199804 362176
rect 199658 292768 199714 292777
rect 199658 292703 199714 292712
rect 199566 291000 199622 291009
rect 199566 290935 199622 290944
rect 199764 288425 199792 362170
rect 199750 288416 199806 288425
rect 199750 288351 199806 288360
rect 200316 271726 200344 468522
rect 200408 380526 200436 482394
rect 200960 480254 200988 488022
rect 201052 484158 201080 488036
rect 201528 487830 201556 488036
rect 201696 488022 201986 488050
rect 202064 488022 202446 488050
rect 202922 488022 203012 488050
rect 203290 488022 203656 488050
rect 203750 488022 203840 488050
rect 201516 487824 201568 487830
rect 201516 487766 201568 487772
rect 201500 485036 201552 485042
rect 201500 484978 201552 484984
rect 201512 484945 201540 484978
rect 201498 484936 201554 484945
rect 201498 484871 201554 484880
rect 201040 484152 201092 484158
rect 201040 484094 201092 484100
rect 201500 484152 201552 484158
rect 201500 484094 201552 484100
rect 200960 480226 201080 480254
rect 200764 479596 200816 479602
rect 200764 479538 200816 479544
rect 200488 471572 200540 471578
rect 200488 471514 200540 471520
rect 200396 380520 200448 380526
rect 200396 380462 200448 380468
rect 200500 377194 200528 471514
rect 200580 465928 200632 465934
rect 200580 465870 200632 465876
rect 200592 380050 200620 465870
rect 200672 465044 200724 465050
rect 200672 464986 200724 464992
rect 200684 380458 200712 464986
rect 200672 380452 200724 380458
rect 200672 380394 200724 380400
rect 200580 380044 200632 380050
rect 200580 379986 200632 379992
rect 200488 377188 200540 377194
rect 200488 377130 200540 377136
rect 200776 271726 200804 479538
rect 200856 471844 200908 471850
rect 200856 471786 200908 471792
rect 200868 273562 200896 471786
rect 200948 465588 201000 465594
rect 200948 465530 201000 465536
rect 200960 284306 200988 465530
rect 201052 380322 201080 480226
rect 201040 380316 201092 380322
rect 201040 380258 201092 380264
rect 201314 379536 201370 379545
rect 201314 379471 201370 379480
rect 200948 284300 201000 284306
rect 200948 284242 201000 284248
rect 200856 273556 200908 273562
rect 200856 273498 200908 273504
rect 200304 271720 200356 271726
rect 200304 271662 200356 271668
rect 200764 271720 200816 271726
rect 200764 271662 200816 271668
rect 199212 209746 199424 209774
rect 199396 186425 199424 209746
rect 199382 186416 199438 186425
rect 199382 186351 199438 186360
rect 199290 184920 199346 184929
rect 199290 184855 199346 184864
rect 199106 183424 199162 183433
rect 199106 183359 199162 183368
rect 199014 180704 199070 180713
rect 199014 180639 199070 180648
rect 199028 179489 199056 180639
rect 199014 179480 199070 179489
rect 199014 179415 199070 179424
rect 198830 139224 198886 139233
rect 198830 139159 198886 139168
rect 199120 76401 199148 183359
rect 199198 179480 199254 179489
rect 199198 179415 199254 179424
rect 199106 76392 199162 76401
rect 199106 76327 199162 76336
rect 198738 74896 198794 74905
rect 198738 74831 198794 74840
rect 199212 73681 199240 179415
rect 199304 77761 199332 184855
rect 199396 79393 199424 186351
rect 199382 79384 199438 79393
rect 199382 79319 199438 79328
rect 199290 77752 199346 77761
rect 199290 77687 199346 77696
rect 199198 73672 199254 73681
rect 199198 73607 199254 73616
rect 201328 59022 201356 379471
rect 201512 376650 201540 484094
rect 201696 480254 201724 488022
rect 201776 487824 201828 487830
rect 201776 487766 201828 487772
rect 201604 480226 201724 480254
rect 201604 378010 201632 480226
rect 201684 471300 201736 471306
rect 201684 471242 201736 471248
rect 201592 378004 201644 378010
rect 201592 377946 201644 377952
rect 201500 376644 201552 376650
rect 201500 376586 201552 376592
rect 201500 359508 201552 359514
rect 201500 359450 201552 359456
rect 201512 282878 201540 359450
rect 201592 358080 201644 358086
rect 201592 358022 201644 358028
rect 201500 282872 201552 282878
rect 201500 282814 201552 282820
rect 201512 282418 201540 282814
rect 201420 282390 201540 282418
rect 201420 253910 201448 282390
rect 201604 271182 201632 358022
rect 201696 271658 201724 471242
rect 201788 380186 201816 487766
rect 202064 484158 202092 488022
rect 202052 484152 202104 484158
rect 202052 484094 202104 484100
rect 202880 484152 202932 484158
rect 202880 484094 202932 484100
rect 202236 474224 202288 474230
rect 202236 474166 202288 474172
rect 201868 470688 201920 470694
rect 201868 470630 201920 470636
rect 201776 380180 201828 380186
rect 201776 380122 201828 380128
rect 201880 377262 201908 470630
rect 202144 467492 202196 467498
rect 202144 467434 202196 467440
rect 201868 377256 201920 377262
rect 201868 377198 201920 377204
rect 202156 376106 202184 467434
rect 202144 376100 202196 376106
rect 202144 376042 202196 376048
rect 201684 271652 201736 271658
rect 201684 271594 201736 271600
rect 201592 271176 201644 271182
rect 201592 271118 201644 271124
rect 201604 258074 201632 271118
rect 201512 258046 201632 258074
rect 201408 253904 201460 253910
rect 201408 253846 201460 253852
rect 201512 167006 201540 258046
rect 202144 176180 202196 176186
rect 202144 176122 202196 176128
rect 201500 167000 201552 167006
rect 201500 166942 201552 166948
rect 202156 145586 202184 176122
rect 202144 145580 202196 145586
rect 202144 145522 202196 145528
rect 202248 70378 202276 474166
rect 202420 472796 202472 472802
rect 202420 472738 202472 472744
rect 202326 469024 202382 469033
rect 202326 468959 202382 468968
rect 202340 166326 202368 468959
rect 202432 271182 202460 472738
rect 202512 468376 202564 468382
rect 202512 468318 202564 468324
rect 202524 272746 202552 468318
rect 202892 380769 202920 484094
rect 202878 380760 202934 380769
rect 202878 380695 202934 380704
rect 202892 380526 202920 380695
rect 202880 380520 202932 380526
rect 202880 380462 202932 380468
rect 202984 380458 203012 488022
rect 203628 485081 203656 488022
rect 203614 485072 203670 485081
rect 203614 485007 203670 485016
rect 203812 484090 203840 488022
rect 203904 488022 204194 488050
rect 204272 488022 204654 488050
rect 204732 488022 205022 488050
rect 205192 488022 205482 488050
rect 203904 484158 203932 488022
rect 203892 484152 203944 484158
rect 203892 484094 203944 484100
rect 203800 484084 203852 484090
rect 203800 484026 203852 484032
rect 203156 482384 203208 482390
rect 203156 482326 203208 482332
rect 203064 468512 203116 468518
rect 203064 468454 203116 468460
rect 202972 380452 203024 380458
rect 202972 380394 203024 380400
rect 202786 379536 202842 379545
rect 202786 379471 202842 379480
rect 202604 360256 202656 360262
rect 202604 360198 202656 360204
rect 202616 359514 202644 360198
rect 202604 359508 202656 359514
rect 202604 359450 202656 359456
rect 202512 272740 202564 272746
rect 202512 272682 202564 272688
rect 202420 271176 202472 271182
rect 202420 271118 202472 271124
rect 202328 166320 202380 166326
rect 202328 166262 202380 166268
rect 202236 70372 202288 70378
rect 202236 70314 202288 70320
rect 201316 59016 201368 59022
rect 201316 58958 201368 58964
rect 202800 58886 202828 379471
rect 203076 271794 203104 468454
rect 203168 376582 203196 482326
rect 203892 481160 203944 481166
rect 203892 481102 203944 481108
rect 203706 471472 203762 471481
rect 203706 471407 203762 471416
rect 203522 471336 203578 471345
rect 203522 471271 203578 471280
rect 203156 376576 203208 376582
rect 203156 376518 203208 376524
rect 203064 271788 203116 271794
rect 203064 271730 203116 271736
rect 202880 253904 202932 253910
rect 202880 253846 202932 253852
rect 202892 176662 202920 253846
rect 202880 176656 202932 176662
rect 202880 176598 202932 176604
rect 202892 176186 202920 176598
rect 202880 176180 202932 176186
rect 202880 176122 202932 176128
rect 203536 166802 203564 471271
rect 203614 466032 203670 466041
rect 203614 465967 203670 465976
rect 203524 166796 203576 166802
rect 203524 166738 203576 166744
rect 203628 166462 203656 465967
rect 203720 166734 203748 471407
rect 203800 466132 203852 466138
rect 203800 466074 203852 466080
rect 203812 282810 203840 466074
rect 203904 389162 203932 481102
rect 203984 465520 204036 465526
rect 203984 465462 204036 465468
rect 203892 389156 203944 389162
rect 203892 389098 203944 389104
rect 203890 380352 203946 380361
rect 203890 380287 203946 380296
rect 203904 358766 203932 380287
rect 203996 376582 204024 465462
rect 204272 379574 204300 488022
rect 204352 484152 204404 484158
rect 204732 484106 204760 488022
rect 204904 484900 204956 484906
rect 204904 484842 204956 484848
rect 204352 484094 204404 484100
rect 204364 413982 204392 484094
rect 204456 484078 204760 484106
rect 204456 476814 204484 484078
rect 204536 482316 204588 482322
rect 204536 482258 204588 482264
rect 204444 476808 204496 476814
rect 204444 476750 204496 476756
rect 204444 471504 204496 471510
rect 204444 471446 204496 471452
rect 204352 413976 204404 413982
rect 204352 413918 204404 413924
rect 204456 380662 204484 471446
rect 204444 380656 204496 380662
rect 204444 380598 204496 380604
rect 204548 380390 204576 482258
rect 204536 380384 204588 380390
rect 204536 380326 204588 380332
rect 204260 379568 204312 379574
rect 204260 379510 204312 379516
rect 204272 376718 204300 379510
rect 204810 378584 204866 378593
rect 204810 378519 204866 378528
rect 204824 378185 204852 378519
rect 204810 378176 204866 378185
rect 204810 378111 204866 378120
rect 204260 376712 204312 376718
rect 204260 376654 204312 376660
rect 203984 376576 204036 376582
rect 203984 376518 204036 376524
rect 203892 358760 203944 358766
rect 203892 358702 203944 358708
rect 203800 282804 203852 282810
rect 203800 282746 203852 282752
rect 203708 166728 203760 166734
rect 203708 166670 203760 166676
rect 204916 166666 204944 484842
rect 205192 484158 205220 488022
rect 205640 485648 205692 485654
rect 205638 485616 205640 485625
rect 205692 485616 205694 485625
rect 205638 485551 205694 485560
rect 205732 485580 205784 485586
rect 205732 485522 205784 485528
rect 205640 485444 205692 485450
rect 205640 485386 205692 485392
rect 205652 485217 205680 485386
rect 205638 485208 205694 485217
rect 205638 485143 205694 485152
rect 205744 484537 205772 485522
rect 205730 484528 205786 484537
rect 205730 484463 205786 484472
rect 205928 484430 205956 488036
rect 206020 488022 206402 488050
rect 206480 488022 206862 488050
rect 207246 488022 207520 488050
rect 205916 484424 205968 484430
rect 205916 484366 205968 484372
rect 205180 484152 205232 484158
rect 205180 484094 205232 484100
rect 205732 484152 205784 484158
rect 205732 484094 205784 484100
rect 205088 475448 205140 475454
rect 205088 475390 205140 475396
rect 204996 467356 205048 467362
rect 204996 467298 205048 467304
rect 205008 178022 205036 467298
rect 205100 271522 205128 475390
rect 205180 471980 205232 471986
rect 205180 471922 205232 471928
rect 205192 272678 205220 471922
rect 205272 466200 205324 466206
rect 205272 466142 205324 466148
rect 205284 273290 205312 466142
rect 205456 465724 205508 465730
rect 205456 465666 205508 465672
rect 205468 378185 205496 465666
rect 205744 416770 205772 484094
rect 205824 474020 205876 474026
rect 205824 473962 205876 473968
rect 205732 416764 205784 416770
rect 205732 416706 205784 416712
rect 205640 414724 205692 414730
rect 205640 414666 205692 414672
rect 205546 413944 205602 413953
rect 205546 413879 205602 413888
rect 205454 378176 205510 378185
rect 205454 378111 205510 378120
rect 205272 273284 205324 273290
rect 205272 273226 205324 273232
rect 205180 272672 205232 272678
rect 205180 272614 205232 272620
rect 205088 271516 205140 271522
rect 205088 271458 205140 271464
rect 204996 178016 205048 178022
rect 204996 177958 205048 177964
rect 204904 166660 204956 166666
rect 204904 166602 204956 166608
rect 203616 166456 203668 166462
rect 203616 166398 203668 166404
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204916 67658 204944 145522
rect 204904 67652 204956 67658
rect 204904 67594 204956 67600
rect 202788 58880 202840 58886
rect 202788 58822 202840 58828
rect 198648 58744 198700 58750
rect 198648 58686 198700 58692
rect 204916 57934 204944 67594
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 183192 57792 183244 57798
rect 183190 57760 183192 57769
rect 197360 57792 197412 57798
rect 183244 57760 183246 57769
rect 197360 57734 197412 57740
rect 183190 57695 183246 57704
rect 205560 57662 205588 413879
rect 205652 376310 205680 414666
rect 205732 378956 205784 378962
rect 205732 378898 205784 378904
rect 205744 378554 205772 378898
rect 205732 378548 205784 378554
rect 205732 378490 205784 378496
rect 205836 377534 205864 473962
rect 205916 465792 205968 465798
rect 205916 465734 205968 465740
rect 205928 380594 205956 465734
rect 206020 413302 206048 488022
rect 206480 484158 206508 488022
rect 206928 485376 206980 485382
rect 206928 485318 206980 485324
rect 206468 484152 206520 484158
rect 206468 484094 206520 484100
rect 206560 483744 206612 483750
rect 206560 483686 206612 483692
rect 206376 479528 206428 479534
rect 206376 479470 206428 479476
rect 206008 413296 206060 413302
rect 206008 413238 206060 413244
rect 206284 389224 206336 389230
rect 206284 389166 206336 389172
rect 205916 380588 205968 380594
rect 205916 380530 205968 380536
rect 206190 379536 206246 379545
rect 206190 379471 206246 379480
rect 205916 379092 205968 379098
rect 205916 379034 205968 379040
rect 205928 378282 205956 379034
rect 205916 378276 205968 378282
rect 205916 378218 205968 378224
rect 205824 377528 205876 377534
rect 205824 377470 205876 377476
rect 205640 376304 205692 376310
rect 205640 376246 205692 376252
rect 206204 58818 206232 379471
rect 206296 360262 206324 389166
rect 206284 360256 206336 360262
rect 206284 360198 206336 360204
rect 206388 165238 206416 479470
rect 206466 468888 206522 468897
rect 206466 468823 206522 468832
rect 206480 166530 206508 468823
rect 206572 271250 206600 483686
rect 206652 466404 206704 466410
rect 206652 466346 206704 466352
rect 206560 271244 206612 271250
rect 206560 271186 206612 271192
rect 206664 270473 206692 466346
rect 206744 464568 206796 464574
rect 206744 464510 206796 464516
rect 206756 272950 206784 464510
rect 206836 413976 206888 413982
rect 206836 413918 206888 413924
rect 206848 410582 206876 413918
rect 206836 410576 206888 410582
rect 206836 410518 206888 410524
rect 206836 378956 206888 378962
rect 206836 378898 206888 378904
rect 206744 272944 206796 272950
rect 206744 272886 206796 272892
rect 206650 270464 206706 270473
rect 206650 270399 206706 270408
rect 206848 268394 206876 378898
rect 206940 378282 206968 485318
rect 207112 484220 207164 484226
rect 207112 484162 207164 484168
rect 207020 466472 207072 466478
rect 207020 466414 207072 466420
rect 207032 390522 207060 466414
rect 207020 390516 207072 390522
rect 207020 390458 207072 390464
rect 207032 389230 207060 390458
rect 207020 389224 207072 389230
rect 207020 389166 207072 389172
rect 207124 383654 207152 484162
rect 207204 484152 207256 484158
rect 207204 484094 207256 484100
rect 207216 417450 207244 484094
rect 207296 474088 207348 474094
rect 207296 474030 207348 474036
rect 207204 417444 207256 417450
rect 207204 417386 207256 417392
rect 207204 416764 207256 416770
rect 207204 416706 207256 416712
rect 207216 414730 207244 416706
rect 207204 414724 207256 414730
rect 207204 414666 207256 414672
rect 207032 383626 207152 383654
rect 207032 380633 207060 383626
rect 207018 380624 207074 380633
rect 207018 380559 207020 380568
rect 207072 380559 207074 380568
rect 207020 380530 207072 380536
rect 207018 380216 207074 380225
rect 207018 380151 207074 380160
rect 207032 379710 207060 380151
rect 207020 379704 207072 379710
rect 207020 379646 207072 379652
rect 206928 378276 206980 378282
rect 206928 378218 206980 378224
rect 207308 377398 207336 474030
rect 207388 471436 207440 471442
rect 207388 471378 207440 471384
rect 207400 380118 207428 471378
rect 207492 466478 207520 488022
rect 207584 488022 207690 488050
rect 207768 488022 208150 488050
rect 208504 488022 208610 488050
rect 209086 488022 209360 488050
rect 207584 484158 207612 488022
rect 207664 484424 207716 484430
rect 207664 484366 207716 484372
rect 207572 484152 207624 484158
rect 207572 484094 207624 484100
rect 207676 475454 207704 484366
rect 207768 484226 207796 488022
rect 208216 485716 208268 485722
rect 208216 485658 208268 485664
rect 207756 484220 207808 484226
rect 207756 484162 207808 484168
rect 207664 475448 207716 475454
rect 207664 475390 207716 475396
rect 207756 474360 207808 474366
rect 207756 474302 207808 474308
rect 207664 468852 207716 468858
rect 207664 468794 207716 468800
rect 207480 466472 207532 466478
rect 207480 466414 207532 466420
rect 207388 380112 207440 380118
rect 207388 380054 207440 380060
rect 207296 377392 207348 377398
rect 207296 377334 207348 377340
rect 207020 375216 207072 375222
rect 207020 375158 207072 375164
rect 207032 374814 207060 375158
rect 207020 374808 207072 374814
rect 207020 374750 207072 374756
rect 206836 268388 206888 268394
rect 206836 268330 206888 268336
rect 207676 175234 207704 468794
rect 207768 271017 207796 474302
rect 207940 466472 207992 466478
rect 207940 466414 207992 466420
rect 207848 466336 207900 466342
rect 207848 466278 207900 466284
rect 207860 272610 207888 466278
rect 207952 422958 207980 466414
rect 207940 422952 207992 422958
rect 207940 422894 207992 422900
rect 208124 414860 208176 414866
rect 208124 414802 208176 414808
rect 207938 380624 207994 380633
rect 207938 380559 207994 380568
rect 207952 377641 207980 380559
rect 208030 378992 208086 379001
rect 208030 378927 208086 378936
rect 207938 377632 207994 377641
rect 207938 377567 207994 377576
rect 207848 272604 207900 272610
rect 207848 272546 207900 272552
rect 207754 271008 207810 271017
rect 207754 270943 207810 270952
rect 207952 268666 207980 377567
rect 208044 269793 208072 378927
rect 208136 374814 208164 414802
rect 208228 378826 208256 485658
rect 208400 485648 208452 485654
rect 208398 485616 208400 485625
rect 208452 485616 208454 485625
rect 208398 485551 208454 485560
rect 208400 484152 208452 484158
rect 208400 484094 208452 484100
rect 208412 380610 208440 484094
rect 208320 380582 208440 380610
rect 208320 380202 208348 380582
rect 208398 380488 208454 380497
rect 208504 380474 208532 488022
rect 209332 485450 209360 488022
rect 209320 485444 209372 485450
rect 209320 485386 209372 485392
rect 209424 484158 209452 488036
rect 209884 485790 209912 488036
rect 209976 488022 210358 488050
rect 210436 488022 210818 488050
rect 211202 488022 211476 488050
rect 211662 488022 211752 488050
rect 209780 485784 209832 485790
rect 209780 485726 209832 485732
rect 209872 485784 209924 485790
rect 209872 485726 209924 485732
rect 209792 485654 209820 485726
rect 209780 485648 209832 485654
rect 209780 485590 209832 485596
rect 209504 485308 209556 485314
rect 209504 485250 209556 485256
rect 209412 484152 209464 484158
rect 209412 484094 209464 484100
rect 209516 482746 209544 485250
rect 209976 484106 210004 488022
rect 209596 484084 209648 484090
rect 209596 484026 209648 484032
rect 209792 484078 210004 484106
rect 209424 482718 209544 482746
rect 209044 482656 209096 482662
rect 209044 482598 209096 482604
rect 208584 466608 208636 466614
rect 208584 466550 208636 466556
rect 208454 380446 208532 380474
rect 208398 380423 208454 380432
rect 208412 380390 208440 380423
rect 208400 380384 208452 380390
rect 208400 380326 208452 380332
rect 208320 380174 208440 380202
rect 208308 379704 208360 379710
rect 208308 379646 208360 379652
rect 208216 378820 208268 378826
rect 208216 378762 208268 378768
rect 208124 374808 208176 374814
rect 208124 374750 208176 374756
rect 208228 272542 208256 378762
rect 208320 375222 208348 379646
rect 208412 379506 208440 380174
rect 208400 379500 208452 379506
rect 208400 379442 208452 379448
rect 208412 378418 208440 379442
rect 208490 379128 208546 379137
rect 208490 379063 208546 379072
rect 208504 378457 208532 379063
rect 208490 378448 208546 378457
rect 208400 378412 208452 378418
rect 208490 378383 208546 378392
rect 208400 378354 208452 378360
rect 208308 375216 208360 375222
rect 208308 375158 208360 375164
rect 208596 359582 208624 466550
rect 208952 464772 209004 464778
rect 208952 464714 209004 464720
rect 208964 375970 208992 464714
rect 208952 375964 209004 375970
rect 208952 375906 209004 375912
rect 208584 359576 208636 359582
rect 208584 359518 208636 359524
rect 208216 272536 208268 272542
rect 208216 272478 208268 272484
rect 208030 269784 208086 269793
rect 208030 269719 208086 269728
rect 207940 268660 207992 268666
rect 207940 268602 207992 268608
rect 207664 175228 207716 175234
rect 207664 175170 207716 175176
rect 206468 166524 206520 166530
rect 206468 166466 206520 166472
rect 209056 165578 209084 482598
rect 209228 478304 209280 478310
rect 209228 478246 209280 478252
rect 209134 468752 209190 468761
rect 209134 468687 209190 468696
rect 209148 166394 209176 468687
rect 209240 271318 209268 478246
rect 209320 471776 209372 471782
rect 209320 471718 209372 471724
rect 209332 272882 209360 471718
rect 209424 379710 209452 482718
rect 209608 470594 209636 484026
rect 209516 470566 209636 470594
rect 209516 391950 209544 470566
rect 209504 391944 209556 391950
rect 209504 391886 209556 391892
rect 209686 390688 209742 390697
rect 209686 390623 209742 390632
rect 209412 379704 209464 379710
rect 209412 379646 209464 379652
rect 209502 379128 209558 379137
rect 209502 379063 209558 379072
rect 209410 378448 209466 378457
rect 209410 378383 209466 378392
rect 209320 272876 209372 272882
rect 209320 272818 209372 272824
rect 209228 271312 209280 271318
rect 209228 271254 209280 271260
rect 209318 269784 209374 269793
rect 209424 269754 209452 378383
rect 209318 269719 209374 269728
rect 209412 269748 209464 269754
rect 209136 166388 209188 166394
rect 209136 166330 209188 166336
rect 209044 165572 209096 165578
rect 209044 165514 209096 165520
rect 206376 165232 206428 165238
rect 206376 165174 206428 165180
rect 209332 144906 209360 269719
rect 209412 269690 209464 269696
rect 209516 268530 209544 379063
rect 209596 378480 209648 378486
rect 209596 378422 209648 378428
rect 209504 268524 209556 268530
rect 209504 268466 209556 268472
rect 209608 268462 209636 378422
rect 209596 268456 209648 268462
rect 209596 268398 209648 268404
rect 209320 144900 209372 144906
rect 209320 144842 209372 144848
rect 206192 58812 206244 58818
rect 206192 58754 206244 58760
rect 209700 57866 209728 390623
rect 209792 379370 209820 484078
rect 210436 483970 210464 488022
rect 211252 485648 211304 485654
rect 211252 485590 211304 485596
rect 211160 485580 211212 485586
rect 211160 485522 211212 485528
rect 211172 484945 211200 485522
rect 211158 484936 211214 484945
rect 211158 484871 211214 484880
rect 211264 484809 211292 485590
rect 211250 484800 211306 484809
rect 211250 484735 211306 484744
rect 211252 484152 211304 484158
rect 211252 484094 211304 484100
rect 209884 483942 210464 483970
rect 209780 379364 209832 379370
rect 209780 379306 209832 379312
rect 209884 379302 209912 483942
rect 210700 482724 210752 482730
rect 210700 482666 210752 482672
rect 210424 481024 210476 481030
rect 210424 480966 210476 480972
rect 210332 468988 210384 468994
rect 210332 468930 210384 468936
rect 210240 464840 210292 464846
rect 210240 464782 210292 464788
rect 209872 379296 209924 379302
rect 209872 379238 209924 379244
rect 210252 376446 210280 464782
rect 210240 376440 210292 376446
rect 210240 376382 210292 376388
rect 210344 273018 210372 468930
rect 210332 273012 210384 273018
rect 210332 272954 210384 272960
rect 210436 164966 210464 480966
rect 210516 472660 210568 472666
rect 210516 472602 210568 472608
rect 210528 165034 210556 472602
rect 210606 468616 210662 468625
rect 210606 468551 210662 468560
rect 210620 166598 210648 468551
rect 210712 271046 210740 482666
rect 210884 471708 210936 471714
rect 210884 471650 210936 471656
rect 210792 470008 210844 470014
rect 210792 469950 210844 469956
rect 210804 271454 210832 469950
rect 210896 272814 210924 471650
rect 211264 468314 211292 484094
rect 211252 468308 211304 468314
rect 211252 468250 211304 468256
rect 211068 379364 211120 379370
rect 211068 379306 211120 379312
rect 210974 379264 211030 379273
rect 210974 379199 211030 379208
rect 210884 272808 210936 272814
rect 210884 272750 210936 272756
rect 210884 272536 210936 272542
rect 210884 272478 210936 272484
rect 210896 271930 210924 272478
rect 210884 271924 210936 271930
rect 210884 271866 210936 271872
rect 210792 271448 210844 271454
rect 210792 271390 210844 271396
rect 210700 271040 210752 271046
rect 210700 270982 210752 270988
rect 210792 269748 210844 269754
rect 210792 269690 210844 269696
rect 210608 166592 210660 166598
rect 210608 166534 210660 166540
rect 210516 165028 210568 165034
rect 210516 164970 210568 164976
rect 210424 164960 210476 164966
rect 210424 164902 210476 164908
rect 210804 147558 210832 269690
rect 210792 147552 210844 147558
rect 210792 147494 210844 147500
rect 210896 145761 210924 271866
rect 210882 145752 210938 145761
rect 210882 145687 210938 145696
rect 210988 57934 211016 379199
rect 211080 379166 211108 379306
rect 211068 379160 211120 379166
rect 211068 379102 211120 379108
rect 211448 379098 211476 488022
rect 211724 484430 211752 488022
rect 211816 488022 212106 488050
rect 211712 484424 211764 484430
rect 211712 484366 211764 484372
rect 211816 484158 211844 488022
rect 212356 485172 212408 485178
rect 212356 485114 212408 485120
rect 211804 484152 211856 484158
rect 211804 484094 211856 484100
rect 211896 478236 211948 478242
rect 211896 478178 211948 478184
rect 211804 476876 211856 476882
rect 211804 476818 211856 476824
rect 211528 471164 211580 471170
rect 211528 471106 211580 471112
rect 211436 379092 211488 379098
rect 211436 379034 211488 379040
rect 211066 378584 211122 378593
rect 211066 378519 211122 378528
rect 210976 57928 211028 57934
rect 210976 57870 211028 57876
rect 209688 57860 209740 57866
rect 209688 57802 209740 57808
rect 205548 57656 205600 57662
rect 157338 57624 157394 57633
rect 157338 57559 157394 57568
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 165618 57624 165674 57633
rect 205548 57598 205600 57604
rect 165618 57559 165674 57568
rect 153290 56400 153346 56409
rect 153290 56335 153346 56344
rect 119066 56128 119122 56137
rect 119066 56063 119122 56072
rect 116124 55140 116176 55146
rect 116124 55082 116176 55088
rect 110420 55072 110472 55078
rect 157352 55049 157380 57559
rect 110420 55014 110472 55020
rect 157338 55040 157394 55049
rect 157338 54975 157394 54984
rect 106280 54936 106332 54942
rect 160112 54913 160140 57559
rect 165632 55185 165660 57559
rect 211080 57458 211108 378519
rect 211434 377904 211490 377913
rect 211434 377839 211490 377848
rect 211448 377641 211476 377839
rect 211434 377632 211490 377641
rect 211434 377567 211490 377576
rect 211540 376242 211568 471106
rect 211620 378412 211672 378418
rect 211620 378354 211672 378360
rect 211528 376236 211580 376242
rect 211528 376178 211580 376184
rect 211632 270434 211660 378354
rect 211712 378276 211764 378282
rect 211712 378218 211764 378224
rect 211724 270502 211752 378218
rect 211712 270496 211764 270502
rect 211712 270438 211764 270444
rect 211620 270428 211672 270434
rect 211620 270370 211672 270376
rect 211068 57452 211120 57458
rect 211068 57394 211120 57400
rect 211816 57322 211844 476818
rect 211908 165374 211936 478178
rect 212080 476944 212132 476950
rect 212080 476886 212132 476892
rect 211986 471608 212042 471617
rect 211986 471543 212042 471552
rect 211896 165368 211948 165374
rect 211896 165310 211948 165316
rect 212000 164218 212028 471543
rect 212092 271794 212120 476886
rect 212172 468920 212224 468926
rect 212172 468862 212224 468868
rect 212080 271788 212132 271794
rect 212080 271730 212132 271736
rect 212184 271114 212212 468862
rect 212264 464500 212316 464506
rect 212264 464442 212316 464448
rect 212276 272542 212304 464442
rect 212368 377398 212396 485114
rect 212448 465792 212500 465798
rect 212448 465734 212500 465740
rect 212460 378593 212488 465734
rect 212552 379914 212580 488036
rect 212736 488022 213026 488050
rect 212632 484152 212684 484158
rect 212632 484094 212684 484100
rect 212644 380633 212672 484094
rect 212630 380624 212686 380633
rect 212630 380559 212686 380568
rect 212540 379908 212592 379914
rect 212540 379850 212592 379856
rect 212446 378584 212502 378593
rect 212446 378519 212502 378528
rect 212460 378321 212488 378519
rect 212446 378312 212502 378321
rect 212446 378247 212502 378256
rect 212446 377904 212502 377913
rect 212446 377839 212502 377848
rect 212356 377392 212408 377398
rect 212356 377334 212408 377340
rect 212354 376680 212410 376689
rect 212354 376615 212410 376624
rect 212264 272536 212316 272542
rect 212264 272478 212316 272484
rect 212172 271108 212224 271114
rect 212172 271050 212224 271056
rect 212172 270496 212224 270502
rect 212172 270438 212224 270444
rect 212184 269618 212212 270438
rect 212262 270056 212318 270065
rect 212262 269991 212318 270000
rect 212172 269612 212224 269618
rect 212172 269554 212224 269560
rect 212080 268388 212132 268394
rect 212080 268330 212132 268336
rect 211988 164212 212040 164218
rect 211988 164154 212040 164160
rect 212092 148374 212120 268330
rect 212080 148368 212132 148374
rect 212080 148310 212132 148316
rect 212184 147626 212212 269554
rect 212276 148646 212304 269991
rect 212264 148640 212316 148646
rect 212264 148582 212316 148588
rect 212172 147620 212224 147626
rect 212172 147562 212224 147568
rect 212368 58954 212396 376615
rect 212460 59090 212488 377839
rect 212552 376174 212580 379850
rect 212736 379710 212764 488022
rect 213380 484430 213408 488036
rect 213472 488022 213854 488050
rect 214024 488022 214314 488050
rect 214790 488022 214880 488050
rect 212816 484424 212868 484430
rect 212816 484366 212868 484372
rect 213368 484424 213420 484430
rect 213368 484366 213420 484372
rect 212724 379704 212776 379710
rect 212724 379646 212776 379652
rect 212736 377641 212764 379646
rect 212828 379438 212856 484366
rect 213472 484158 213500 488022
rect 213460 484152 213512 484158
rect 213460 484094 213512 484100
rect 213920 484152 213972 484158
rect 213920 484094 213972 484100
rect 213368 471232 213420 471238
rect 213368 471174 213420 471180
rect 213184 467424 213236 467430
rect 213184 467366 213236 467372
rect 212908 467220 212960 467226
rect 212908 467162 212960 467168
rect 212920 381041 212948 467162
rect 213092 465656 213144 465662
rect 213092 465598 213144 465604
rect 212906 381032 212962 381041
rect 212906 380967 212962 380976
rect 212816 379432 212868 379438
rect 212816 379374 212868 379380
rect 212722 377632 212778 377641
rect 212722 377567 212778 377576
rect 213104 376718 213132 465598
rect 213092 376712 213144 376718
rect 213092 376654 213144 376660
rect 212540 376168 212592 376174
rect 212540 376110 212592 376116
rect 212908 274712 212960 274718
rect 212908 274654 212960 274660
rect 212920 148442 212948 274654
rect 213196 271862 213224 467366
rect 213274 377632 213330 377641
rect 213274 377567 213330 377576
rect 213184 271856 213236 271862
rect 213184 271798 213236 271804
rect 213092 270428 213144 270434
rect 213092 270370 213144 270376
rect 213104 269890 213132 270370
rect 213092 269884 213144 269890
rect 213092 269826 213144 269832
rect 212908 148436 212960 148442
rect 212908 148378 212960 148384
rect 213000 147756 213052 147762
rect 213000 147698 213052 147704
rect 212448 59084 212500 59090
rect 212448 59026 212500 59032
rect 212356 58948 212408 58954
rect 212356 58890 212408 58896
rect 211804 57316 211856 57322
rect 211804 57258 211856 57264
rect 213012 55758 213040 147698
rect 213104 144770 213132 269826
rect 213288 268938 213316 377567
rect 213380 376310 213408 471174
rect 213736 380588 213788 380594
rect 213736 380530 213788 380536
rect 213748 379846 213776 380530
rect 213828 380520 213880 380526
rect 213828 380462 213880 380468
rect 213840 380050 213868 380462
rect 213828 380044 213880 380050
rect 213828 379986 213880 379992
rect 213736 379840 213788 379846
rect 213736 379782 213788 379788
rect 213748 379624 213776 379782
rect 213564 379596 213776 379624
rect 213460 378752 213512 378758
rect 213460 378694 213512 378700
rect 213368 376304 213420 376310
rect 213368 376246 213420 376252
rect 213472 273426 213500 378694
rect 213460 273420 213512 273426
rect 213460 273362 213512 273368
rect 213564 269006 213592 379596
rect 213840 379522 213868 379986
rect 213748 379494 213868 379522
rect 213644 378616 213696 378622
rect 213644 378558 213696 378564
rect 213656 270434 213684 378558
rect 213748 271998 213776 379494
rect 213828 379432 213880 379438
rect 213828 379374 213880 379380
rect 213840 379234 213868 379374
rect 213828 379228 213880 379234
rect 213828 379170 213880 379176
rect 213826 377904 213882 377913
rect 213826 377839 213882 377848
rect 213736 271992 213788 271998
rect 213736 271934 213788 271940
rect 213644 270428 213696 270434
rect 213644 270370 213696 270376
rect 213552 269000 213604 269006
rect 213552 268942 213604 268948
rect 213276 268932 213328 268938
rect 213276 268874 213328 268880
rect 213460 268524 213512 268530
rect 213460 268466 213512 268472
rect 213368 268456 213420 268462
rect 213368 268398 213420 268404
rect 213184 148708 213236 148714
rect 213184 148650 213236 148656
rect 213196 147558 213224 148650
rect 213380 148578 213408 268398
rect 213368 148572 213420 148578
rect 213368 148514 213420 148520
rect 213184 147552 213236 147558
rect 213184 147494 213236 147500
rect 213092 144764 213144 144770
rect 213092 144706 213144 144712
rect 213196 55894 213224 147494
rect 213274 145888 213330 145897
rect 213274 145823 213330 145832
rect 213288 144906 213316 145823
rect 213276 144900 213328 144906
rect 213276 144842 213328 144848
rect 213184 55888 213236 55894
rect 213184 55830 213236 55836
rect 213000 55752 213052 55758
rect 213000 55694 213052 55700
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 106280 54878 106332 54884
rect 160098 54904 160154 54913
rect 160098 54839 160154 54848
rect 91468 54732 91520 54738
rect 91468 54674 91520 54680
rect 81440 54664 81492 54670
rect 81440 54606 81492 54612
rect 78680 54596 78732 54602
rect 78680 54538 78732 54544
rect 213288 54398 213316 144842
rect 213472 144838 213500 268466
rect 213564 144906 213592 268942
rect 213736 148368 213788 148374
rect 213736 148310 213788 148316
rect 213644 147688 213696 147694
rect 213644 147630 213696 147636
rect 213552 144900 213604 144906
rect 213552 144842 213604 144848
rect 213460 144832 213512 144838
rect 213460 144774 213512 144780
rect 213276 54392 213328 54398
rect 213276 54334 213328 54340
rect 213656 54330 213684 147630
rect 213748 55146 213776 148310
rect 213840 57594 213868 377839
rect 213932 375358 213960 484094
rect 214024 376174 214052 488022
rect 214852 484537 214880 488022
rect 214944 488022 215234 488050
rect 215312 488022 215602 488050
rect 215680 488022 216062 488050
rect 216232 488022 216522 488050
rect 216998 488022 217088 488050
rect 214838 484528 214894 484537
rect 214838 484463 214894 484472
rect 214944 484158 214972 488022
rect 215024 484424 215076 484430
rect 215024 484366 215076 484372
rect 214932 484152 214984 484158
rect 214932 484094 214984 484100
rect 214840 481092 214892 481098
rect 214840 481034 214892 481040
rect 214564 474156 214616 474162
rect 214564 474098 214616 474104
rect 214380 468444 214432 468450
rect 214380 468386 214432 468392
rect 214392 376378 214420 468386
rect 214472 376508 214524 376514
rect 214472 376450 214524 376456
rect 214380 376372 214432 376378
rect 214380 376314 214432 376320
rect 214012 376168 214064 376174
rect 214012 376110 214064 376116
rect 214024 375902 214052 376110
rect 214012 375896 214064 375902
rect 214012 375838 214064 375844
rect 213920 375352 213972 375358
rect 213920 375294 213972 375300
rect 213932 375154 213960 375294
rect 213920 375148 213972 375154
rect 213920 375090 213972 375096
rect 214380 358556 214432 358562
rect 214380 358498 214432 358504
rect 214392 270337 214420 358498
rect 214378 270328 214434 270337
rect 214378 270263 214434 270272
rect 214484 269074 214512 376450
rect 214472 269068 214524 269074
rect 214472 269010 214524 269016
rect 214472 251932 214524 251938
rect 214472 251874 214524 251880
rect 214484 162722 214512 251874
rect 214576 165442 214604 474098
rect 214656 472728 214708 472734
rect 214656 472670 214708 472676
rect 214668 165510 214696 472670
rect 214746 471200 214802 471209
rect 214746 471135 214802 471144
rect 214760 166870 214788 471135
rect 214852 271658 214880 481034
rect 214932 474292 214984 474298
rect 214932 474234 214984 474240
rect 214840 271652 214892 271658
rect 214840 271594 214892 271600
rect 214944 271590 214972 474234
rect 215036 379778 215064 484366
rect 215116 469056 215168 469062
rect 215116 468998 215168 469004
rect 215024 379772 215076 379778
rect 215024 379714 215076 379720
rect 215036 376514 215064 379714
rect 215024 376508 215076 376514
rect 215024 376450 215076 376456
rect 215128 375902 215156 468998
rect 215312 380066 215340 488022
rect 215680 484106 215708 488022
rect 215496 484078 215708 484106
rect 215496 380769 215524 484078
rect 216232 480254 216260 488022
rect 217060 484430 217088 488022
rect 217152 488022 217442 488050
rect 217048 484424 217100 484430
rect 217048 484366 217100 484372
rect 215588 480226 216260 480254
rect 215588 402974 215616 480226
rect 216036 478372 216088 478378
rect 216036 478314 216088 478320
rect 215852 469192 215904 469198
rect 215852 469134 215904 469140
rect 215588 402946 215708 402974
rect 215482 380760 215538 380769
rect 215482 380695 215538 380704
rect 215312 380038 215524 380066
rect 215300 379976 215352 379982
rect 215300 379918 215352 379924
rect 215312 379574 215340 379918
rect 215300 379568 215352 379574
rect 215300 379510 215352 379516
rect 215392 379432 215444 379438
rect 215392 379374 215444 379380
rect 215404 378350 215432 379374
rect 215392 378344 215444 378350
rect 215392 378286 215444 378292
rect 215206 376680 215262 376689
rect 215206 376615 215262 376624
rect 215116 375896 215168 375902
rect 215116 375838 215168 375844
rect 215116 375284 215168 375290
rect 215116 375226 215168 375232
rect 215128 374746 215156 375226
rect 215116 374740 215168 374746
rect 215116 374682 215168 374688
rect 215024 273420 215076 273426
rect 215024 273362 215076 273368
rect 214932 271584 214984 271590
rect 214932 271526 214984 271532
rect 214930 270328 214986 270337
rect 214930 270263 214986 270272
rect 214840 251864 214892 251870
rect 214840 251806 214892 251812
rect 214748 166864 214800 166870
rect 214748 166806 214800 166812
rect 214656 165504 214708 165510
rect 214656 165446 214708 165452
rect 214564 165436 214616 165442
rect 214564 165378 214616 165384
rect 214472 162716 214524 162722
rect 214472 162658 214524 162664
rect 214484 59158 214512 162658
rect 214852 162654 214880 251806
rect 214840 162648 214892 162654
rect 214840 162590 214892 162596
rect 214852 161474 214880 162590
rect 214760 161446 214880 161474
rect 214564 148640 214616 148646
rect 214564 148582 214616 148588
rect 214472 59152 214524 59158
rect 214472 59094 214524 59100
rect 213828 57588 213880 57594
rect 213828 57530 213880 57536
rect 214576 56574 214604 148582
rect 214656 148572 214708 148578
rect 214656 148514 214708 148520
rect 214564 56568 214616 56574
rect 214564 56510 214616 56516
rect 214668 56370 214696 148514
rect 214760 59226 214788 161446
rect 214944 148918 214972 270263
rect 215036 148986 215064 273362
rect 215128 270502 215156 374682
rect 215116 270496 215168 270502
rect 215116 270438 215168 270444
rect 215116 268252 215168 268258
rect 215116 268194 215168 268200
rect 215024 148980 215076 148986
rect 215024 148922 215076 148928
rect 214932 148912 214984 148918
rect 214932 148854 214984 148860
rect 214840 148436 214892 148442
rect 214840 148378 214892 148384
rect 214852 147506 214880 148378
rect 214944 147694 214972 148854
rect 215036 147762 215064 148922
rect 215024 147756 215076 147762
rect 215024 147698 215076 147704
rect 214932 147688 214984 147694
rect 214932 147630 214984 147636
rect 214852 147478 215064 147506
rect 214930 145616 214986 145625
rect 214930 145551 214986 145560
rect 214944 144838 214972 145551
rect 214932 144832 214984 144838
rect 214932 144774 214984 144780
rect 214748 59220 214800 59226
rect 214748 59162 214800 59168
rect 214656 56364 214708 56370
rect 214656 56306 214708 56312
rect 214944 55185 214972 144774
rect 215036 56438 215064 147478
rect 215128 145858 215156 268194
rect 215116 145852 215168 145858
rect 215116 145794 215168 145800
rect 215024 56432 215076 56438
rect 215024 56374 215076 56380
rect 214930 55176 214986 55185
rect 213736 55140 213788 55146
rect 214930 55111 214986 55120
rect 213736 55082 213788 55088
rect 215128 54602 215156 145794
rect 215220 57798 215248 376615
rect 215404 274718 215432 378286
rect 215496 375290 215524 380038
rect 215574 377904 215630 377913
rect 215574 377839 215630 377848
rect 215484 375284 215536 375290
rect 215484 375226 215536 375232
rect 215588 277386 215616 377839
rect 215680 377777 215708 402946
rect 215666 377768 215722 377777
rect 215666 377703 215722 377712
rect 215864 376514 215892 469134
rect 215944 468784 215996 468790
rect 215944 468726 215996 468732
rect 215852 376508 215904 376514
rect 215852 376450 215904 376456
rect 215668 358148 215720 358154
rect 215668 358090 215720 358096
rect 215496 277358 215616 277386
rect 215392 274712 215444 274718
rect 215392 274654 215444 274660
rect 215404 273494 215432 274654
rect 215392 273488 215444 273494
rect 215392 273430 215444 273436
rect 215496 273170 215524 277358
rect 215404 273142 215524 273170
rect 215404 267734 215432 273142
rect 215680 271810 215708 358090
rect 215852 357536 215904 357542
rect 215852 357478 215904 357484
rect 215864 277394 215892 357478
rect 215772 277366 215892 277394
rect 215772 273358 215800 277366
rect 215760 273352 215812 273358
rect 215760 273294 215812 273300
rect 215588 271782 215708 271810
rect 215588 270065 215616 271782
rect 215668 270428 215720 270434
rect 215668 270370 215720 270376
rect 215574 270056 215630 270065
rect 215574 269991 215630 270000
rect 215680 269958 215708 270370
rect 215668 269952 215720 269958
rect 215668 269894 215720 269900
rect 215404 267706 215616 267734
rect 215208 57792 215260 57798
rect 215208 57734 215260 57740
rect 215588 57526 215616 267706
rect 215680 145654 215708 269894
rect 215772 149054 215800 273294
rect 215852 268932 215904 268938
rect 215852 268874 215904 268880
rect 215864 268734 215892 268874
rect 215852 268728 215904 268734
rect 215852 268670 215904 268676
rect 215864 161474 215892 268670
rect 215956 165102 215984 468726
rect 216048 271697 216076 478314
rect 216220 471912 216272 471918
rect 216220 471854 216272 471860
rect 216128 466064 216180 466070
rect 216128 466006 216180 466012
rect 216034 271688 216090 271697
rect 216034 271623 216090 271632
rect 216140 270978 216168 466006
rect 216232 376038 216260 471854
rect 217152 470594 217180 488022
rect 217796 485722 217824 488036
rect 218072 488022 218270 488050
rect 217784 485716 217836 485722
rect 217784 485658 217836 485664
rect 217508 485240 217560 485246
rect 217508 485182 217560 485188
rect 217416 485104 217468 485110
rect 217416 485046 217468 485052
rect 217324 476808 217376 476814
rect 217324 476750 217376 476756
rect 216876 470566 217180 470594
rect 216678 417888 216734 417897
rect 216678 417823 216734 417832
rect 216692 417450 216720 417823
rect 216680 417444 216732 417450
rect 216680 417386 216732 417392
rect 216692 412634 216720 417386
rect 216876 414866 216904 470566
rect 216864 414860 216916 414866
rect 216864 414802 216916 414808
rect 217046 414760 217102 414769
rect 217046 414695 217048 414704
rect 217100 414695 217102 414704
rect 217048 414666 217100 414672
rect 216862 413808 216918 413817
rect 216862 413743 216918 413752
rect 216876 413302 216904 413743
rect 216864 413296 216916 413302
rect 216864 413238 216916 413244
rect 216692 412606 216812 412634
rect 216678 410952 216734 410961
rect 216678 410887 216734 410896
rect 216692 410582 216720 410887
rect 216680 410576 216732 410582
rect 216680 410518 216732 410524
rect 216680 407516 216732 407522
rect 216680 407458 216732 407464
rect 216692 398154 216720 407458
rect 216784 398274 216812 412606
rect 216772 398268 216824 398274
rect 216772 398210 216824 398216
rect 216692 398126 216812 398154
rect 216680 398064 216732 398070
rect 216680 398006 216732 398012
rect 216692 392086 216720 398006
rect 216680 392080 216732 392086
rect 216680 392022 216732 392028
rect 216680 391944 216732 391950
rect 216680 391886 216732 391892
rect 216692 390969 216720 391886
rect 216678 390960 216734 390969
rect 216678 390895 216734 390904
rect 216680 390516 216732 390522
rect 216680 390458 216732 390464
rect 216692 389337 216720 390458
rect 216678 389328 216734 389337
rect 216678 389263 216734 389272
rect 216680 389156 216732 389162
rect 216680 389098 216732 389104
rect 216692 389065 216720 389098
rect 216678 389056 216734 389065
rect 216678 388991 216734 389000
rect 216784 388498 216812 398126
rect 216692 388470 216812 388498
rect 216692 380866 216720 388470
rect 216772 388408 216824 388414
rect 216772 388350 216824 388356
rect 216680 380860 216732 380866
rect 216680 380802 216732 380808
rect 216586 380760 216642 380769
rect 216586 380695 216642 380704
rect 216404 379976 216456 379982
rect 216404 379918 216456 379924
rect 216312 376168 216364 376174
rect 216312 376110 216364 376116
rect 216220 376032 216272 376038
rect 216220 375974 216272 375980
rect 216324 375630 216352 376110
rect 216312 375624 216364 375630
rect 216312 375566 216364 375572
rect 216220 271992 216272 271998
rect 216220 271934 216272 271940
rect 216128 270972 216180 270978
rect 216128 270914 216180 270920
rect 216036 269068 216088 269074
rect 216036 269010 216088 269016
rect 216048 268598 216076 269010
rect 216036 268592 216088 268598
rect 216036 268534 216088 268540
rect 215944 165096 215996 165102
rect 215944 165038 215996 165044
rect 216048 162858 216076 268534
rect 216232 164014 216260 271934
rect 216324 268326 216352 375566
rect 216416 271425 216444 379918
rect 216494 376680 216550 376689
rect 216494 376615 216550 376624
rect 216508 375698 216536 376615
rect 216600 375766 216628 380695
rect 216588 375760 216640 375766
rect 216588 375702 216640 375708
rect 216496 375692 216548 375698
rect 216496 375634 216548 375640
rect 216402 271416 216458 271425
rect 216402 271351 216458 271360
rect 216404 270496 216456 270502
rect 216404 270438 216456 270444
rect 216416 269550 216444 270438
rect 216404 269544 216456 269550
rect 216404 269486 216456 269492
rect 216312 268320 216364 268326
rect 216312 268262 216364 268268
rect 216220 164008 216272 164014
rect 216220 163950 216272 163956
rect 216036 162852 216088 162858
rect 216036 162794 216088 162800
rect 216220 161560 216272 161566
rect 216220 161502 216272 161508
rect 216232 161474 216260 161502
rect 215864 161446 216260 161474
rect 215760 149048 215812 149054
rect 215760 148990 215812 148996
rect 215852 148504 215904 148510
rect 215852 148446 215904 148452
rect 215864 147642 215892 148446
rect 215864 147626 215984 147642
rect 215852 147620 215984 147626
rect 215904 147614 215984 147620
rect 215852 147562 215904 147568
rect 215864 147531 215892 147562
rect 215668 145648 215720 145654
rect 215668 145590 215720 145596
rect 215850 145072 215906 145081
rect 215850 145007 215906 145016
rect 215864 59430 215892 145007
rect 215852 59424 215904 59430
rect 215852 59366 215904 59372
rect 215576 57520 215628 57526
rect 215576 57462 215628 57468
rect 215956 55078 215984 147614
rect 216128 145716 216180 145722
rect 216128 145658 216180 145664
rect 216036 144900 216088 144906
rect 216036 144842 216088 144848
rect 215944 55072 215996 55078
rect 215944 55014 215996 55020
rect 215116 54596 215168 54602
rect 215116 54538 215168 54544
rect 216048 54466 216076 144842
rect 216140 56030 216168 145658
rect 216232 59634 216260 161446
rect 216416 146169 216444 269486
rect 216508 268870 216536 375634
rect 216692 309097 216720 380802
rect 216784 378078 216812 388350
rect 216876 380798 216904 413238
rect 216956 410576 217008 410582
rect 216956 410518 217008 410524
rect 216864 380792 216916 380798
rect 216864 380734 216916 380740
rect 216772 378072 216824 378078
rect 216772 378014 216824 378020
rect 216678 309088 216734 309097
rect 216678 309023 216734 309032
rect 216876 307737 216904 380734
rect 216968 380730 216996 410518
rect 217060 407522 217088 414666
rect 217336 409193 217364 476750
rect 217322 409184 217378 409193
rect 217322 409119 217378 409128
rect 217048 407516 217100 407522
rect 217048 407458 217100 407464
rect 217048 392080 217100 392086
rect 217048 392022 217100 392028
rect 217060 388414 217088 392022
rect 217048 388408 217100 388414
rect 217048 388350 217100 388356
rect 216956 380724 217008 380730
rect 216956 380666 217008 380672
rect 216968 379574 216996 380666
rect 216956 379568 217008 379574
rect 216956 379510 217008 379516
rect 217138 379536 217194 379545
rect 217138 379471 217194 379480
rect 217048 358624 217100 358630
rect 217048 358566 217100 358572
rect 216954 309904 217010 309913
rect 216954 309839 217010 309848
rect 216862 307728 216918 307737
rect 216862 307663 216918 307672
rect 216680 284300 216732 284306
rect 216680 284242 216732 284248
rect 216692 284073 216720 284242
rect 216678 284064 216734 284073
rect 216678 283999 216734 284008
rect 216680 282872 216732 282878
rect 216680 282814 216732 282820
rect 216692 282441 216720 282814
rect 216772 282804 216824 282810
rect 216772 282746 216824 282752
rect 216678 282432 216734 282441
rect 216678 282367 216734 282376
rect 216784 282169 216812 282746
rect 216770 282160 216826 282169
rect 216770 282095 216826 282104
rect 216586 271416 216642 271425
rect 216586 271351 216642 271360
rect 216496 268864 216548 268870
rect 216496 268806 216548 268812
rect 216600 164082 216628 271351
rect 216680 270428 216732 270434
rect 216680 270370 216732 270376
rect 216692 176746 216720 270370
rect 216862 270328 216918 270337
rect 216862 270263 216918 270272
rect 216772 270156 216824 270162
rect 216772 270098 216824 270104
rect 216784 176866 216812 270098
rect 216876 270065 216904 270263
rect 216862 270056 216918 270065
rect 216862 269991 216918 270000
rect 216862 203960 216918 203969
rect 216862 203895 216918 203904
rect 216772 176860 216824 176866
rect 216772 176802 216824 176808
rect 216692 176718 216812 176746
rect 216680 176656 216732 176662
rect 216680 176598 216732 176604
rect 216692 175409 216720 176598
rect 216678 175400 216734 175409
rect 216678 175335 216734 175344
rect 216784 175250 216812 176718
rect 216692 175222 216812 175250
rect 216588 164076 216640 164082
rect 216588 164018 216640 164024
rect 216692 163538 216720 175222
rect 216772 175160 216824 175166
rect 216772 175102 216824 175108
rect 216680 163532 216732 163538
rect 216680 163474 216732 163480
rect 216496 149048 216548 149054
rect 216496 148990 216548 148996
rect 216402 146160 216458 146169
rect 216402 146095 216458 146104
rect 216312 145648 216364 145654
rect 216312 145590 216364 145596
rect 216324 145382 216352 145590
rect 216312 145376 216364 145382
rect 216312 145318 216364 145324
rect 216220 59628 216272 59634
rect 216220 59570 216272 59576
rect 216128 56024 216180 56030
rect 216128 55966 216180 55972
rect 216324 55962 216352 145318
rect 216416 145081 216444 146095
rect 216402 145072 216458 145081
rect 216402 145007 216458 145016
rect 216404 144968 216456 144974
rect 216404 144910 216456 144916
rect 216312 55956 216364 55962
rect 216312 55898 216364 55904
rect 216416 54670 216444 144910
rect 216508 55214 216536 148990
rect 216588 145648 216640 145654
rect 216588 145590 216640 145596
rect 216600 144906 216628 145590
rect 216784 145178 216812 175102
rect 216772 145172 216824 145178
rect 216772 145114 216824 145120
rect 216588 144900 216640 144906
rect 216588 144842 216640 144848
rect 216876 96937 216904 203895
rect 216968 203017 216996 309839
rect 217060 270094 217088 358566
rect 217152 302161 217180 379471
rect 217324 378072 217376 378078
rect 217324 378014 217376 378020
rect 217336 377330 217364 378014
rect 217428 377534 217456 485046
rect 217520 378078 217548 485182
rect 217692 475448 217744 475454
rect 217692 475390 217744 475396
rect 217600 466268 217652 466274
rect 217600 466210 217652 466216
rect 217612 380934 217640 466210
rect 217704 412049 217732 475390
rect 217784 469124 217836 469130
rect 217784 469066 217836 469072
rect 217690 412040 217746 412049
rect 217690 411975 217746 411984
rect 217600 380928 217652 380934
rect 217600 380870 217652 380876
rect 217600 379568 217652 379574
rect 217600 379510 217652 379516
rect 217508 378072 217560 378078
rect 217508 378014 217560 378020
rect 217416 377528 217468 377534
rect 217416 377470 217468 377476
rect 217324 377324 217376 377330
rect 217324 377266 217376 377272
rect 217232 375760 217284 375766
rect 217232 375702 217284 375708
rect 217138 302152 217194 302161
rect 217138 302087 217194 302096
rect 217048 270088 217100 270094
rect 217048 270030 217100 270036
rect 216954 203008 217010 203017
rect 216954 202943 217010 202952
rect 216862 96928 216918 96937
rect 216862 96863 216918 96872
rect 216968 95985 216996 202943
rect 217152 195265 217180 302087
rect 217244 270434 217272 375702
rect 217336 311001 217364 377266
rect 217508 375148 217560 375154
rect 217508 375090 217560 375096
rect 217520 375057 217548 375090
rect 217506 375048 217562 375057
rect 217506 374983 217562 374992
rect 217322 310992 217378 311001
rect 217322 310927 217378 310936
rect 217506 310992 217562 311001
rect 217506 310927 217562 310936
rect 217414 307728 217470 307737
rect 217414 307663 217470 307672
rect 217428 306785 217456 307663
rect 217414 306776 217470 306785
rect 217414 306711 217470 306720
rect 217232 270428 217284 270434
rect 217232 270370 217284 270376
rect 217428 199889 217456 306711
rect 217520 203969 217548 310927
rect 217612 303929 217640 379510
rect 217704 377058 217732 411975
rect 217796 411466 217824 469066
rect 217968 422952 218020 422958
rect 217968 422894 218020 422900
rect 217980 416945 218008 422894
rect 217966 416936 218022 416945
rect 217966 416871 218022 416880
rect 217784 411460 217836 411466
rect 217784 411402 217836 411408
rect 217874 409184 217930 409193
rect 217874 409119 217930 409128
rect 217888 380905 217916 409119
rect 217874 380896 217930 380905
rect 217874 380831 217930 380840
rect 217784 379908 217836 379914
rect 217784 379850 217836 379856
rect 217796 379642 217824 379850
rect 217784 379636 217836 379642
rect 217784 379578 217836 379584
rect 217888 379545 217916 380831
rect 217874 379536 217930 379545
rect 217874 379471 217930 379480
rect 217692 377052 217744 377058
rect 217692 376994 217744 377000
rect 217704 373994 217732 376994
rect 217876 374808 217928 374814
rect 217876 374750 217928 374756
rect 217704 373966 217824 373994
rect 217690 309088 217746 309097
rect 217690 309023 217746 309032
rect 217704 307873 217732 309023
rect 217690 307864 217746 307873
rect 217690 307799 217746 307808
rect 217598 303920 217654 303929
rect 217598 303855 217654 303864
rect 217506 203960 217562 203969
rect 217506 203895 217562 203904
rect 217414 199880 217470 199889
rect 217414 199815 217470 199824
rect 217230 197024 217286 197033
rect 217230 196959 217286 196968
rect 217138 195256 217194 195265
rect 217138 195191 217194 195200
rect 217048 178016 217100 178022
rect 217048 177958 217100 177964
rect 217060 177041 217088 177958
rect 217046 177032 217102 177041
rect 217046 176967 217102 176976
rect 217048 176860 217100 176866
rect 217048 176802 217100 176808
rect 217060 175166 217088 176802
rect 217140 175228 217192 175234
rect 217140 175170 217192 175176
rect 217048 175160 217100 175166
rect 217152 175137 217180 175170
rect 217048 175102 217100 175108
rect 217138 175128 217194 175137
rect 217138 175063 217194 175072
rect 217140 162852 217192 162858
rect 217140 162794 217192 162800
rect 217152 161498 217180 162794
rect 217140 161492 217192 161498
rect 217140 161434 217192 161440
rect 217048 145580 217100 145586
rect 217048 145522 217100 145528
rect 216954 95976 217010 95985
rect 216954 95911 217010 95920
rect 216680 70372 216732 70378
rect 216680 70314 216732 70320
rect 216692 70009 216720 70314
rect 216678 70000 216734 70009
rect 216678 69935 216734 69944
rect 216678 68368 216734 68377
rect 216678 68303 216734 68312
rect 216692 67658 216720 68303
rect 216680 67652 216732 67658
rect 216680 67594 216732 67600
rect 216496 55208 216548 55214
rect 216496 55150 216548 55156
rect 217060 54806 217088 145522
rect 217152 59566 217180 161434
rect 217244 90001 217272 196959
rect 217428 92857 217456 199815
rect 217506 197432 217562 197441
rect 217506 197367 217562 197376
rect 217414 92848 217470 92857
rect 217414 92783 217470 92792
rect 217520 91089 217548 197367
rect 217612 197033 217640 303855
rect 217704 200841 217732 307799
rect 217796 305017 217824 373966
rect 217782 305008 217838 305017
rect 217782 304943 217838 304952
rect 217690 200832 217746 200841
rect 217690 200767 217746 200776
rect 217598 197024 217654 197033
rect 217598 196959 217654 196968
rect 217598 195256 217654 195265
rect 217598 195191 217654 195200
rect 217506 91080 217562 91089
rect 217506 91015 217562 91024
rect 217230 89992 217286 90001
rect 217230 89927 217286 89936
rect 217612 88233 217640 195191
rect 217704 93809 217732 200767
rect 217796 198121 217824 304943
rect 217888 269822 217916 374750
rect 217980 309913 218008 416871
rect 218072 379545 218100 488022
rect 218716 485353 218744 488036
rect 219072 485444 219124 485450
rect 219072 485386 219124 485392
rect 218702 485344 218758 485353
rect 218702 485279 218758 485288
rect 218152 484424 218204 484430
rect 218152 484366 218204 484372
rect 218164 380474 218192 484366
rect 219084 480254 219112 485386
rect 219176 485382 219204 488036
rect 219452 488022 219558 488050
rect 219636 488022 220018 488050
rect 220096 488022 220478 488050
rect 220832 488022 220938 488050
rect 221016 488022 221398 488050
rect 219164 485376 219216 485382
rect 219164 485318 219216 485324
rect 219084 480226 219204 480254
rect 218796 475380 218848 475386
rect 218796 475322 218848 475328
rect 218244 467288 218296 467294
rect 218244 467230 218296 467236
rect 218256 466546 218284 467230
rect 218704 467152 218756 467158
rect 218704 467094 218756 467100
rect 218244 466540 218296 466546
rect 218244 466482 218296 466488
rect 218256 380610 218284 466482
rect 218256 380582 218560 380610
rect 218164 380446 218284 380474
rect 218152 380384 218204 380390
rect 218152 380326 218204 380332
rect 218164 379914 218192 380326
rect 218152 379908 218204 379914
rect 218152 379850 218204 379856
rect 218058 379536 218114 379545
rect 218058 379471 218114 379480
rect 218256 375358 218284 380446
rect 218532 380361 218560 380582
rect 218518 380352 218574 380361
rect 218518 380287 218574 380296
rect 218336 379908 218388 379914
rect 218336 379850 218388 379856
rect 218060 375352 218112 375358
rect 218060 375294 218112 375300
rect 218244 375352 218296 375358
rect 218244 375294 218296 375300
rect 218072 375086 218100 375294
rect 218060 375080 218112 375086
rect 218060 375022 218112 375028
rect 217966 309904 218022 309913
rect 217966 309839 218022 309848
rect 217876 269816 217928 269822
rect 217876 269758 217928 269764
rect 217968 269476 218020 269482
rect 217968 269418 218020 269424
rect 217782 198112 217838 198121
rect 217782 198047 217838 198056
rect 217796 197441 217824 198047
rect 217782 197432 217838 197441
rect 217782 197367 217838 197376
rect 217874 162752 217930 162761
rect 217874 162687 217876 162696
rect 217928 162687 217930 162696
rect 217876 162658 217928 162664
rect 217876 145988 217928 145994
rect 217876 145930 217928 145936
rect 217888 145178 217916 145930
rect 217980 145790 218008 269418
rect 218348 268258 218376 379850
rect 218520 358760 218572 358766
rect 218520 358702 218572 358708
rect 218426 273320 218482 273329
rect 218426 273255 218482 273264
rect 218336 268252 218388 268258
rect 218336 268194 218388 268200
rect 217968 145784 218020 145790
rect 217968 145726 218020 145732
rect 217876 145172 217928 145178
rect 217876 145114 217928 145120
rect 217690 93800 217746 93809
rect 217690 93735 217746 93744
rect 217598 88224 217654 88233
rect 217598 88159 217654 88168
rect 217140 59560 217192 59566
rect 217140 59502 217192 59508
rect 217048 54800 217100 54806
rect 217048 54742 217100 54748
rect 217888 54738 217916 145114
rect 217980 144974 218008 145726
rect 217968 144968 218020 144974
rect 217968 144910 218020 144916
rect 217966 68368 218022 68377
rect 217966 68303 218022 68312
rect 217980 59362 218008 68303
rect 218336 61124 218388 61130
rect 218336 61066 218388 61072
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218348 56098 218376 61066
rect 218440 57390 218468 273255
rect 218532 269278 218560 358702
rect 218612 269816 218664 269822
rect 218612 269758 218664 269764
rect 218520 269272 218572 269278
rect 218520 269214 218572 269220
rect 218520 268660 218572 268666
rect 218520 268602 218572 268608
rect 218532 162654 218560 268602
rect 218520 162648 218572 162654
rect 218520 162590 218572 162596
rect 218624 162178 218652 269758
rect 218612 162172 218664 162178
rect 218612 162114 218664 162120
rect 218520 145512 218572 145518
rect 218520 145454 218572 145460
rect 218532 59702 218560 145454
rect 218612 145104 218664 145110
rect 218612 145046 218664 145052
rect 218624 61130 218652 145046
rect 218612 61124 218664 61130
rect 218612 61066 218664 61072
rect 218716 61010 218744 467094
rect 218808 165170 218836 475322
rect 219072 469940 219124 469946
rect 219072 469882 219124 469888
rect 218888 465860 218940 465866
rect 218888 465802 218940 465808
rect 218796 165164 218848 165170
rect 218796 165106 218848 165112
rect 218900 164898 218928 465802
rect 218978 465760 219034 465769
rect 218978 465695 219034 465704
rect 218992 165306 219020 465695
rect 219084 271386 219112 469882
rect 219176 378894 219204 480226
rect 219256 411460 219308 411466
rect 219256 411402 219308 411408
rect 219164 378888 219216 378894
rect 219164 378830 219216 378836
rect 219176 378622 219204 378830
rect 219164 378616 219216 378622
rect 219164 378558 219216 378564
rect 219268 376174 219296 411402
rect 219452 379438 219480 488022
rect 219636 484242 219664 488022
rect 220096 485874 220124 488022
rect 219544 484214 219664 484242
rect 219820 485846 220124 485874
rect 219440 379432 219492 379438
rect 219440 379374 219492 379380
rect 219440 379160 219492 379166
rect 219440 379102 219492 379108
rect 219256 376168 219308 376174
rect 219256 376110 219308 376116
rect 219348 375352 219400 375358
rect 219348 375294 219400 375300
rect 219256 358692 219308 358698
rect 219256 358634 219308 358640
rect 219164 358284 219216 358290
rect 219164 358226 219216 358232
rect 219072 271380 219124 271386
rect 219072 271322 219124 271328
rect 219176 270366 219204 358226
rect 219164 270360 219216 270366
rect 219164 270302 219216 270308
rect 219072 270088 219124 270094
rect 219072 270030 219124 270036
rect 218980 165300 219032 165306
rect 218980 165242 219032 165248
rect 218888 164892 218940 164898
rect 218888 164834 218940 164840
rect 218888 163532 218940 163538
rect 218888 163474 218940 163480
rect 218796 144764 218848 144770
rect 218796 144706 218848 144712
rect 218624 60982 218744 61010
rect 218520 59696 218572 59702
rect 218520 59638 218572 59644
rect 218428 57384 218480 57390
rect 218428 57326 218480 57332
rect 218624 57254 218652 60982
rect 218702 60616 218758 60625
rect 218702 60551 218758 60560
rect 218716 57730 218744 60551
rect 218704 57724 218756 57730
rect 218704 57666 218756 57672
rect 218612 57248 218664 57254
rect 218612 57190 218664 57196
rect 218336 56092 218388 56098
rect 218336 56034 218388 56040
rect 217876 54732 217928 54738
rect 217876 54674 217928 54680
rect 216404 54664 216456 54670
rect 216404 54606 216456 54612
rect 218808 54534 218836 144706
rect 218900 59498 218928 163474
rect 218980 162648 219032 162654
rect 218980 162590 219032 162596
rect 218888 59492 218940 59498
rect 218888 59434 218940 59440
rect 218992 59294 219020 162590
rect 219084 146062 219112 270030
rect 219176 151814 219204 270302
rect 219268 270026 219296 358634
rect 219360 273630 219388 375294
rect 219348 273624 219400 273630
rect 219348 273566 219400 273572
rect 219452 270494 219480 379102
rect 219544 378962 219572 484214
rect 219820 470594 219848 485846
rect 219900 485784 219952 485790
rect 219900 485726 219952 485732
rect 219636 470566 219848 470594
rect 219636 402974 219664 470566
rect 219636 402946 219848 402974
rect 219716 379636 219768 379642
rect 219716 379578 219768 379584
rect 219624 379296 219676 379302
rect 219624 379238 219676 379244
rect 219532 378956 219584 378962
rect 219532 378898 219584 378904
rect 219360 270466 219480 270494
rect 219360 270230 219388 270466
rect 219348 270224 219400 270230
rect 219348 270166 219400 270172
rect 219256 270020 219308 270026
rect 219256 269962 219308 269968
rect 219268 269346 219296 269962
rect 219256 269340 219308 269346
rect 219256 269282 219308 269288
rect 219176 151786 219296 151814
rect 219268 146198 219296 151786
rect 219256 146192 219308 146198
rect 219256 146134 219308 146140
rect 219072 146056 219124 146062
rect 219072 145998 219124 146004
rect 219084 145586 219112 145998
rect 219072 145580 219124 145586
rect 219072 145522 219124 145528
rect 219072 145444 219124 145450
rect 219072 145386 219124 145392
rect 218980 59288 219032 59294
rect 218980 59230 219032 59236
rect 219084 56506 219112 145386
rect 219268 145110 219296 146134
rect 219360 145926 219388 270166
rect 219636 270162 219664 379238
rect 219624 270156 219676 270162
rect 219624 270098 219676 270104
rect 219624 269272 219676 269278
rect 219624 269214 219676 269220
rect 219636 164150 219664 269214
rect 219728 269074 219756 379578
rect 219820 378758 219848 402946
rect 219808 378752 219860 378758
rect 219808 378694 219860 378700
rect 219912 378604 219940 485726
rect 220176 484424 220228 484430
rect 220176 484366 220228 484372
rect 220188 470594 220216 484366
rect 220832 480282 220860 488022
rect 221016 484242 221044 488022
rect 221752 485314 221780 488036
rect 222242 488022 222608 488050
rect 221740 485308 221792 485314
rect 221740 485250 221792 485256
rect 220924 484214 221044 484242
rect 220820 480276 220872 480282
rect 220820 480218 220872 480224
rect 219820 378576 219940 378604
rect 220004 470566 220216 470594
rect 219820 378214 219848 378576
rect 219808 378208 219860 378214
rect 219808 378150 219860 378156
rect 219820 270502 219848 378150
rect 219900 273624 219952 273630
rect 219900 273566 219952 273572
rect 219808 270496 219860 270502
rect 219808 270438 219860 270444
rect 219808 269340 219860 269346
rect 219808 269282 219860 269288
rect 219716 269068 219768 269074
rect 219716 269010 219768 269016
rect 219624 164144 219676 164150
rect 219624 164086 219676 164092
rect 219532 162172 219584 162178
rect 219532 162114 219584 162120
rect 219348 145920 219400 145926
rect 219348 145862 219400 145868
rect 219360 145722 219388 145862
rect 219348 145716 219400 145722
rect 219348 145658 219400 145664
rect 219440 145716 219492 145722
rect 219440 145658 219492 145664
rect 219348 145580 219400 145586
rect 219348 145522 219400 145528
rect 219256 145104 219308 145110
rect 219256 145046 219308 145052
rect 219256 144968 219308 144974
rect 219162 144936 219218 144945
rect 219256 144910 219308 144916
rect 219162 144871 219218 144880
rect 219072 56500 219124 56506
rect 219072 56442 219124 56448
rect 219176 56234 219204 144871
rect 219268 74534 219296 144910
rect 219360 144770 219388 145522
rect 219452 145382 219480 145658
rect 219440 145376 219492 145382
rect 219440 145318 219492 145324
rect 219348 144764 219400 144770
rect 219348 144706 219400 144712
rect 219268 74506 219388 74534
rect 219254 60616 219310 60625
rect 219254 60551 219310 60560
rect 219268 58682 219296 60551
rect 219256 58676 219308 58682
rect 219256 58618 219308 58624
rect 219164 56228 219216 56234
rect 219164 56170 219216 56176
rect 219360 56166 219388 74506
rect 219348 56160 219400 56166
rect 219348 56102 219400 56108
rect 219544 55010 219572 162114
rect 219532 55004 219584 55010
rect 219532 54946 219584 54952
rect 219636 54942 219664 164086
rect 219728 145382 219756 269010
rect 219716 145376 219768 145382
rect 219716 145318 219768 145324
rect 219624 54936 219676 54942
rect 219624 54878 219676 54884
rect 219728 54874 219756 145318
rect 219820 145314 219848 269282
rect 219912 146305 219940 273566
rect 219898 146296 219954 146305
rect 219898 146231 219954 146240
rect 219808 145308 219860 145314
rect 219808 145250 219860 145256
rect 219820 144974 219848 145250
rect 219808 144968 219860 144974
rect 219912 144945 219940 146231
rect 219808 144910 219860 144916
rect 219898 144936 219954 144945
rect 219898 144871 219954 144880
rect 219900 143336 219952 143342
rect 219900 143278 219952 143284
rect 219912 56302 219940 143278
rect 219900 56296 219952 56302
rect 219900 56238 219952 56244
rect 220004 55826 220032 470566
rect 220924 465798 220952 484214
rect 222580 482361 222608 488022
rect 222672 484430 222700 488036
rect 223162 488022 223528 488050
rect 223500 485081 223528 488022
rect 223486 485072 223542 485081
rect 223486 485007 223542 485016
rect 222660 484424 222712 484430
rect 222660 484366 222712 484372
rect 222566 482352 222622 482361
rect 222566 482287 222622 482296
rect 221004 480276 221056 480282
rect 221004 480218 221056 480224
rect 220912 465792 220964 465798
rect 220912 465734 220964 465740
rect 221016 465730 221044 480218
rect 223592 478281 223620 488036
rect 223990 488022 224264 488050
rect 224450 488022 224816 488050
rect 224236 485246 224264 488022
rect 224224 485240 224276 485246
rect 224224 485182 224276 485188
rect 224788 483750 224816 488022
rect 224880 484537 224908 488036
rect 225370 488022 225644 488050
rect 225738 488022 226104 488050
rect 225616 485110 225644 488022
rect 226076 485314 226104 488022
rect 226064 485308 226116 485314
rect 226064 485250 226116 485256
rect 226168 485217 226196 488036
rect 226536 488022 226642 488050
rect 226720 488022 227102 488050
rect 227272 488022 227562 488050
rect 227732 488022 227930 488050
rect 228008 488022 228390 488050
rect 228560 488022 228850 488050
rect 229326 488022 229600 488050
rect 226154 485208 226210 485217
rect 226154 485143 226210 485152
rect 225604 485104 225656 485110
rect 225604 485046 225656 485052
rect 224866 484528 224922 484537
rect 224866 484463 224922 484472
rect 226340 484152 226392 484158
rect 226340 484094 226392 484100
rect 224776 483744 224828 483750
rect 224776 483686 224828 483692
rect 223578 478272 223634 478281
rect 223578 478207 223634 478216
rect 226352 472666 226380 484094
rect 226432 484016 226484 484022
rect 226432 483958 226484 483964
rect 226444 472870 226472 483958
rect 226536 475561 226564 488022
rect 226720 484158 226748 488022
rect 226708 484152 226760 484158
rect 226708 484094 226760 484100
rect 227272 484022 227300 488022
rect 227260 484016 227312 484022
rect 227260 483958 227312 483964
rect 226522 475552 226578 475561
rect 226522 475487 226578 475496
rect 226432 472864 226484 472870
rect 226432 472806 226484 472812
rect 227732 472734 227760 488022
rect 227812 484152 227864 484158
rect 227812 484094 227864 484100
rect 227824 474026 227852 484094
rect 228008 476921 228036 488022
rect 228560 484158 228588 488022
rect 228548 484152 228600 484158
rect 228548 484094 228600 484100
rect 229572 481030 229600 488022
rect 229756 483818 229784 488036
rect 229848 488022 230138 488050
rect 230614 488022 230704 488050
rect 229744 483812 229796 483818
rect 229744 483754 229796 483760
rect 229560 481024 229612 481030
rect 229560 480966 229612 480972
rect 229848 479641 229876 488022
rect 230676 485178 230704 488022
rect 230768 488022 231058 488050
rect 231534 488022 231808 488050
rect 231902 488022 231992 488050
rect 230664 485172 230716 485178
rect 230664 485114 230716 485120
rect 229834 479632 229890 479641
rect 229834 479567 229890 479576
rect 227994 476912 228050 476921
rect 227994 476847 228050 476856
rect 230768 476785 230796 488022
rect 231780 485353 231808 488022
rect 231766 485344 231822 485353
rect 231766 485279 231822 485288
rect 231860 484152 231912 484158
rect 231860 484094 231912 484100
rect 230754 476776 230810 476785
rect 230754 476711 230810 476720
rect 231872 474094 231900 484094
rect 231964 475833 231992 488022
rect 232332 485489 232360 488036
rect 232424 488022 232806 488050
rect 233282 488022 233648 488050
rect 233742 488022 234016 488050
rect 234110 488022 234384 488050
rect 232318 485480 232374 485489
rect 232318 485415 232374 485424
rect 232424 484158 232452 488022
rect 233620 485761 233648 488022
rect 233606 485752 233662 485761
rect 233606 485687 233662 485696
rect 232412 484152 232464 484158
rect 232412 484094 232464 484100
rect 233988 480865 234016 488022
rect 234356 485217 234384 488022
rect 234540 485382 234568 488036
rect 234632 488022 235014 488050
rect 235490 488022 235856 488050
rect 234528 485376 234580 485382
rect 234528 485318 234580 485324
rect 234342 485208 234398 485217
rect 234342 485143 234398 485152
rect 233974 480856 234030 480865
rect 233974 480791 234030 480800
rect 234632 478417 234660 488022
rect 235828 485625 235856 488022
rect 235814 485616 235870 485625
rect 235814 485551 235870 485560
rect 235920 484945 235948 488036
rect 236318 488022 236408 488050
rect 235906 484936 235962 484945
rect 235906 484871 235962 484880
rect 236000 484152 236052 484158
rect 236000 484094 236052 484100
rect 234618 478408 234674 478417
rect 234618 478343 234674 478352
rect 231950 475824 232006 475833
rect 231950 475759 232006 475768
rect 231860 474088 231912 474094
rect 231860 474030 231912 474036
rect 227812 474020 227864 474026
rect 227812 473962 227864 473968
rect 227720 472728 227772 472734
rect 227720 472670 227772 472676
rect 226340 472660 226392 472666
rect 226340 472602 226392 472608
rect 236012 465798 236040 484094
rect 236380 482497 236408 488022
rect 236472 488022 236762 488050
rect 236840 488022 237222 488050
rect 237392 488022 237682 488050
rect 237760 488022 238142 488050
rect 238220 488022 238510 488050
rect 238772 488022 238970 488050
rect 239446 488022 239720 488050
rect 239906 488022 240088 488050
rect 236366 482488 236422 482497
rect 236366 482423 236422 482432
rect 236472 479534 236500 488022
rect 236840 484158 236868 488022
rect 236828 484152 236880 484158
rect 236828 484094 236880 484100
rect 236460 479528 236512 479534
rect 236460 479470 236512 479476
rect 237392 472802 237420 488022
rect 237760 484106 237788 488022
rect 237484 484078 237788 484106
rect 237484 476814 237512 484078
rect 238220 478174 238248 488022
rect 238208 478168 238260 478174
rect 238208 478110 238260 478116
rect 238772 476882 238800 488022
rect 239692 485518 239720 488022
rect 239680 485512 239732 485518
rect 239680 485454 239732 485460
rect 240060 485450 240088 488022
rect 240152 488022 240258 488050
rect 240336 488022 240718 488050
rect 240888 488022 241178 488050
rect 240048 485444 240100 485450
rect 240048 485386 240100 485392
rect 238760 476876 238812 476882
rect 238760 476818 238812 476824
rect 237472 476808 237524 476814
rect 237472 476750 237524 476756
rect 240152 473074 240180 488022
rect 240232 484152 240284 484158
rect 240232 484094 240284 484100
rect 240140 473068 240192 473074
rect 240140 473010 240192 473016
rect 240244 472938 240272 484094
rect 240336 475697 240364 488022
rect 240888 484158 240916 488022
rect 240876 484152 240928 484158
rect 240876 484094 240928 484100
rect 241520 484152 241572 484158
rect 241520 484094 241572 484100
rect 240322 475688 240378 475697
rect 240322 475623 240378 475632
rect 240232 472932 240284 472938
rect 240232 472874 240284 472880
rect 237380 472796 237432 472802
rect 237380 472738 237432 472744
rect 241532 465866 241560 484094
rect 241624 473006 241652 488036
rect 241716 488022 242098 488050
rect 242176 488022 242466 488050
rect 241716 476950 241744 488022
rect 242176 484158 242204 488022
rect 242928 487778 242956 488036
rect 243188 488022 243386 488050
rect 243464 488022 243846 488050
rect 244322 488022 244596 488050
rect 244690 488022 245056 488050
rect 245150 488022 245240 488050
rect 242928 487750 243124 487778
rect 242164 484152 242216 484158
rect 242164 484094 242216 484100
rect 243096 481098 243124 487750
rect 243084 481092 243136 481098
rect 243084 481034 243136 481040
rect 243188 480978 243216 488022
rect 242912 480950 243216 480978
rect 241704 476944 241756 476950
rect 241704 476886 241756 476892
rect 241612 473000 241664 473006
rect 241612 472942 241664 472948
rect 241520 465860 241572 465866
rect 241520 465802 241572 465808
rect 236000 465792 236052 465798
rect 236000 465734 236052 465740
rect 242912 465730 242940 480950
rect 243464 474230 243492 488022
rect 244568 485586 244596 488022
rect 244556 485580 244608 485586
rect 244556 485522 244608 485528
rect 245028 482322 245056 488022
rect 245212 483954 245240 488022
rect 245304 488022 245594 488050
rect 245948 488022 246054 488050
rect 246132 488022 246422 488050
rect 246592 488022 246882 488050
rect 245200 483948 245252 483954
rect 245200 483890 245252 483896
rect 245016 482316 245068 482322
rect 245016 482258 245068 482264
rect 243452 474224 243504 474230
rect 243452 474166 243504 474172
rect 245304 470594 245332 488022
rect 245660 480888 245712 480894
rect 245660 480830 245712 480836
rect 245672 474366 245700 480830
rect 245948 479602 245976 488022
rect 245936 479596 245988 479602
rect 245936 479538 245988 479544
rect 246132 476114 246160 488022
rect 246592 480894 246620 488022
rect 247328 481001 247356 488036
rect 247420 488022 247802 488050
rect 248278 488022 248368 488050
rect 248646 488022 248736 488050
rect 247314 480992 247370 481001
rect 247314 480927 247370 480936
rect 246580 480888 246632 480894
rect 246580 480830 246632 480836
rect 247420 478242 247448 488022
rect 248340 483886 248368 488022
rect 248512 487076 248564 487082
rect 248512 487018 248564 487024
rect 248328 483880 248380 483886
rect 248328 483822 248380 483828
rect 248420 480888 248472 480894
rect 248420 480830 248472 480836
rect 247408 478236 247460 478242
rect 247408 478178 247460 478184
rect 245764 476086 246160 476114
rect 245764 475386 245792 476086
rect 245752 475380 245804 475386
rect 245752 475322 245804 475328
rect 245660 474360 245712 474366
rect 245660 474302 245712 474308
rect 244292 470566 245332 470594
rect 244292 465934 244320 470566
rect 248432 466002 248460 480830
rect 248524 466070 248552 487018
rect 248708 485774 248736 488022
rect 248800 488022 249090 488050
rect 249168 488022 249550 488050
rect 249812 488022 250010 488050
rect 250088 488022 250470 488050
rect 250548 488022 250838 488050
rect 248800 487082 248828 488022
rect 248788 487076 248840 487082
rect 248788 487018 248840 487024
rect 248708 485746 248828 485774
rect 248800 476114 248828 485746
rect 249168 480894 249196 488022
rect 249156 480888 249208 480894
rect 249156 480830 249208 480836
rect 248616 476086 248828 476114
rect 248616 466138 248644 476086
rect 249812 468654 249840 488022
rect 250088 476114 250116 488022
rect 249904 476086 250116 476114
rect 249800 468648 249852 468654
rect 249800 468590 249852 468596
rect 249904 468586 249932 476086
rect 250548 471306 250576 488022
rect 251180 481160 251232 481166
rect 251180 481102 251232 481108
rect 250536 471300 250588 471306
rect 250536 471242 250588 471248
rect 249892 468580 249944 468586
rect 249892 468522 249944 468528
rect 251192 467294 251220 481102
rect 251284 480978 251312 488036
rect 251376 488022 251758 488050
rect 251928 488022 252218 488050
rect 251376 481166 251404 488022
rect 251364 481160 251416 481166
rect 251364 481102 251416 481108
rect 251284 480950 251404 480978
rect 251272 480888 251324 480894
rect 251272 480830 251324 480836
rect 251180 467288 251232 467294
rect 251180 467230 251232 467236
rect 251284 467226 251312 480830
rect 251376 474434 251404 480950
rect 251928 480894 251956 488022
rect 251916 480888 251968 480894
rect 251916 480830 251968 480836
rect 251364 474428 251416 474434
rect 251364 474370 251416 474376
rect 251272 467220 251324 467226
rect 251272 467162 251324 467168
rect 252572 467158 252600 488036
rect 252756 488022 253046 488050
rect 253216 488022 253506 488050
rect 253982 488022 254072 488050
rect 252652 480888 252704 480894
rect 252652 480830 252704 480836
rect 252664 468518 252692 480830
rect 252756 474298 252784 488022
rect 253216 480894 253244 488022
rect 253204 480888 253256 480894
rect 253204 480830 253256 480836
rect 253940 480888 253992 480894
rect 253940 480830 253992 480836
rect 252744 474292 252796 474298
rect 252744 474234 252796 474240
rect 252652 468512 252704 468518
rect 252652 468454 252704 468460
rect 253952 467498 253980 480830
rect 254044 474162 254072 488022
rect 254136 488022 254426 488050
rect 254504 488022 254794 488050
rect 254872 488022 255254 488050
rect 255332 488022 255714 488050
rect 255792 488022 256174 488050
rect 256344 488022 256634 488050
rect 256712 488022 257002 488050
rect 257478 488022 257752 488050
rect 257938 488022 258028 488050
rect 254136 475969 254164 488022
rect 254504 480894 254532 488022
rect 254492 480888 254544 480894
rect 254492 480830 254544 480836
rect 254872 477086 254900 488022
rect 254860 477080 254912 477086
rect 254860 477022 254912 477028
rect 254122 475960 254178 475969
rect 254122 475895 254178 475904
rect 254032 474156 254084 474162
rect 254032 474098 254084 474104
rect 255332 468858 255360 488022
rect 255792 479806 255820 488022
rect 255780 479800 255832 479806
rect 256344 479777 256372 488022
rect 255780 479742 255832 479748
rect 256330 479768 256386 479777
rect 256712 479738 256740 488022
rect 257724 482458 257752 488022
rect 258000 484090 258028 488022
rect 258092 488022 258382 488050
rect 258460 488022 258842 488050
rect 258920 488022 259210 488050
rect 259564 488022 259670 488050
rect 259748 488022 260130 488050
rect 260208 488022 260590 488050
rect 260974 488022 261248 488050
rect 261434 488022 261800 488050
rect 261894 488022 262168 488050
rect 257988 484084 258040 484090
rect 257988 484026 258040 484032
rect 257712 482452 257764 482458
rect 257712 482394 257764 482400
rect 256330 479703 256386 479712
rect 256700 479732 256752 479738
rect 256700 479674 256752 479680
rect 255320 468852 255372 468858
rect 255320 468794 255372 468800
rect 253940 467492 253992 467498
rect 253940 467434 253992 467440
rect 258092 467362 258120 488022
rect 258460 479670 258488 488022
rect 258448 479664 258500 479670
rect 258448 479606 258500 479612
rect 258920 477154 258948 488022
rect 259564 485774 259592 488022
rect 259748 485774 259776 488022
rect 259472 485746 259592 485774
rect 259656 485746 259776 485774
rect 259472 480894 259500 485746
rect 259656 481114 259684 485746
rect 259564 481086 259684 481114
rect 259460 480888 259512 480894
rect 259460 480830 259512 480836
rect 259460 479460 259512 479466
rect 259460 479402 259512 479408
rect 258908 477148 258960 477154
rect 258908 477090 258960 477096
rect 258080 467356 258132 467362
rect 258080 467298 258132 467304
rect 252560 467152 252612 467158
rect 252560 467094 252612 467100
rect 259472 466274 259500 479402
rect 259564 471374 259592 481086
rect 259644 480888 259696 480894
rect 259644 480830 259696 480836
rect 259656 475454 259684 480830
rect 260208 479466 260236 488022
rect 261220 481166 261248 488022
rect 261772 482390 261800 488022
rect 262140 484022 262168 488022
rect 262128 484016 262180 484022
rect 262128 483958 262180 483964
rect 261760 482384 261812 482390
rect 261760 482326 261812 482332
rect 261208 481160 261260 481166
rect 261208 481102 261260 481108
rect 262220 480888 262272 480894
rect 262220 480830 262272 480836
rect 260196 479460 260248 479466
rect 260196 479402 260248 479408
rect 259644 475448 259696 475454
rect 259644 475390 259696 475396
rect 259552 471368 259604 471374
rect 259552 471310 259604 471316
rect 259460 466268 259512 466274
rect 259460 466210 259512 466216
rect 262232 466206 262260 480830
rect 262324 467430 262352 488036
rect 262416 488022 262798 488050
rect 262876 488022 263166 488050
rect 262416 480894 262444 488022
rect 262404 480888 262456 480894
rect 262404 480830 262456 480836
rect 262876 473142 262904 488022
rect 263612 474570 263640 488036
rect 263796 488022 264086 488050
rect 264256 488022 264546 488050
rect 263692 484152 263744 484158
rect 263692 484094 263744 484100
rect 263704 477222 263732 484094
rect 263692 477216 263744 477222
rect 263692 477158 263744 477164
rect 263796 477018 263824 488022
rect 264256 484158 264284 488022
rect 264244 484152 264296 484158
rect 264244 484094 264296 484100
rect 263784 477012 263836 477018
rect 263784 476954 263836 476960
rect 263600 474564 263652 474570
rect 263600 474506 263652 474512
rect 262864 473136 262916 473142
rect 262864 473078 262916 473084
rect 262312 467424 262364 467430
rect 262312 467366 262364 467372
rect 262220 466200 262272 466206
rect 262220 466142 262272 466148
rect 248604 466132 248656 466138
rect 248604 466074 248656 466080
rect 248512 466064 248564 466070
rect 248512 466006 248564 466012
rect 248420 465996 248472 466002
rect 248420 465938 248472 465944
rect 244280 465928 244332 465934
rect 244280 465870 244332 465876
rect 221004 465724 221056 465730
rect 221004 465666 221056 465672
rect 242900 465724 242952 465730
rect 242900 465666 242952 465672
rect 264992 464370 265020 488036
rect 265176 488022 265374 488050
rect 265452 488022 265834 488050
rect 265912 488022 266294 488050
rect 266464 488022 266754 488050
rect 266832 488022 267122 488050
rect 267200 488022 267582 488050
rect 267844 488022 268042 488050
rect 268120 488022 268502 488050
rect 268672 488022 268962 488050
rect 269132 488022 269330 488050
rect 269408 488022 269790 488050
rect 269960 488022 270250 488050
rect 270604 488022 270710 488050
rect 270880 488022 271170 488050
rect 271248 488022 271538 488050
rect 271892 488022 271998 488050
rect 272076 488022 272458 488050
rect 272536 488022 272918 488050
rect 273302 488022 273392 488050
rect 265072 484152 265124 484158
rect 265072 484094 265124 484100
rect 265084 468489 265112 484094
rect 265176 468790 265204 488022
rect 265452 470594 265480 488022
rect 265912 484158 265940 488022
rect 265900 484152 265952 484158
rect 265900 484094 265952 484100
rect 266360 484152 266412 484158
rect 266360 484094 266412 484100
rect 265268 470566 265480 470594
rect 265268 469878 265296 470566
rect 265256 469872 265308 469878
rect 265256 469814 265308 469820
rect 266372 468994 266400 484094
rect 266360 468988 266412 468994
rect 266360 468930 266412 468936
rect 266464 468926 266492 488022
rect 266832 484158 266860 488022
rect 266820 484152 266872 484158
rect 266820 484094 266872 484100
rect 267200 470594 267228 488022
rect 267740 484152 267792 484158
rect 267740 484094 267792 484100
rect 266556 470566 267228 470594
rect 266452 468920 266504 468926
rect 266452 468862 266504 468868
rect 265164 468784 265216 468790
rect 265164 468726 265216 468732
rect 266556 468722 266584 470566
rect 266544 468716 266596 468722
rect 266544 468658 266596 468664
rect 265070 468480 265126 468489
rect 265070 468415 265126 468424
rect 267752 466342 267780 484094
rect 267844 470150 267872 488022
rect 268120 474502 268148 488022
rect 268672 484158 268700 488022
rect 268660 484152 268712 484158
rect 268660 484094 268712 484100
rect 268108 474496 268160 474502
rect 268108 474438 268160 474444
rect 267832 470144 267884 470150
rect 267832 470086 267884 470092
rect 269132 469130 269160 488022
rect 269212 484152 269264 484158
rect 269212 484094 269264 484100
rect 269224 478514 269252 484094
rect 269212 478508 269264 478514
rect 269212 478450 269264 478456
rect 269408 478446 269436 488022
rect 269960 484158 269988 488022
rect 269948 484152 270000 484158
rect 269948 484094 270000 484100
rect 270500 484152 270552 484158
rect 270500 484094 270552 484100
rect 269396 478440 269448 478446
rect 269396 478382 269448 478388
rect 270512 475522 270540 484094
rect 270604 478310 270632 488022
rect 270880 478378 270908 488022
rect 271248 484158 271276 488022
rect 271236 484152 271288 484158
rect 271236 484094 271288 484100
rect 270868 478372 270920 478378
rect 270868 478314 270920 478320
rect 270592 478304 270644 478310
rect 270592 478246 270644 478252
rect 270500 475516 270552 475522
rect 270500 475458 270552 475464
rect 269120 469124 269172 469130
rect 269120 469066 269172 469072
rect 267740 466336 267792 466342
rect 267740 466278 267792 466284
rect 271892 464438 271920 488022
rect 271972 484152 272024 484158
rect 271972 484094 272024 484100
rect 271984 474638 272012 484094
rect 272076 479874 272104 488022
rect 272536 484158 272564 488022
rect 272524 484152 272576 484158
rect 272524 484094 272576 484100
rect 273260 484152 273312 484158
rect 273260 484094 273312 484100
rect 272064 479868 272116 479874
rect 272064 479810 272116 479816
rect 271972 474632 272024 474638
rect 271972 474574 272024 474580
rect 273272 467634 273300 484094
rect 273260 467628 273312 467634
rect 273260 467570 273312 467576
rect 273364 467566 273392 488022
rect 273456 488022 273746 488050
rect 273824 488022 274206 488050
rect 273456 469062 273484 488022
rect 273824 484158 273852 488022
rect 274668 487830 274696 488036
rect 274744 488022 275126 488050
rect 275204 488022 275494 488050
rect 275664 488022 275954 488050
rect 276032 488022 276414 488050
rect 276890 488022 277164 488050
rect 274656 487824 274708 487830
rect 274656 487766 274708 487772
rect 273812 484152 273864 484158
rect 273812 484094 273864 484100
rect 274640 484152 274692 484158
rect 274640 484094 274692 484100
rect 273444 469056 273496 469062
rect 273444 468998 273496 469004
rect 273352 467560 273404 467566
rect 273352 467502 273404 467508
rect 274652 466410 274680 484094
rect 274744 477290 274772 488022
rect 274824 487824 274876 487830
rect 274824 487766 274876 487772
rect 274836 482662 274864 487766
rect 275204 484158 275232 488022
rect 275192 484152 275244 484158
rect 275192 484094 275244 484100
rect 274824 482656 274876 482662
rect 274824 482598 274876 482604
rect 275664 479942 275692 488022
rect 275652 479936 275704 479942
rect 275652 479878 275704 479884
rect 274732 477284 274784 477290
rect 274732 477226 274784 477232
rect 276032 474706 276060 488022
rect 277136 482633 277164 488022
rect 277122 482624 277178 482633
rect 277122 482559 277178 482568
rect 277320 482526 277348 488036
rect 277504 488022 277702 488050
rect 277400 484152 277452 484158
rect 277400 484094 277452 484100
rect 277308 482520 277360 482526
rect 277308 482462 277360 482468
rect 276020 474700 276072 474706
rect 276020 474642 276072 474648
rect 277412 467702 277440 484094
rect 277504 469198 277532 488022
rect 278148 482594 278176 488036
rect 278240 488022 278622 488050
rect 278884 488022 279082 488050
rect 279160 488022 279542 488050
rect 279926 488022 280108 488050
rect 280386 488022 280752 488050
rect 280846 488022 281120 488050
rect 281306 488022 281488 488050
rect 278240 484158 278268 488022
rect 278228 484152 278280 484158
rect 278228 484094 278280 484100
rect 278780 484152 278832 484158
rect 278780 484094 278832 484100
rect 278136 482588 278188 482594
rect 278136 482530 278188 482536
rect 278792 477358 278820 484094
rect 278884 480010 278912 488022
rect 279160 484158 279188 488022
rect 280080 484226 280108 488022
rect 280068 484220 280120 484226
rect 280068 484162 280120 484168
rect 279148 484152 279200 484158
rect 279148 484094 279200 484100
rect 280724 481137 280752 488022
rect 281092 481234 281120 488022
rect 281460 481302 281488 488022
rect 281552 488022 281658 488050
rect 281736 488022 282118 488050
rect 282288 488022 282578 488050
rect 283054 488022 283144 488050
rect 281448 481296 281500 481302
rect 281448 481238 281500 481244
rect 281080 481228 281132 481234
rect 281080 481170 281132 481176
rect 280710 481128 280766 481137
rect 280710 481063 280766 481072
rect 278872 480004 278924 480010
rect 278872 479946 278924 479952
rect 278780 477352 278832 477358
rect 278780 477294 278832 477300
rect 281552 470354 281580 488022
rect 281632 484152 281684 484158
rect 281632 484094 281684 484100
rect 281540 470348 281592 470354
rect 281540 470290 281592 470296
rect 281644 470014 281672 484094
rect 281736 470218 281764 488022
rect 282288 484158 282316 488022
rect 282276 484152 282328 484158
rect 282276 484094 282328 484100
rect 282920 484152 282972 484158
rect 282920 484094 282972 484100
rect 282932 470422 282960 484094
rect 283012 481364 283064 481370
rect 283012 481306 283064 481312
rect 282920 470416 282972 470422
rect 282920 470358 282972 470364
rect 281724 470212 281776 470218
rect 281724 470154 281776 470160
rect 281632 470008 281684 470014
rect 281632 469950 281684 469956
rect 283024 469810 283052 481306
rect 283116 470490 283144 488022
rect 283208 488022 283498 488050
rect 283576 488022 283866 488050
rect 283208 484158 283236 488022
rect 283196 484152 283248 484158
rect 283196 484094 283248 484100
rect 283576 481370 283604 488022
rect 283564 481364 283616 481370
rect 283564 481306 283616 481312
rect 283104 470484 283156 470490
rect 283104 470426 283156 470432
rect 284312 469946 284340 488036
rect 284802 488022 285168 488050
rect 285262 488022 285536 488050
rect 285140 482730 285168 488022
rect 285508 484362 285536 488022
rect 285496 484356 285548 484362
rect 285496 484298 285548 484304
rect 285128 482724 285180 482730
rect 285128 482666 285180 482672
rect 285692 470082 285720 488036
rect 285864 484288 285916 484294
rect 285864 484230 285916 484236
rect 285772 484152 285824 484158
rect 285772 484094 285824 484100
rect 285784 471986 285812 484094
rect 285772 471980 285824 471986
rect 285772 471922 285824 471928
rect 285876 471442 285904 484230
rect 286060 480298 286088 488036
rect 286152 488022 286534 488050
rect 286704 488022 286994 488050
rect 286152 484294 286180 488022
rect 286140 484288 286192 484294
rect 286140 484230 286192 484236
rect 286704 484158 286732 488022
rect 286692 484152 286744 484158
rect 286692 484094 286744 484100
rect 287060 484152 287112 484158
rect 287060 484094 287112 484100
rect 285968 480270 286088 480298
rect 285968 473210 285996 480270
rect 285956 473204 286008 473210
rect 285956 473146 286008 473152
rect 285864 471436 285916 471442
rect 285864 471378 285916 471384
rect 285680 470076 285732 470082
rect 285680 470018 285732 470024
rect 284300 469940 284352 469946
rect 284300 469882 284352 469888
rect 283012 469804 283064 469810
rect 283012 469746 283064 469752
rect 277492 469192 277544 469198
rect 277492 469134 277544 469140
rect 277400 467696 277452 467702
rect 277400 467638 277452 467644
rect 274640 466404 274692 466410
rect 274640 466346 274692 466352
rect 287072 464506 287100 484094
rect 287440 483614 287468 488036
rect 287532 488022 287822 488050
rect 287992 488022 288282 488050
rect 288544 488022 288742 488050
rect 288912 488022 289202 488050
rect 289678 488022 289768 488050
rect 287428 483608 287480 483614
rect 287428 483550 287480 483556
rect 287532 471918 287560 488022
rect 287992 484158 288020 488022
rect 287980 484152 288032 484158
rect 287980 484094 288032 484100
rect 288440 484152 288492 484158
rect 288440 484094 288492 484100
rect 287520 471912 287572 471918
rect 287520 471854 287572 471860
rect 288452 465662 288480 484094
rect 288544 473958 288572 488022
rect 288912 484158 288940 488022
rect 289740 484294 289768 488022
rect 289832 488022 290030 488050
rect 290200 488022 290490 488050
rect 290568 488022 290950 488050
rect 289728 484288 289780 484294
rect 289728 484230 289780 484236
rect 288900 484152 288952 484158
rect 288900 484094 288952 484100
rect 288532 473952 288584 473958
rect 288532 473894 288584 473900
rect 289832 470558 289860 488022
rect 289912 484152 289964 484158
rect 289912 484094 289964 484100
rect 289924 473890 289952 484094
rect 290200 475658 290228 488022
rect 290568 484158 290596 488022
rect 291200 484288 291252 484294
rect 291200 484230 291252 484236
rect 290556 484152 290608 484158
rect 290556 484094 290608 484100
rect 290188 475652 290240 475658
rect 290188 475594 290240 475600
rect 289912 473884 289964 473890
rect 289912 473826 289964 473832
rect 289820 470552 289872 470558
rect 289820 470494 289872 470500
rect 291212 467770 291240 484230
rect 291292 484152 291344 484158
rect 291292 484094 291344 484100
rect 291304 477494 291332 484094
rect 291292 477488 291344 477494
rect 291292 477430 291344 477436
rect 291396 477426 291424 488036
rect 291488 488022 291870 488050
rect 291948 488022 292238 488050
rect 292592 488022 292698 488050
rect 292776 488022 293158 488050
rect 293328 488022 293618 488050
rect 294002 488022 294092 488050
rect 291488 484158 291516 488022
rect 291948 484294 291976 488022
rect 291936 484288 291988 484294
rect 291936 484230 291988 484236
rect 291476 484152 291528 484158
rect 291476 484094 291528 484100
rect 291384 477420 291436 477426
rect 291384 477362 291436 477368
rect 291200 467764 291252 467770
rect 291200 467706 291252 467712
rect 292592 465769 292620 488022
rect 292672 480344 292724 480350
rect 292672 480286 292724 480292
rect 292684 471578 292712 480286
rect 292776 475590 292804 488022
rect 293328 480350 293356 488022
rect 294064 481370 294092 488022
rect 294156 488022 294446 488050
rect 294616 488022 294906 488050
rect 294052 481364 294104 481370
rect 294052 481306 294104 481312
rect 293316 480344 293368 480350
rect 293316 480286 293368 480292
rect 294156 478122 294184 488022
rect 294236 481364 294288 481370
rect 294236 481306 294288 481312
rect 293972 478094 294184 478122
rect 292764 475584 292816 475590
rect 292764 475526 292816 475532
rect 292672 471572 292724 471578
rect 292672 471514 292724 471520
rect 293972 468450 294000 478094
rect 294248 473354 294276 481306
rect 294616 480078 294644 488022
rect 294604 480072 294656 480078
rect 294604 480014 294656 480020
rect 294064 473326 294276 473354
rect 294064 471510 294092 473326
rect 295352 471646 295380 488036
rect 295536 488022 295826 488050
rect 295904 488022 296194 488050
rect 296272 488022 296654 488050
rect 296824 488022 297114 488050
rect 297192 488022 297574 488050
rect 297744 488022 298034 488050
rect 298204 488022 298402 488050
rect 298480 488022 298862 488050
rect 299032 488022 299322 488050
rect 299492 488022 299782 488050
rect 295432 480888 295484 480894
rect 295432 480830 295484 480836
rect 295444 471782 295472 480830
rect 295536 471850 295564 488022
rect 295904 480894 295932 488022
rect 295892 480888 295944 480894
rect 295892 480830 295944 480836
rect 295524 471844 295576 471850
rect 295524 471786 295576 471792
rect 295432 471776 295484 471782
rect 295432 471718 295484 471724
rect 296272 471714 296300 488022
rect 296720 480888 296772 480894
rect 296720 480830 296772 480836
rect 296260 471708 296312 471714
rect 296260 471650 296312 471656
rect 295340 471640 295392 471646
rect 295340 471582 295392 471588
rect 294052 471504 294104 471510
rect 294052 471446 294104 471452
rect 293960 468444 294012 468450
rect 293960 468386 294012 468392
rect 296732 468382 296760 480830
rect 296824 470286 296852 488022
rect 297192 478553 297220 488022
rect 297364 484152 297416 484158
rect 297364 484094 297416 484100
rect 297376 483614 297404 484094
rect 297364 483608 297416 483614
rect 297364 483550 297416 483556
rect 297744 480894 297772 488022
rect 297732 480888 297784 480894
rect 297732 480830 297784 480836
rect 298100 480888 298152 480894
rect 298100 480830 298152 480836
rect 297178 478544 297234 478553
rect 297178 478479 297234 478488
rect 296812 470280 296864 470286
rect 296812 470222 296864 470228
rect 296720 468376 296772 468382
rect 296720 468318 296772 468324
rect 292578 465760 292634 465769
rect 292578 465695 292634 465704
rect 288440 465656 288492 465662
rect 288440 465598 288492 465604
rect 298112 465594 298140 480830
rect 298204 471209 298232 488022
rect 298480 480894 298508 488022
rect 298468 480888 298520 480894
rect 298468 480830 298520 480836
rect 299032 473278 299060 488022
rect 299020 473272 299072 473278
rect 299020 473214 299072 473220
rect 299492 471238 299520 488022
rect 312556 482225 312584 623766
rect 312648 563990 312676 641038
rect 315304 640960 315356 640966
rect 315304 640902 315356 640908
rect 314016 640688 314068 640694
rect 314016 640630 314068 640636
rect 313924 632120 313976 632126
rect 313924 632062 313976 632068
rect 312636 563984 312688 563990
rect 312636 563926 312688 563932
rect 312912 552560 312964 552566
rect 312912 552502 312964 552508
rect 312728 552492 312780 552498
rect 312728 552434 312780 552440
rect 312636 552084 312688 552090
rect 312636 552026 312688 552032
rect 312648 522986 312676 552026
rect 312636 522980 312688 522986
rect 312636 522922 312688 522928
rect 312740 522918 312768 552434
rect 312820 551132 312872 551138
rect 312820 551074 312872 551080
rect 312832 524278 312860 551074
rect 312924 527134 312952 552502
rect 313004 552424 313056 552430
rect 313004 552366 313056 552372
rect 313016 528562 313044 552366
rect 313096 551200 313148 551206
rect 313096 551142 313148 551148
rect 313004 528556 313056 528562
rect 313004 528498 313056 528504
rect 313108 528494 313136 551142
rect 313096 528488 313148 528494
rect 313096 528430 313148 528436
rect 312912 527128 312964 527134
rect 312912 527070 312964 527076
rect 313936 526318 313964 632062
rect 314028 559706 314056 640630
rect 314016 559700 314068 559706
rect 314016 559642 314068 559648
rect 315316 556850 315344 640902
rect 316684 640892 316736 640898
rect 316684 640834 316736 640840
rect 315304 556844 315356 556850
rect 315304 556786 315356 556792
rect 316696 552906 316724 640834
rect 316868 640620 316920 640626
rect 316868 640562 316920 640568
rect 316776 636880 316828 636886
rect 316776 636822 316828 636828
rect 316788 575657 316816 636822
rect 316774 575648 316830 575657
rect 316774 575583 316830 575592
rect 316774 570888 316830 570897
rect 316774 570823 316830 570832
rect 316684 552900 316736 552906
rect 316684 552842 316736 552848
rect 315396 552356 315448 552362
rect 315396 552298 315448 552304
rect 315304 552220 315356 552226
rect 315304 552162 315356 552168
rect 314016 550928 314068 550934
rect 314016 550870 314068 550876
rect 313924 526312 313976 526318
rect 313924 526254 313976 526260
rect 314028 524822 314056 550870
rect 314016 524816 314068 524822
rect 314016 524758 314068 524764
rect 312820 524272 312872 524278
rect 312820 524214 312872 524220
rect 312728 522912 312780 522918
rect 312728 522854 312780 522860
rect 315316 522850 315344 552162
rect 315408 526590 315436 552298
rect 316684 550792 316736 550798
rect 316684 550734 316736 550740
rect 315488 549568 315540 549574
rect 315488 549510 315540 549516
rect 315500 526930 315528 549510
rect 315672 548820 315724 548826
rect 315672 548762 315724 548768
rect 315578 548040 315634 548049
rect 315578 547975 315634 547984
rect 315592 527066 315620 547975
rect 315684 528426 315712 548762
rect 315672 528420 315724 528426
rect 315672 528362 315724 528368
rect 315580 527060 315632 527066
rect 315580 527002 315632 527008
rect 315488 526924 315540 526930
rect 315488 526866 315540 526872
rect 315396 526584 315448 526590
rect 315396 526526 315448 526532
rect 316696 525434 316724 550734
rect 316684 525428 316736 525434
rect 316684 525370 316736 525376
rect 315304 522844 315356 522850
rect 315304 522786 315356 522792
rect 316788 483682 316816 570823
rect 316880 554130 316908 640562
rect 316960 640484 317012 640490
rect 316960 640426 317012 640432
rect 316972 565350 317000 640426
rect 317064 568002 317092 643146
rect 318800 642388 318852 642394
rect 318800 642330 318852 642336
rect 318246 640520 318302 640529
rect 318246 640455 318302 640464
rect 318156 640416 318208 640422
rect 318156 640358 318208 640364
rect 317970 638208 318026 638217
rect 317970 638143 318026 638152
rect 317984 637702 318012 638143
rect 317972 637696 318024 637702
rect 317972 637638 318024 637644
rect 318062 633448 318118 633457
rect 318062 633383 318118 633392
rect 317694 628688 317750 628697
rect 317694 628623 317750 628632
rect 317708 627978 317736 628623
rect 317696 627972 317748 627978
rect 317696 627914 317748 627920
rect 317418 623928 317474 623937
rect 317418 623863 317474 623872
rect 317432 623830 317460 623863
rect 317420 623824 317472 623830
rect 317420 623766 317472 623772
rect 317602 619168 317658 619177
rect 317602 619103 317658 619112
rect 317616 618322 317644 619103
rect 317604 618316 317656 618322
rect 317604 618258 317656 618264
rect 317970 614408 318026 614417
rect 317970 614343 318026 614352
rect 317984 614174 318012 614343
rect 317972 614168 318024 614174
rect 317972 614110 318024 614116
rect 317970 609648 318026 609657
rect 317970 609583 318026 609592
rect 317984 608666 318012 609583
rect 317972 608660 318024 608666
rect 317972 608602 318024 608608
rect 317970 604888 318026 604897
rect 317970 604823 318026 604832
rect 317984 604518 318012 604823
rect 317972 604512 318024 604518
rect 317972 604454 318024 604460
rect 317970 595368 318026 595377
rect 317970 595303 318026 595312
rect 317984 594862 318012 595303
rect 317972 594856 318024 594862
rect 317972 594798 318024 594804
rect 317970 590608 318026 590617
rect 317970 590543 318026 590552
rect 317984 589354 318012 590543
rect 317972 589348 318024 589354
rect 317972 589290 318024 589296
rect 317970 585848 318026 585857
rect 317970 585783 318026 585792
rect 317984 585206 318012 585783
rect 317972 585200 318024 585206
rect 317972 585142 318024 585148
rect 317970 580408 318026 580417
rect 317970 580343 318026 580352
rect 317984 579698 318012 580343
rect 317972 579692 318024 579698
rect 317972 579634 318024 579640
rect 317052 567996 317104 568002
rect 317052 567938 317104 567944
rect 317970 566128 318026 566137
rect 317970 566063 318026 566072
rect 317984 565894 318012 566063
rect 317972 565888 318024 565894
rect 317972 565830 318024 565836
rect 316960 565344 317012 565350
rect 316960 565286 317012 565292
rect 317970 561368 318026 561377
rect 317970 561303 318026 561312
rect 317984 560318 318012 561303
rect 317972 560312 318024 560318
rect 317972 560254 318024 560260
rect 318076 557534 318104 633383
rect 318168 559774 318196 640358
rect 318260 563854 318288 640455
rect 318340 639396 318392 639402
rect 318340 639338 318392 639344
rect 318352 596834 318380 639338
rect 318812 600137 318840 642330
rect 378600 641232 378652 641238
rect 378600 641174 378652 641180
rect 332876 641164 332928 641170
rect 332876 641106 332928 641112
rect 319628 641028 319680 641034
rect 319628 640970 319680 640976
rect 319536 640348 319588 640354
rect 319536 640290 319588 640296
rect 319444 639328 319496 639334
rect 319444 639270 319496 639276
rect 318798 600128 318854 600137
rect 318798 600063 318854 600072
rect 318340 596828 318392 596834
rect 318340 596770 318392 596776
rect 318248 563848 318300 563854
rect 318248 563790 318300 563796
rect 318156 559768 318208 559774
rect 318156 559710 318208 559716
rect 317420 557524 317472 557530
rect 317420 557466 317472 557472
rect 317984 557506 318104 557534
rect 317432 556617 317460 557466
rect 317418 556608 317474 556617
rect 317418 556543 317474 556552
rect 316868 554124 316920 554130
rect 316868 554066 316920 554072
rect 316868 552288 316920 552294
rect 316868 552230 316920 552236
rect 316880 522782 316908 552230
rect 317984 551410 318012 557506
rect 318524 552628 318576 552634
rect 318524 552570 318576 552576
rect 318432 552152 318484 552158
rect 318432 552094 318484 552100
rect 318062 551848 318118 551857
rect 318062 551783 318118 551792
rect 318076 551478 318104 551783
rect 318064 551472 318116 551478
rect 318064 551414 318116 551420
rect 317972 551404 318024 551410
rect 317972 551346 318024 551352
rect 318248 551268 318300 551274
rect 318248 551210 318300 551216
rect 318156 550860 318208 550866
rect 318156 550802 318208 550808
rect 318062 549944 318118 549953
rect 318062 549879 318118 549888
rect 316960 549500 317012 549506
rect 316960 549442 317012 549448
rect 316972 526386 317000 549442
rect 317972 547868 318024 547874
rect 317972 547810 318024 547816
rect 317984 547097 318012 547810
rect 317970 547088 318026 547097
rect 317970 547023 318026 547032
rect 317972 542360 318024 542366
rect 317970 542328 317972 542337
rect 318024 542328 318026 542337
rect 317970 542263 318026 542272
rect 318076 528086 318104 549879
rect 318064 528080 318116 528086
rect 318064 528022 318116 528028
rect 316960 526380 317012 526386
rect 316960 526322 317012 526328
rect 318168 525230 318196 550802
rect 318260 525570 318288 551210
rect 318340 550996 318392 551002
rect 318340 550938 318392 550944
rect 318248 525564 318300 525570
rect 318248 525506 318300 525512
rect 318156 525224 318208 525230
rect 318156 525166 318208 525172
rect 318352 524890 318380 550938
rect 318444 527814 318472 552094
rect 318536 527882 318564 552570
rect 319456 549982 319484 639270
rect 319548 554198 319576 640290
rect 319640 559638 319668 640970
rect 319812 640756 319864 640762
rect 319812 640698 319864 640704
rect 319718 640656 319774 640665
rect 319718 640591 319774 640600
rect 319732 562494 319760 640591
rect 319824 565214 319852 640698
rect 323860 640348 323912 640354
rect 323860 640290 323912 640296
rect 323872 638996 323900 640290
rect 328366 639296 328422 639305
rect 328366 639231 328422 639240
rect 328380 638996 328408 639231
rect 332888 638996 332916 641106
rect 337384 641096 337436 641102
rect 337384 641038 337436 641044
rect 337396 638996 337424 641038
rect 355416 641028 355468 641034
rect 355416 640970 355468 640976
rect 350908 640824 350960 640830
rect 350908 640766 350960 640772
rect 341892 639668 341944 639674
rect 341892 639610 341944 639616
rect 341904 638996 341932 639610
rect 346398 639160 346454 639169
rect 346398 639095 346454 639104
rect 346412 638996 346440 639095
rect 350920 638996 350948 640766
rect 355428 638996 355456 640970
rect 359924 640960 359976 640966
rect 359924 640902 359976 640908
rect 359936 638996 359964 640902
rect 364432 640892 364484 640898
rect 364432 640834 364484 640840
rect 364444 638996 364472 640834
rect 373448 640756 373500 640762
rect 373448 640698 373500 640704
rect 368940 640688 368992 640694
rect 368940 640630 368992 640636
rect 368952 638996 368980 640630
rect 373460 638996 373488 640698
rect 378612 638996 378640 641174
rect 392122 640656 392178 640665
rect 387616 640620 387668 640626
rect 392122 640591 392178 640600
rect 387616 640562 387668 640568
rect 383108 640552 383160 640558
rect 383108 640494 383160 640500
rect 383120 638996 383148 640494
rect 387628 638996 387656 640562
rect 392136 638996 392164 640591
rect 396632 640484 396684 640490
rect 396632 640426 396684 640432
rect 396644 638996 396672 640426
rect 401152 638996 401180 646478
rect 423680 643748 423732 643754
rect 423680 643690 423732 643696
rect 419170 640520 419226 640529
rect 419170 640455 419226 640464
rect 414664 640348 414716 640354
rect 414664 640290 414716 640296
rect 409880 639056 409932 639062
rect 405370 639024 405426 639033
rect 405426 638982 405674 639010
rect 414676 639010 414704 640290
rect 409932 639004 410182 639010
rect 409880 638998 410182 639004
rect 409892 638982 410182 638998
rect 414584 638996 414704 639010
rect 419184 638996 419212 640455
rect 423692 638996 423720 643690
rect 428188 640416 428240 640422
rect 428188 640358 428240 640364
rect 428200 638996 428228 640358
rect 428464 639600 428516 639606
rect 428464 639542 428516 639548
rect 414584 638994 414690 638996
rect 414572 638988 414690 638994
rect 405370 638959 405426 638968
rect 414624 638982 414690 638988
rect 414572 638930 414624 638936
rect 428476 629950 428504 639542
rect 428464 629944 428516 629950
rect 428464 629886 428516 629892
rect 428370 566264 428426 566273
rect 428370 566199 428426 566208
rect 319812 565208 319864 565214
rect 319812 565150 319864 565156
rect 319720 562488 319772 562494
rect 319720 562430 319772 562436
rect 319628 559632 319680 559638
rect 319628 559574 319680 559580
rect 319536 554192 319588 554198
rect 319536 554134 319588 554140
rect 319720 550180 319772 550186
rect 319720 550122 319772 550128
rect 319444 549976 319496 549982
rect 319444 549918 319496 549924
rect 319732 549930 319760 550122
rect 319812 550112 319864 550118
rect 319864 550060 319944 550066
rect 319812 550054 319944 550060
rect 319824 550038 319944 550054
rect 319732 549902 319852 549930
rect 319536 549432 319588 549438
rect 319536 549374 319588 549380
rect 318708 548616 318760 548622
rect 318708 548558 318760 548564
rect 318616 548548 318668 548554
rect 318616 548490 318668 548496
rect 318628 532817 318656 548490
rect 318720 537577 318748 548558
rect 319444 548140 319496 548146
rect 319444 548082 319496 548088
rect 318706 537568 318762 537577
rect 318706 537503 318762 537512
rect 318614 532808 318670 532817
rect 318614 532743 318670 532752
rect 318524 527876 318576 527882
rect 318524 527818 318576 527824
rect 318432 527808 318484 527814
rect 318432 527750 318484 527756
rect 319456 525094 319484 548082
rect 319548 526862 319576 549374
rect 319628 548208 319680 548214
rect 319628 548150 319680 548156
rect 319536 526856 319588 526862
rect 319536 526798 319588 526804
rect 319640 525774 319668 548150
rect 319720 548072 319772 548078
rect 319720 548014 319772 548020
rect 319628 525768 319680 525774
rect 319628 525710 319680 525716
rect 319732 525706 319760 548014
rect 319824 527950 319852 549902
rect 319916 528018 319944 550038
rect 427818 528592 427874 528601
rect 427818 528527 427874 528536
rect 320022 528278 320220 528306
rect 319904 528012 319956 528018
rect 319904 527954 319956 527960
rect 319812 527944 319864 527950
rect 319812 527886 319864 527892
rect 319720 525700 319772 525706
rect 319720 525642 319772 525648
rect 320088 525632 320140 525638
rect 320192 525620 320220 528278
rect 356086 528142 356284 528170
rect 324530 528006 324912 528034
rect 324884 526454 324912 528006
rect 328656 528006 329038 528034
rect 333256 528006 333546 528034
rect 337672 528006 338054 528034
rect 342272 528006 342562 528034
rect 346688 528006 347070 528034
rect 351288 528006 351578 528034
rect 324872 526448 324924 526454
rect 324872 526390 324924 526396
rect 328656 526250 328684 528006
rect 328644 526244 328696 526250
rect 328644 526186 328696 526192
rect 320456 525700 320508 525706
rect 320456 525642 320508 525648
rect 320140 525592 320220 525620
rect 320468 525586 320496 525642
rect 333256 525638 333284 528006
rect 337672 526318 337700 528006
rect 337660 526312 337712 526318
rect 337660 526254 337712 526260
rect 320088 525574 320140 525580
rect 320284 525570 320496 525586
rect 333244 525632 333296 525638
rect 333244 525574 333296 525580
rect 320272 525564 320496 525570
rect 320324 525558 320496 525564
rect 320548 525564 320600 525570
rect 320272 525506 320324 525512
rect 320548 525506 320600 525512
rect 320560 525450 320588 525506
rect 320376 525434 320588 525450
rect 320364 525428 320588 525434
rect 320416 525422 320588 525428
rect 320640 525428 320692 525434
rect 320364 525370 320416 525376
rect 320640 525370 320692 525376
rect 319444 525088 319496 525094
rect 319444 525030 319496 525036
rect 318340 524884 318392 524890
rect 318340 524826 318392 524832
rect 320652 524822 320680 525370
rect 342272 524958 342300 528006
rect 346688 525026 346716 528006
rect 351288 526386 351316 528006
rect 351276 526380 351328 526386
rect 351276 526322 351328 526328
rect 356256 525162 356284 528142
rect 360304 528006 360594 528034
rect 364720 528006 365102 528034
rect 369320 528006 369610 528034
rect 374472 528006 374762 528034
rect 378152 528006 379270 528034
rect 383672 528006 383778 528034
rect 387904 528006 388286 528034
rect 391952 528006 392794 528034
rect 396920 528006 397302 528034
rect 401612 528006 401810 528034
rect 405936 528006 406318 528034
rect 410536 528006 410826 528034
rect 414952 528006 415334 528034
rect 419552 528006 419842 528034
rect 423968 528006 424350 528034
rect 356244 525156 356296 525162
rect 356244 525098 356296 525104
rect 360304 525094 360332 528006
rect 364720 525298 364748 528006
rect 369320 527270 369348 528006
rect 369308 527264 369360 527270
rect 369308 527206 369360 527212
rect 364708 525292 364760 525298
rect 364708 525234 364760 525240
rect 374472 525230 374500 528006
rect 374460 525224 374512 525230
rect 374460 525166 374512 525172
rect 360292 525088 360344 525094
rect 360292 525030 360344 525036
rect 346676 525020 346728 525026
rect 346676 524962 346728 524968
rect 342260 524952 342312 524958
rect 342260 524894 342312 524900
rect 320640 524816 320692 524822
rect 320640 524758 320692 524764
rect 316868 522776 316920 522782
rect 316868 522718 316920 522724
rect 378152 486470 378180 528006
rect 383672 525366 383700 528006
rect 387904 525502 387932 528006
rect 387892 525496 387944 525502
rect 387892 525438 387944 525444
rect 383660 525360 383712 525366
rect 383660 525302 383712 525308
rect 391952 489161 391980 528006
rect 396920 527202 396948 528006
rect 396908 527196 396960 527202
rect 396908 527138 396960 527144
rect 401612 525434 401640 528006
rect 405936 525570 405964 528006
rect 405924 525564 405976 525570
rect 405924 525506 405976 525512
rect 401600 525428 401652 525434
rect 401600 525370 401652 525376
rect 410536 524890 410564 528006
rect 414952 526522 414980 528006
rect 414940 526516 414992 526522
rect 414940 526458 414992 526464
rect 419552 525706 419580 528006
rect 423968 525774 423996 528006
rect 423956 525768 424008 525774
rect 423956 525710 424008 525716
rect 419540 525700 419592 525706
rect 419540 525642 419592 525648
rect 410524 524884 410576 524890
rect 410524 524826 410576 524832
rect 427832 522782 427860 528527
rect 428384 527814 428412 566199
rect 428372 527808 428424 527814
rect 428372 527750 428424 527756
rect 429212 526454 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429384 647896 429436 647902
rect 429384 647838 429436 647844
rect 429290 591288 429346 591297
rect 429290 591223 429346 591232
rect 429200 526448 429252 526454
rect 429200 526390 429252 526396
rect 427820 522776 427872 522782
rect 427820 522718 427872 522724
rect 391938 489152 391994 489161
rect 391938 489087 391994 489096
rect 378140 486464 378192 486470
rect 378140 486406 378192 486412
rect 356796 485580 356848 485586
rect 356796 485522 356848 485528
rect 356704 485308 356756 485314
rect 356704 485250 356756 485256
rect 316776 483676 316828 483682
rect 316776 483618 316828 483624
rect 312542 482216 312598 482225
rect 312542 482151 312598 482160
rect 299480 471232 299532 471238
rect 298190 471200 298246 471209
rect 299480 471174 299532 471180
rect 298190 471135 298246 471144
rect 339408 466608 339460 466614
rect 338486 466576 338542 466585
rect 339408 466550 339460 466556
rect 339774 466576 339830 466585
rect 338486 466511 338542 466520
rect 338500 466478 338528 466511
rect 339420 466478 339448 466550
rect 339774 466511 339776 466520
rect 339828 466511 339830 466520
rect 350998 466576 351054 466585
rect 350998 466511 351054 466520
rect 339776 466482 339828 466488
rect 351012 466478 351040 466511
rect 338488 466472 338540 466478
rect 338488 466414 338540 466420
rect 339408 466472 339460 466478
rect 339408 466414 339460 466420
rect 351000 466472 351052 466478
rect 351000 466414 351052 466420
rect 298100 465588 298152 465594
rect 298100 465530 298152 465536
rect 287060 464500 287112 464506
rect 287060 464442 287112 464448
rect 271880 464432 271932 464438
rect 271880 464374 271932 464380
rect 264980 464364 265032 464370
rect 264980 464306 265032 464312
rect 276020 380928 276072 380934
rect 235998 380896 236054 380905
rect 235998 380831 236054 380840
rect 237102 380896 237158 380905
rect 237102 380831 237158 380840
rect 243082 380896 243138 380905
rect 243082 380831 243138 380840
rect 245382 380896 245438 380905
rect 245382 380831 245438 380840
rect 247590 380896 247646 380905
rect 247590 380831 247646 380840
rect 254490 380896 254546 380905
rect 254490 380831 254546 380840
rect 255870 380896 255926 380905
rect 255870 380831 255926 380840
rect 256974 380896 257030 380905
rect 256974 380831 257030 380840
rect 276018 380896 276020 380905
rect 276072 380896 276074 380905
rect 276018 380831 276074 380840
rect 236012 380050 236040 380831
rect 236000 380044 236052 380050
rect 236000 379986 236052 379992
rect 237116 379982 237144 380831
rect 237104 379976 237156 379982
rect 237104 379918 237156 379924
rect 239956 379976 240008 379982
rect 239956 379918 240008 379924
rect 220728 379772 220780 379778
rect 220728 379714 220780 379720
rect 220740 379642 220768 379714
rect 220728 379636 220780 379642
rect 220728 379578 220780 379584
rect 221832 379568 221884 379574
rect 221832 379510 221884 379516
rect 220636 379500 220688 379506
rect 220636 379442 220688 379448
rect 220544 379296 220596 379302
rect 220544 379238 220596 379244
rect 220176 379160 220228 379166
rect 220176 379102 220228 379108
rect 220452 379160 220504 379166
rect 220452 379102 220504 379108
rect 220188 378690 220216 379102
rect 220176 378684 220228 378690
rect 220176 378626 220228 378632
rect 220464 378214 220492 379102
rect 220556 378554 220584 379238
rect 220648 378758 220676 379442
rect 220728 379364 220780 379370
rect 220728 379306 220780 379312
rect 220740 378962 220768 379306
rect 220820 379228 220872 379234
rect 220820 379170 220872 379176
rect 220728 378956 220780 378962
rect 220728 378898 220780 378904
rect 220636 378752 220688 378758
rect 220636 378694 220688 378700
rect 220544 378548 220596 378554
rect 220544 378490 220596 378496
rect 220452 378208 220504 378214
rect 220452 378150 220504 378156
rect 220832 358630 220860 379170
rect 221556 379092 221608 379098
rect 221556 379034 221608 379040
rect 220912 379024 220964 379030
rect 220912 378966 220964 378972
rect 220924 358698 220952 378966
rect 221002 378720 221058 378729
rect 221002 378655 221058 378664
rect 220912 358692 220964 358698
rect 220912 358634 220964 358640
rect 220820 358624 220872 358630
rect 220820 358566 220872 358572
rect 221016 358562 221044 378655
rect 221568 378622 221596 379034
rect 221646 378856 221702 378865
rect 221646 378791 221702 378800
rect 221096 378616 221148 378622
rect 221556 378616 221608 378622
rect 221096 378558 221148 378564
rect 221278 378584 221334 378593
rect 221004 358556 221056 358562
rect 221004 358498 221056 358504
rect 221108 358290 221136 378558
rect 221556 378558 221608 378564
rect 221278 378519 221334 378528
rect 221186 378312 221242 378321
rect 221186 378247 221242 378256
rect 221096 358284 221148 358290
rect 221096 358226 221148 358232
rect 221200 358154 221228 378247
rect 221188 358148 221240 358154
rect 221188 358090 221240 358096
rect 221292 357542 221320 378519
rect 221660 378321 221688 378791
rect 221646 378312 221702 378321
rect 221646 378247 221702 378256
rect 221844 377777 221872 379510
rect 221924 379228 221976 379234
rect 221924 379170 221976 379176
rect 221936 378350 221964 379170
rect 222014 379128 222070 379137
rect 222014 379063 222070 379072
rect 222028 378729 222056 379063
rect 222108 379024 222160 379030
rect 222108 378966 222160 378972
rect 222014 378720 222070 378729
rect 222014 378655 222070 378664
rect 221924 378344 221976 378350
rect 221924 378286 221976 378292
rect 222120 378214 222148 378966
rect 233882 378720 233938 378729
rect 233882 378655 233938 378664
rect 233896 378457 233924 378655
rect 233882 378448 233938 378457
rect 233882 378383 233938 378392
rect 222108 378208 222160 378214
rect 222108 378150 222160 378156
rect 221370 377768 221426 377777
rect 221370 377703 221426 377712
rect 221830 377768 221886 377777
rect 221830 377703 221886 377712
rect 221384 358766 221412 377703
rect 239968 375834 239996 379918
rect 243096 379846 243124 380831
rect 244278 380352 244334 380361
rect 244278 380287 244334 380296
rect 244292 379914 244320 380287
rect 244280 379908 244332 379914
rect 244280 379850 244332 379856
rect 243084 379840 243136 379846
rect 243084 379782 243136 379788
rect 245396 378894 245424 380831
rect 245658 379264 245714 379273
rect 245658 379199 245714 379208
rect 245384 378888 245436 378894
rect 245384 378830 245436 378836
rect 245672 378418 245700 379199
rect 247604 378962 247632 380831
rect 254504 379778 254532 380831
rect 254492 379772 254544 379778
rect 254492 379714 254544 379720
rect 255884 379642 255912 380831
rect 256988 379710 257016 380831
rect 259458 380624 259514 380633
rect 259458 380559 259514 380568
rect 265254 380624 265310 380633
rect 265254 380559 265310 380568
rect 270958 380624 271014 380633
rect 270958 380559 271014 380568
rect 259472 379982 259500 380559
rect 259460 379976 259512 379982
rect 259460 379918 259512 379924
rect 256976 379704 257028 379710
rect 256976 379646 257028 379652
rect 255872 379636 255924 379642
rect 255872 379578 255924 379584
rect 265268 379574 265296 380559
rect 265256 379568 265308 379574
rect 265256 379510 265308 379516
rect 268658 379400 268714 379409
rect 268658 379335 268714 379344
rect 248602 379264 248658 379273
rect 248602 379199 248658 379208
rect 250074 379264 250130 379273
rect 250074 379199 250130 379208
rect 251178 379264 251234 379273
rect 251178 379199 251234 379208
rect 252282 379264 252338 379273
rect 252282 379199 252338 379208
rect 253386 379264 253442 379273
rect 253386 379199 253442 379208
rect 261666 379264 261722 379273
rect 261666 379199 261722 379208
rect 247592 378956 247644 378962
rect 247592 378898 247644 378904
rect 248616 378690 248644 379199
rect 248604 378684 248656 378690
rect 248604 378626 248656 378632
rect 250088 378554 250116 379199
rect 251192 378622 251220 379199
rect 251180 378616 251232 378622
rect 251180 378558 251232 378564
rect 250076 378548 250128 378554
rect 250076 378490 250128 378496
rect 248234 378448 248290 378457
rect 245660 378412 245712 378418
rect 248234 378383 248290 378392
rect 250626 378448 250682 378457
rect 250626 378383 250682 378392
rect 245660 378354 245712 378360
rect 248248 376106 248276 378383
rect 248236 376100 248288 376106
rect 248236 376042 248288 376048
rect 250640 375902 250668 378383
rect 252296 378350 252324 379199
rect 253202 379128 253258 379137
rect 253202 379063 253258 379072
rect 252284 378344 252336 378350
rect 253216 378321 253244 379063
rect 252284 378286 252336 378292
rect 253202 378312 253258 378321
rect 253202 378247 253258 378256
rect 253400 378214 253428 379199
rect 253570 378448 253626 378457
rect 253570 378383 253626 378392
rect 255962 378448 256018 378457
rect 255962 378383 256018 378392
rect 258354 378448 258410 378457
rect 258354 378383 258410 378392
rect 260930 378448 260986 378457
rect 260930 378383 260986 378392
rect 253388 378208 253440 378214
rect 253388 378150 253440 378156
rect 253584 375970 253612 378383
rect 255976 376038 256004 378383
rect 258368 376242 258396 378383
rect 260944 376310 260972 378383
rect 260932 376304 260984 376310
rect 260932 376246 260984 376252
rect 258356 376236 258408 376242
rect 258356 376178 258408 376184
rect 255964 376032 256016 376038
rect 255964 375974 256016 375980
rect 253572 375964 253624 375970
rect 253572 375906 253624 375912
rect 250628 375896 250680 375902
rect 250628 375838 250680 375844
rect 239956 375828 240008 375834
rect 239956 375770 240008 375776
rect 261680 375154 261708 379199
rect 268672 378826 268700 379335
rect 268660 378820 268712 378826
rect 268660 378762 268712 378768
rect 263598 378448 263654 378457
rect 263598 378383 263654 378392
rect 265346 378448 265402 378457
rect 265346 378383 265402 378392
rect 268106 378448 268162 378457
rect 268106 378383 268162 378392
rect 262770 378312 262826 378321
rect 262770 378247 262826 378256
rect 262784 375290 262812 378247
rect 263612 376446 263640 378383
rect 263600 376440 263652 376446
rect 263600 376382 263652 376388
rect 265360 376174 265388 378383
rect 266358 378312 266414 378321
rect 266358 378247 266414 378256
rect 267554 378312 267610 378321
rect 267554 378247 267610 378256
rect 265348 376168 265400 376174
rect 265348 376110 265400 376116
rect 266372 375358 266400 378247
rect 266360 375352 266412 375358
rect 266360 375294 266412 375300
rect 262772 375284 262824 375290
rect 262772 375226 262824 375232
rect 261668 375148 261720 375154
rect 261668 375090 261720 375096
rect 267568 374746 267596 378247
rect 268120 376378 268148 378383
rect 270972 376514 271000 380559
rect 274640 380452 274692 380458
rect 274640 380394 274692 380400
rect 274652 379506 274680 380394
rect 295340 380316 295392 380322
rect 295340 380258 295392 380264
rect 274640 379500 274692 379506
rect 274640 379442 274692 379448
rect 295352 379438 295380 380258
rect 301504 380248 301556 380254
rect 301504 380190 301556 380196
rect 273260 379432 273312 379438
rect 271050 379400 271106 379409
rect 271050 379335 271106 379344
rect 271970 379400 272026 379409
rect 271970 379335 272026 379344
rect 273258 379400 273260 379409
rect 275652 379432 275704 379438
rect 273312 379400 273314 379409
rect 273258 379335 273314 379344
rect 274362 379400 274418 379409
rect 274362 379335 274364 379344
rect 271064 378486 271092 379335
rect 271052 378480 271104 378486
rect 271052 378422 271104 378428
rect 271984 378282 272012 379335
rect 274416 379335 274418 379344
rect 275650 379400 275652 379409
rect 295340 379432 295392 379438
rect 275704 379400 275706 379409
rect 275650 379335 275706 379344
rect 285954 379400 286010 379409
rect 285954 379335 286010 379344
rect 287610 379400 287666 379409
rect 287610 379335 287666 379344
rect 290922 379400 290978 379409
rect 290922 379335 290978 379344
rect 293314 379400 293370 379409
rect 295340 379374 295392 379380
rect 295890 379400 295946 379409
rect 293314 379335 293370 379344
rect 295890 379335 295946 379344
rect 298098 379400 298154 379409
rect 298098 379335 298154 379344
rect 300858 379400 300914 379409
rect 301516 379370 301544 380190
rect 311808 380180 311860 380186
rect 311808 380122 311860 380128
rect 311820 379438 311848 380122
rect 323308 379500 323360 379506
rect 323308 379442 323360 379448
rect 310980 379432 311032 379438
rect 303066 379400 303122 379409
rect 300858 379335 300914 379344
rect 301504 379364 301556 379370
rect 274364 379306 274416 379312
rect 273442 379264 273498 379273
rect 273442 379199 273498 379208
rect 277030 379264 277086 379273
rect 277030 379199 277086 379208
rect 277858 379264 277914 379273
rect 277858 379199 277914 379208
rect 279146 379264 279202 379273
rect 279146 379199 279202 379208
rect 280802 379264 280858 379273
rect 280802 379199 280858 379208
rect 283010 379264 283066 379273
rect 283010 379199 283066 379208
rect 271972 378276 272024 378282
rect 271972 378218 272024 378224
rect 273260 378208 273312 378214
rect 273260 378150 273312 378156
rect 273272 378049 273300 378150
rect 273258 378040 273314 378049
rect 273258 377975 273314 377984
rect 273456 376582 273484 379199
rect 277044 378282 277072 379199
rect 276020 378276 276072 378282
rect 276020 378218 276072 378224
rect 277032 378276 277084 378282
rect 277032 378218 277084 378224
rect 276032 378185 276060 378218
rect 276018 378176 276074 378185
rect 276018 378111 276074 378120
rect 277872 377466 277900 379199
rect 277860 377460 277912 377466
rect 277860 377402 277912 377408
rect 273444 376576 273496 376582
rect 273444 376518 273496 376524
rect 270960 376508 271012 376514
rect 270960 376450 271012 376456
rect 268108 376372 268160 376378
rect 268108 376314 268160 376320
rect 279160 375222 279188 379199
rect 280816 377398 280844 379199
rect 280804 377392 280856 377398
rect 280804 377334 280856 377340
rect 283024 376718 283052 379199
rect 285968 377602 285996 379335
rect 287624 378146 287652 379335
rect 287612 378140 287664 378146
rect 287612 378082 287664 378088
rect 290936 377670 290964 379335
rect 293328 377738 293356 379335
rect 295904 377806 295932 379335
rect 298112 377874 298140 379335
rect 300872 377942 300900 379335
rect 303066 379335 303122 379344
rect 305734 379400 305790 379409
rect 305734 379335 305790 379344
rect 308402 379400 308458 379409
rect 308402 379335 308458 379344
rect 310978 379400 310980 379409
rect 311808 379432 311860 379438
rect 311032 379400 311034 379409
rect 315764 379432 315816 379438
rect 311808 379374 311860 379380
rect 313370 379400 313426 379409
rect 310978 379335 311034 379344
rect 313370 379335 313372 379344
rect 301504 379306 301556 379312
rect 303080 378214 303108 379335
rect 303068 378208 303120 378214
rect 303068 378150 303120 378156
rect 300860 377936 300912 377942
rect 300860 377878 300912 377884
rect 298100 377868 298152 377874
rect 298100 377810 298152 377816
rect 295892 377800 295944 377806
rect 295892 377742 295944 377748
rect 293316 377732 293368 377738
rect 293316 377674 293368 377680
rect 290924 377664 290976 377670
rect 290924 377606 290976 377612
rect 285956 377596 286008 377602
rect 285956 377538 286008 377544
rect 305748 377534 305776 379335
rect 308416 378078 308444 379335
rect 313424 379335 313426 379344
rect 315762 379400 315764 379409
rect 323320 379409 323348 379442
rect 315816 379400 315818 379409
rect 315762 379335 315818 379344
rect 318338 379400 318394 379409
rect 318338 379335 318394 379344
rect 323306 379400 323362 379409
rect 323306 379335 323362 379344
rect 313372 379306 313424 379312
rect 308404 378072 308456 378078
rect 308404 378014 308456 378020
rect 318352 378010 318380 379335
rect 325882 379264 325938 379273
rect 325882 379199 325938 379208
rect 320914 378584 320970 378593
rect 320914 378519 320970 378528
rect 318340 378004 318392 378010
rect 318340 377946 318392 377952
rect 305736 377528 305788 377534
rect 305736 377470 305788 377476
rect 283012 376712 283064 376718
rect 283012 376654 283064 376660
rect 320928 376650 320956 378519
rect 320916 376644 320968 376650
rect 320916 376586 320968 376592
rect 325896 375329 325924 379199
rect 343178 378448 343234 378457
rect 343178 378383 343234 378392
rect 343192 378350 343220 378383
rect 342260 378344 342312 378350
rect 342260 378286 342312 378292
rect 343180 378344 343232 378350
rect 343180 378286 343232 378292
rect 343546 378312 343602 378321
rect 325882 375320 325938 375329
rect 325882 375255 325938 375264
rect 279148 375216 279200 375222
rect 279148 375158 279200 375164
rect 267556 374740 267608 374746
rect 267556 374682 267608 374688
rect 342272 374678 342300 378286
rect 343546 378247 343602 378256
rect 356612 378276 356664 378282
rect 343560 378214 343588 378247
rect 356612 378218 356664 378224
rect 343548 378208 343600 378214
rect 343548 378150 343600 378156
rect 342260 374672 342312 374678
rect 342260 374614 342312 374620
rect 339868 359576 339920 359582
rect 339868 359518 339920 359524
rect 339880 358873 339908 359518
rect 343560 358902 343588 378150
rect 351736 359508 351788 359514
rect 351736 359450 351788 359456
rect 342260 358896 342312 358902
rect 338486 358864 338542 358873
rect 338486 358799 338488 358808
rect 338540 358799 338542 358808
rect 339866 358864 339922 358873
rect 342260 358838 342312 358844
rect 343548 358896 343600 358902
rect 351748 358873 351776 359450
rect 343548 358838 343600 358844
rect 351734 358864 351790 358873
rect 339866 358799 339922 358808
rect 338488 358770 338540 358776
rect 221372 358760 221424 358766
rect 221372 358702 221424 358708
rect 342272 358086 342300 358838
rect 351734 358799 351790 358808
rect 342260 358080 342312 358086
rect 342260 358022 342312 358028
rect 221280 357536 221332 357542
rect 221280 357478 221332 357484
rect 266358 273728 266414 273737
rect 266358 273663 266414 273672
rect 278042 273728 278098 273737
rect 278042 273663 278098 273672
rect 266372 273630 266400 273663
rect 266360 273624 266412 273630
rect 250718 273592 250774 273601
rect 266360 273566 266412 273572
rect 273350 273592 273406 273601
rect 250718 273527 250720 273536
rect 250772 273527 250774 273536
rect 273350 273527 273406 273536
rect 275742 273592 275798 273601
rect 275742 273527 275798 273536
rect 250720 273498 250772 273504
rect 273364 273494 273392 273527
rect 273352 273488 273404 273494
rect 273352 273430 273404 273436
rect 275756 273426 275784 273527
rect 275744 273420 275796 273426
rect 275744 273362 275796 273368
rect 278056 273358 278084 273663
rect 283470 273592 283526 273601
rect 283470 273527 283526 273536
rect 278044 273352 278096 273358
rect 278044 273294 278096 273300
rect 283484 273290 283512 273527
rect 285954 273320 286010 273329
rect 283472 273284 283524 273290
rect 285954 273255 286010 273264
rect 283472 273226 283524 273232
rect 285968 272950 285996 273255
rect 288164 273012 288216 273018
rect 288164 272954 288216 272960
rect 285956 272944 286008 272950
rect 288176 272921 288204 272954
rect 285956 272886 286008 272892
rect 287978 272912 288034 272921
rect 287978 272847 288034 272856
rect 288162 272912 288218 272921
rect 288162 272847 288218 272856
rect 290922 272912 290978 272921
rect 290922 272847 290924 272856
rect 287992 272649 288020 272847
rect 290976 272847 290978 272856
rect 293314 272912 293370 272921
rect 293314 272847 293370 272856
rect 300858 272912 300914 272921
rect 300858 272847 300914 272856
rect 290924 272818 290976 272824
rect 293328 272746 293356 272847
rect 300872 272814 300900 272847
rect 300860 272808 300912 272814
rect 298466 272776 298522 272785
rect 293316 272740 293368 272746
rect 300860 272750 300912 272756
rect 298466 272711 298522 272720
rect 293316 272682 293368 272688
rect 298480 272678 298508 272711
rect 298468 272672 298520 272678
rect 287978 272640 288034 272649
rect 298468 272614 298520 272620
rect 305826 272640 305882 272649
rect 287978 272575 288034 272584
rect 305826 272575 305828 272584
rect 305880 272575 305882 272584
rect 320914 272640 320970 272649
rect 320914 272575 320970 272584
rect 305828 272546 305880 272552
rect 320928 272542 320956 272575
rect 320916 272536 320968 272542
rect 320916 272478 320968 272484
rect 235998 272232 236054 272241
rect 235998 272167 236054 272176
rect 265162 272232 265218 272241
rect 265162 272167 265218 272176
rect 236012 271998 236040 272167
rect 236000 271992 236052 271998
rect 236000 271934 236052 271940
rect 258262 271552 258318 271561
rect 258262 271487 258318 271496
rect 263598 271552 263654 271561
rect 263598 271487 263654 271496
rect 264978 271552 265034 271561
rect 264978 271487 264980 271496
rect 252558 271280 252614 271289
rect 252558 271215 252614 271224
rect 252572 271182 252600 271215
rect 252560 271176 252612 271182
rect 247038 271144 247094 271153
rect 252560 271118 252612 271124
rect 255318 271144 255374 271153
rect 247038 271079 247094 271088
rect 258276 271114 258304 271487
rect 263612 271318 263640 271487
rect 265032 271487 265034 271496
rect 264980 271458 265032 271464
rect 263600 271312 263652 271318
rect 260838 271280 260894 271289
rect 263600 271254 263652 271260
rect 260838 271215 260840 271224
rect 260892 271215 260894 271224
rect 260840 271186 260892 271192
rect 255318 271079 255374 271088
rect 258264 271108 258316 271114
rect 247052 270978 247080 271079
rect 255332 271046 255360 271079
rect 258264 271050 258316 271056
rect 255320 271040 255372 271046
rect 255320 270982 255372 270988
rect 247040 270972 247092 270978
rect 247040 270914 247092 270920
rect 253938 270872 253994 270881
rect 253938 270807 253994 270816
rect 244370 270736 244426 270745
rect 244370 270671 244426 270680
rect 251270 270736 251326 270745
rect 251270 270671 251326 270680
rect 239126 270600 239182 270609
rect 239126 270535 239182 270544
rect 242898 270600 242954 270609
rect 242898 270535 242954 270544
rect 244278 270600 244334 270609
rect 244278 270535 244334 270544
rect 220636 270496 220688 270502
rect 220636 270438 220688 270444
rect 220648 269482 220676 270438
rect 220728 270292 220780 270298
rect 220728 270234 220780 270240
rect 220740 270162 220768 270234
rect 220728 270156 220780 270162
rect 220728 270098 220780 270104
rect 224224 270156 224276 270162
rect 224224 270098 224276 270104
rect 224132 269952 224184 269958
rect 224132 269894 224184 269900
rect 224144 269686 224172 269894
rect 224236 269890 224264 270098
rect 224408 269952 224460 269958
rect 224408 269894 224460 269900
rect 224224 269884 224276 269890
rect 224224 269826 224276 269832
rect 224316 269884 224368 269890
rect 224316 269826 224368 269832
rect 224132 269680 224184 269686
rect 224132 269622 224184 269628
rect 224328 269550 224356 269826
rect 224316 269544 224368 269550
rect 224316 269486 224368 269492
rect 220636 269476 220688 269482
rect 220636 269418 220688 269424
rect 224420 269278 224448 269894
rect 239140 269754 239168 270535
rect 239128 269748 239180 269754
rect 239128 269690 239180 269696
rect 224408 269272 224460 269278
rect 224408 269214 224460 269220
rect 242912 269006 242940 270535
rect 244292 269686 244320 270535
rect 244280 269680 244332 269686
rect 244280 269622 244332 269628
rect 242900 269000 242952 269006
rect 242900 268942 242952 268948
rect 231860 268932 231912 268938
rect 231860 268874 231912 268880
rect 230480 268864 230532 268870
rect 230480 268806 230532 268812
rect 229192 268796 229244 268802
rect 229192 268738 229244 268744
rect 229204 268433 229232 268738
rect 229190 268424 229246 268433
rect 229190 268359 229246 268368
rect 229204 258074 229232 268359
rect 229112 258046 229232 258074
rect 229112 251938 229140 258046
rect 229100 251932 229152 251938
rect 229100 251874 229152 251880
rect 230492 251870 230520 268806
rect 231872 268326 231900 268874
rect 231860 268320 231912 268326
rect 231860 268262 231912 268268
rect 230480 251864 230532 251870
rect 231872 251841 231900 268262
rect 244384 268258 244412 270671
rect 245658 270600 245714 270609
rect 245658 270535 245714 270544
rect 247038 270600 247094 270609
rect 247038 270535 247094 270544
rect 248510 270600 248566 270609
rect 248510 270535 248566 270544
rect 249798 270600 249854 270609
rect 249798 270535 249854 270544
rect 251178 270600 251234 270609
rect 251178 270535 251234 270544
rect 245672 270162 245700 270535
rect 247052 270502 247080 270535
rect 247040 270496 247092 270502
rect 247040 270438 247092 270444
rect 248524 270230 248552 270535
rect 249812 270298 249840 270535
rect 251192 270366 251220 270535
rect 251180 270360 251232 270366
rect 251180 270302 251232 270308
rect 249800 270292 249852 270298
rect 249800 270234 249852 270240
rect 248512 270224 248564 270230
rect 248512 270166 248564 270172
rect 245660 270156 245712 270162
rect 245660 270098 245712 270104
rect 251284 270094 251312 270671
rect 252558 270600 252614 270609
rect 252558 270535 252614 270544
rect 251272 270088 251324 270094
rect 251272 270030 251324 270036
rect 252572 270026 252600 270535
rect 252560 270020 252612 270026
rect 252560 269962 252612 269968
rect 253952 269074 253980 270807
rect 255318 270736 255374 270745
rect 255318 270671 255374 270680
rect 259550 270736 259606 270745
rect 259550 270671 259606 270680
rect 253940 269068 253992 269074
rect 253940 269010 253992 269016
rect 255332 268734 255360 270671
rect 256698 270600 256754 270609
rect 256698 270535 256754 270544
rect 258078 270600 258134 270609
rect 258078 270535 258134 270544
rect 259458 270600 259514 270609
rect 259458 270535 259514 270544
rect 255320 268728 255372 268734
rect 255320 268670 255372 268676
rect 256712 268598 256740 270535
rect 258092 268666 258120 270535
rect 259472 268938 259500 270535
rect 259460 268932 259512 268938
rect 259460 268874 259512 268880
rect 259564 268870 259592 270671
rect 260838 270600 260894 270609
rect 260838 270535 260894 270544
rect 262218 270600 262274 270609
rect 262218 270535 262274 270544
rect 263598 270600 263654 270609
rect 263598 270535 263654 270544
rect 259552 268864 259604 268870
rect 259552 268806 259604 268812
rect 260852 268802 260880 270535
rect 262232 269890 262260 270535
rect 263612 270434 263640 270535
rect 263600 270428 263652 270434
rect 263600 270370 263652 270376
rect 265176 269958 265204 272167
rect 268200 271924 268252 271930
rect 268200 271866 268252 271872
rect 268212 271833 268240 271866
rect 313280 271856 313332 271862
rect 268198 271824 268254 271833
rect 268198 271759 268254 271768
rect 270498 271824 270554 271833
rect 270498 271759 270554 271768
rect 276018 271824 276074 271833
rect 276018 271759 276074 271768
rect 280158 271824 280214 271833
rect 280158 271759 280214 271768
rect 307758 271824 307814 271833
rect 307758 271759 307760 271768
rect 268016 271720 268068 271726
rect 268016 271662 268068 271668
rect 268028 271561 268056 271662
rect 268014 271552 268070 271561
rect 268014 271487 268070 271496
rect 270512 271454 270540 271759
rect 276032 271590 276060 271759
rect 280172 271658 280200 271759
rect 307812 271759 307814 271768
rect 313278 271824 313280 271833
rect 343548 271856 343600 271862
rect 313332 271824 313334 271833
rect 313278 271759 313334 271768
rect 343546 271824 343548 271833
rect 343600 271824 343602 271833
rect 343546 271759 343602 271768
rect 307760 271730 307812 271736
rect 280160 271652 280212 271658
rect 280160 271594 280212 271600
rect 276020 271584 276072 271590
rect 271878 271552 271934 271561
rect 276020 271526 276072 271532
rect 277122 271552 277178 271561
rect 271878 271487 271934 271496
rect 277122 271487 277178 271496
rect 343546 271552 343602 271561
rect 343546 271487 343602 271496
rect 270500 271448 270552 271454
rect 270500 271390 270552 271396
rect 266358 270600 266414 270609
rect 266358 270535 266414 270544
rect 269118 270600 269174 270609
rect 269118 270535 269174 270544
rect 270498 270600 270554 270609
rect 270498 270535 270554 270544
rect 265164 269952 265216 269958
rect 265164 269894 265216 269900
rect 262220 269884 262272 269890
rect 262220 269826 262272 269832
rect 266372 269822 266400 270535
rect 266360 269816 266412 269822
rect 266360 269758 266412 269764
rect 260840 268796 260892 268802
rect 260840 268738 260892 268744
rect 258080 268660 258132 268666
rect 258080 268602 258132 268608
rect 256700 268592 256752 268598
rect 256700 268534 256752 268540
rect 269132 268530 269160 270535
rect 269120 268524 269172 268530
rect 269120 268466 269172 268472
rect 270512 268462 270540 270535
rect 271892 269618 271920 271487
rect 277136 271182 277164 271487
rect 277674 271416 277730 271425
rect 277674 271351 277676 271360
rect 277728 271351 277730 271360
rect 277676 271322 277728 271328
rect 343560 271250 343588 271487
rect 343548 271244 343600 271250
rect 343548 271186 343600 271192
rect 356624 271182 356652 378218
rect 277124 271176 277176 271182
rect 277124 271118 277176 271124
rect 356612 271176 356664 271182
rect 356612 271118 356664 271124
rect 280066 270872 280122 270881
rect 280066 270807 280122 270816
rect 273166 270600 273222 270609
rect 273166 270535 273222 270544
rect 271880 269612 271932 269618
rect 271880 269554 271932 269560
rect 270500 268456 270552 268462
rect 270500 268398 270552 268404
rect 273180 268394 273208 270535
rect 280080 270502 280108 270807
rect 280068 270496 280120 270502
rect 280068 270438 280120 270444
rect 356612 270496 356664 270502
rect 356612 270438 356664 270444
rect 273168 268388 273220 268394
rect 273168 268330 273220 268336
rect 244372 268252 244424 268258
rect 244372 268194 244424 268200
rect 340788 253904 340840 253910
rect 340788 253846 340840 253852
rect 340800 253473 340828 253846
rect 340786 253464 340842 253473
rect 340786 253399 340842 253408
rect 339408 253292 339460 253298
rect 339408 253234 339460 253240
rect 339420 253065 339448 253234
rect 351828 253224 351880 253230
rect 351826 253192 351828 253201
rect 351880 253192 351882 253201
rect 351826 253127 351882 253136
rect 339406 253056 339462 253065
rect 339406 252991 339462 253000
rect 230480 251806 230532 251812
rect 231858 251832 231914 251841
rect 231858 251767 231914 251776
rect 260932 166864 260984 166870
rect 260932 166806 260984 166812
rect 260944 166569 260972 166806
rect 265900 166796 265952 166802
rect 265900 166738 265952 166744
rect 265912 166569 265940 166738
rect 270868 166728 270920 166734
rect 270868 166670 270920 166676
rect 285954 166696 286010 166705
rect 270880 166569 270908 166670
rect 285954 166631 285956 166640
rect 286008 166631 286010 166640
rect 291014 166696 291070 166705
rect 291014 166631 291070 166640
rect 293406 166696 293462 166705
rect 293406 166631 293462 166640
rect 295890 166696 295946 166705
rect 295890 166631 295946 166640
rect 298466 166696 298522 166705
rect 298466 166631 298522 166640
rect 305918 166696 305974 166705
rect 305918 166631 305974 166640
rect 285956 166602 286008 166608
rect 260930 166560 260986 166569
rect 260930 166495 260986 166504
rect 265898 166560 265954 166569
rect 265898 166495 265954 166504
rect 270866 166560 270922 166569
rect 270866 166495 270922 166504
rect 291028 166462 291056 166631
rect 293420 166530 293448 166631
rect 295904 166598 295932 166631
rect 295892 166592 295944 166598
rect 295892 166534 295944 166540
rect 293408 166524 293460 166530
rect 293408 166466 293460 166472
rect 291016 166456 291068 166462
rect 291016 166398 291068 166404
rect 298480 166394 298508 166631
rect 298468 166388 298520 166394
rect 298468 166330 298520 166336
rect 305932 166326 305960 166631
rect 305920 166320 305972 166326
rect 305920 166262 305972 166268
rect 235998 165608 236054 165617
rect 235998 165543 236054 165552
rect 238758 165608 238814 165617
rect 238758 165543 238814 165552
rect 242898 165608 242954 165617
rect 242898 165543 242954 165552
rect 247038 165608 247094 165617
rect 247038 165543 247094 165552
rect 247682 165608 247738 165617
rect 247682 165543 247738 165552
rect 249798 165608 249854 165617
rect 249798 165543 249854 165552
rect 252558 165608 252614 165617
rect 252558 165543 252614 165552
rect 258078 165608 258134 165617
rect 258078 165543 258134 165552
rect 260838 165608 260894 165617
rect 260838 165543 260894 165552
rect 264978 165608 265034 165617
rect 264978 165543 265034 165552
rect 267646 165608 267702 165617
rect 267922 165608 267978 165617
rect 267702 165566 267872 165594
rect 267646 165543 267702 165552
rect 236012 164014 236040 165543
rect 236090 164248 236146 164257
rect 236090 164183 236146 164192
rect 237378 164248 237434 164257
rect 237378 164183 237434 164192
rect 236104 164082 236132 164183
rect 236092 164076 236144 164082
rect 236092 164018 236144 164024
rect 236000 164008 236052 164014
rect 236000 163950 236052 163956
rect 235264 161560 235316 161566
rect 235264 161502 235316 161508
rect 235276 146266 235304 161502
rect 235264 146260 235316 146266
rect 235264 146202 235316 146208
rect 220082 145752 220138 145761
rect 220082 145687 220138 145696
rect 220096 143342 220124 145687
rect 236012 145450 236040 163950
rect 236104 145518 236132 164018
rect 236644 161492 236696 161498
rect 236644 161434 236696 161440
rect 236656 146198 236684 161434
rect 236644 146192 236696 146198
rect 236644 146134 236696 146140
rect 237392 145897 237420 164183
rect 238772 148714 238800 165543
rect 240138 164248 240194 164257
rect 240138 164183 240194 164192
rect 241518 164248 241574 164257
rect 241518 164183 241574 164192
rect 240152 148918 240180 164183
rect 240140 148912 240192 148918
rect 240140 148854 240192 148860
rect 238760 148708 238812 148714
rect 238760 148650 238812 148656
rect 241532 148646 241560 164183
rect 241520 148640 241572 148646
rect 241520 148582 241572 148588
rect 237378 145888 237434 145897
rect 237378 145823 237434 145832
rect 242912 145654 242940 165543
rect 244278 164520 244334 164529
rect 244278 164455 244334 164464
rect 244292 145858 244320 164455
rect 244370 164248 244426 164257
rect 244370 164183 244426 164192
rect 245658 164248 245714 164257
rect 245658 164183 245714 164192
rect 244280 145852 244332 145858
rect 244280 145794 244332 145800
rect 244384 145722 244412 164183
rect 244372 145716 244424 145722
rect 244372 145658 244424 145664
rect 242900 145648 242952 145654
rect 242900 145590 242952 145596
rect 245672 145586 245700 164183
rect 247052 145790 247080 165543
rect 247696 164898 247724 165543
rect 249812 164966 249840 165543
rect 252572 165034 252600 165543
rect 258092 165102 258120 165543
rect 258080 165096 258132 165102
rect 258080 165038 258132 165044
rect 252560 165028 252612 165034
rect 252560 164970 252612 164976
rect 249800 164960 249852 164966
rect 249800 164902 249852 164908
rect 247684 164892 247736 164898
rect 247684 164834 247736 164840
rect 251270 164520 251326 164529
rect 251270 164455 251326 164464
rect 259550 164520 259606 164529
rect 259550 164455 259606 164464
rect 248418 164248 248474 164257
rect 248418 164183 248474 164192
rect 249798 164248 249854 164257
rect 249798 164183 249854 164192
rect 251178 164248 251234 164257
rect 251178 164183 251234 164192
rect 248432 145926 248460 164183
rect 249812 145994 249840 164183
rect 251192 146130 251220 164183
rect 251180 146124 251232 146130
rect 251180 146066 251232 146072
rect 251284 146062 251312 164455
rect 252558 164248 252614 164257
rect 252558 164183 252614 164192
rect 253938 164248 253994 164257
rect 253938 164183 253994 164192
rect 255318 164248 255374 164257
rect 255318 164183 255374 164192
rect 256698 164248 256754 164257
rect 256698 164183 256754 164192
rect 258078 164248 258134 164257
rect 258078 164183 258134 164192
rect 259458 164248 259514 164257
rect 259458 164183 259514 164192
rect 251272 146056 251324 146062
rect 251272 145998 251324 146004
rect 249800 145988 249852 145994
rect 249800 145930 249852 145936
rect 248420 145920 248472 145926
rect 248420 145862 248472 145868
rect 247040 145784 247092 145790
rect 247040 145726 247092 145732
rect 245660 145580 245712 145586
rect 245660 145522 245712 145528
rect 236092 145512 236144 145518
rect 236092 145454 236144 145460
rect 236000 145444 236052 145450
rect 236000 145386 236052 145392
rect 252572 145314 252600 164183
rect 253952 145382 253980 164183
rect 255332 146266 255360 164183
rect 255320 146260 255372 146266
rect 255320 146202 255372 146208
rect 256712 146198 256740 164183
rect 258092 162654 258120 164183
rect 259472 162722 259500 164183
rect 259564 162790 259592 164455
rect 260852 162858 260880 165543
rect 263506 164248 263562 164257
rect 263782 164248 263838 164257
rect 263562 164206 263640 164234
rect 263506 164183 263562 164192
rect 260840 162852 260892 162858
rect 260840 162794 260892 162800
rect 259552 162784 259604 162790
rect 259552 162726 259604 162732
rect 259460 162716 259512 162722
rect 259460 162658 259512 162664
rect 258080 162648 258132 162654
rect 258080 162590 258132 162596
rect 256700 146192 256752 146198
rect 263612 146169 263640 164206
rect 263782 164183 263838 164192
rect 263796 163538 263824 164183
rect 264992 164150 265020 165543
rect 266358 164520 266414 164529
rect 266358 164455 266414 164464
rect 264980 164144 265032 164150
rect 264980 164086 265032 164092
rect 263784 163532 263836 163538
rect 263784 163474 263836 163480
rect 266372 162178 266400 164455
rect 267738 164248 267794 164257
rect 267738 164183 267794 164192
rect 266360 162172 266412 162178
rect 266360 162114 266412 162120
rect 256700 146134 256752 146140
rect 263598 146160 263654 146169
rect 263598 146095 263654 146104
rect 267752 145761 267780 164183
rect 267844 146305 267872 165566
rect 267922 165543 267978 165552
rect 280158 165608 280214 165617
rect 280158 165543 280214 165552
rect 283378 165608 283434 165617
rect 283378 165543 283434 165552
rect 300858 165608 300914 165617
rect 300858 165543 300914 165552
rect 308402 165608 308458 165617
rect 308402 165543 308458 165552
rect 323030 165608 323086 165617
rect 323030 165543 323086 165552
rect 325882 165608 325938 165617
rect 325882 165543 325884 165552
rect 267936 165238 267964 165543
rect 280172 165374 280200 165543
rect 280160 165368 280212 165374
rect 280160 165310 280212 165316
rect 283392 165306 283420 165543
rect 300872 165442 300900 165543
rect 308416 165510 308444 165543
rect 308404 165504 308456 165510
rect 308404 165446 308456 165452
rect 300860 165436 300912 165442
rect 300860 165378 300912 165384
rect 283380 165300 283432 165306
rect 283380 165242 283432 165248
rect 267924 165232 267976 165238
rect 267924 165174 267976 165180
rect 271878 165200 271934 165209
rect 271878 165135 271934 165144
rect 275926 165200 275982 165209
rect 277398 165200 277454 165209
rect 275982 165158 276152 165186
rect 275926 165135 275982 165144
rect 269118 164248 269174 164257
rect 269118 164183 269174 164192
rect 270498 164248 270554 164257
rect 270498 164183 270554 164192
rect 267830 146296 267886 146305
rect 267830 146231 267886 146240
rect 267738 145752 267794 145761
rect 267738 145687 267794 145696
rect 269132 145625 269160 164183
rect 270512 148578 270540 164183
rect 270500 148572 270552 148578
rect 270500 148514 270552 148520
rect 271892 148510 271920 165135
rect 274454 164520 274510 164529
rect 274454 164455 274510 164464
rect 274468 164098 274496 164455
rect 274546 164248 274602 164257
rect 276018 164248 276074 164257
rect 274602 164206 274772 164234
rect 274546 164183 274602 164192
rect 274468 164070 274680 164098
rect 271880 148504 271932 148510
rect 271880 148446 271932 148452
rect 274652 148442 274680 164070
rect 274640 148436 274692 148442
rect 274640 148378 274692 148384
rect 274744 148374 274772 164206
rect 276018 164183 276074 164192
rect 274732 148368 274784 148374
rect 274732 148310 274784 148316
rect 276032 146441 276060 164183
rect 276124 148986 276152 165158
rect 277398 165135 277400 165144
rect 277452 165135 277454 165144
rect 280066 165200 280122 165209
rect 280066 165135 280122 165144
rect 277400 165106 277452 165112
rect 278686 164248 278742 164257
rect 278742 164206 278820 164234
rect 278686 164183 278742 164192
rect 278792 149054 278820 164206
rect 278780 149048 278832 149054
rect 278780 148990 278832 148996
rect 276112 148980 276164 148986
rect 276112 148922 276164 148928
rect 276018 146432 276074 146441
rect 276018 146367 276074 146376
rect 276032 146266 276060 146367
rect 276020 146260 276072 146266
rect 276020 146202 276072 146208
rect 269118 145616 269174 145625
rect 280080 145586 280108 165135
rect 323044 164218 323072 165543
rect 325936 165543 325938 165552
rect 343270 165608 343326 165617
rect 343270 165543 343272 165552
rect 325884 165514 325936 165520
rect 343324 165543 343326 165552
rect 343454 165608 343510 165617
rect 343454 165543 343510 165552
rect 343272 165514 343324 165520
rect 343468 164898 343496 165543
rect 343456 164892 343508 164898
rect 343456 164834 343508 164840
rect 323032 164212 323084 164218
rect 323032 164154 323084 164160
rect 338488 146192 338540 146198
rect 338488 146134 338540 146140
rect 269118 145551 269174 145560
rect 280068 145580 280120 145586
rect 280068 145522 280120 145528
rect 307668 145580 307720 145586
rect 307668 145522 307720 145528
rect 253940 145376 253992 145382
rect 253940 145318 253992 145324
rect 252560 145308 252612 145314
rect 252560 145250 252612 145256
rect 307680 144906 307708 145522
rect 338500 144945 338528 146134
rect 340236 146124 340288 146130
rect 340236 146066 340288 146072
rect 340248 144945 340276 146066
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 307668 144900 307720 144906
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 356624 144906 356652 270438
rect 351642 144871 351698 144880
rect 356612 144900 356664 144906
rect 307668 144842 307720 144848
rect 356612 144842 356664 144848
rect 220084 143336 220136 143342
rect 220084 143278 220136 143284
rect 237102 59800 237158 59809
rect 237102 59735 237158 59744
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 256974 59800 257030 59809
rect 256974 59735 257030 59744
rect 262862 59800 262918 59809
rect 262862 59735 262918 59744
rect 263874 59800 263930 59809
rect 263874 59735 263930 59744
rect 237116 59702 237144 59735
rect 237104 59696 237156 59702
rect 237104 59638 237156 59644
rect 255884 59634 255912 59735
rect 255872 59628 255924 59634
rect 255872 59570 255924 59576
rect 256988 59566 257016 59735
rect 258078 59664 258134 59673
rect 258078 59599 258134 59608
rect 260654 59664 260710 59673
rect 260654 59599 260710 59608
rect 261758 59664 261814 59673
rect 261758 59599 261814 59608
rect 256976 59560 257028 59566
rect 256976 59502 257028 59508
rect 258092 59294 258120 59599
rect 258080 59288 258132 59294
rect 258080 59230 258132 59236
rect 260668 59226 260696 59599
rect 260656 59220 260708 59226
rect 260656 59162 260708 59168
rect 261772 59158 261800 59599
rect 262876 59430 262904 59735
rect 263888 59498 263916 59735
rect 308494 59664 308550 59673
rect 308494 59599 308550 59608
rect 315854 59664 315910 59673
rect 315854 59599 315910 59608
rect 263876 59492 263928 59498
rect 263876 59434 263928 59440
rect 262864 59424 262916 59430
rect 262864 59366 262916 59372
rect 279238 59256 279294 59265
rect 279238 59191 279294 59200
rect 290922 59256 290978 59265
rect 290922 59191 290978 59200
rect 300858 59256 300914 59265
rect 300858 59191 300914 59200
rect 279252 59158 279280 59191
rect 261760 59152 261812 59158
rect 261760 59094 261812 59100
rect 279240 59152 279292 59158
rect 279240 59094 279292 59100
rect 290936 59090 290964 59191
rect 290924 59084 290976 59090
rect 290924 59026 290976 59032
rect 300872 59022 300900 59191
rect 300860 59016 300912 59022
rect 300860 58958 300912 58964
rect 308508 58886 308536 59599
rect 315868 58954 315896 59599
rect 320914 59256 320970 59265
rect 320914 59191 320970 59200
rect 325882 59256 325938 59265
rect 325882 59191 325938 59200
rect 315856 58948 315908 58954
rect 315856 58890 315908 58896
rect 308496 58880 308548 58886
rect 308496 58822 308548 58828
rect 320928 58818 320956 59191
rect 320916 58812 320968 58818
rect 320916 58754 320968 58760
rect 325896 58750 325924 59191
rect 356624 59158 356652 144842
rect 356612 59152 356664 59158
rect 356612 59094 356664 59100
rect 356716 58886 356744 485250
rect 356808 166802 356836 485522
rect 358268 485512 358320 485518
rect 358268 485454 358320 485460
rect 358176 485240 358228 485246
rect 358176 485182 358228 485188
rect 358084 484356 358136 484362
rect 358084 484298 358136 484304
rect 356888 479800 356940 479806
rect 356888 479742 356940 479748
rect 356900 272882 356928 479742
rect 357072 478508 357124 478514
rect 357072 478450 357124 478456
rect 356980 466540 357032 466546
rect 356980 466482 357032 466488
rect 356992 359582 357020 466482
rect 357084 377670 357112 478450
rect 357256 474700 357308 474706
rect 357256 474642 357308 474648
rect 357164 471980 357216 471986
rect 357164 471922 357216 471928
rect 357072 377664 357124 377670
rect 357072 377606 357124 377612
rect 357072 375420 357124 375426
rect 357072 375362 357124 375368
rect 356980 359576 357032 359582
rect 356980 359518 357032 359524
rect 356888 272876 356940 272882
rect 356888 272818 356940 272824
rect 356980 271924 357032 271930
rect 356980 271866 357032 271872
rect 356992 271250 357020 271866
rect 356980 271244 357032 271250
rect 356980 271186 357032 271192
rect 356888 271176 356940 271182
rect 356888 271118 356940 271124
rect 356796 166796 356848 166802
rect 356796 166738 356848 166744
rect 356900 146266 356928 271118
rect 356992 165578 357020 271186
rect 357084 270502 357112 375362
rect 357176 374814 357204 471922
rect 357268 378078 357296 474642
rect 357992 470144 358044 470150
rect 357992 470086 358044 470092
rect 357808 469804 357860 469810
rect 357808 469746 357860 469752
rect 357820 411942 357848 469746
rect 357900 465656 357952 465662
rect 357900 465598 357952 465604
rect 357808 411936 357860 411942
rect 357808 411878 357860 411884
rect 357912 378962 357940 465598
rect 357900 378956 357952 378962
rect 357900 378898 357952 378904
rect 357256 378072 357308 378078
rect 357256 378014 357308 378020
rect 358004 377602 358032 470086
rect 358096 417450 358124 484298
rect 358084 417444 358136 417450
rect 358084 417386 358136 417392
rect 358084 389224 358136 389230
rect 358084 389166 358136 389172
rect 357992 377596 358044 377602
rect 357992 377538 358044 377544
rect 357164 374808 357216 374814
rect 357164 374750 357216 374756
rect 357164 359576 357216 359582
rect 357164 359518 357216 359524
rect 357072 270496 357124 270502
rect 357072 270438 357124 270444
rect 357176 253978 357204 359518
rect 358096 359514 358124 389166
rect 358084 359508 358136 359514
rect 358084 359450 358136 359456
rect 358096 282198 358124 359450
rect 358084 282192 358136 282198
rect 358084 282134 358136 282140
rect 357164 253972 357216 253978
rect 357164 253914 357216 253920
rect 357532 253972 357584 253978
rect 357532 253914 357584 253920
rect 356980 165572 357032 165578
rect 356980 165514 357032 165520
rect 357440 165572 357492 165578
rect 357440 165514 357492 165520
rect 356888 146260 356940 146266
rect 356888 146202 356940 146208
rect 356704 58880 356756 58886
rect 356704 58822 356756 58828
rect 325884 58744 325936 58750
rect 325884 58686 325936 58692
rect 323308 57928 323360 57934
rect 235998 57896 236054 57905
rect 235998 57831 236054 57840
rect 237378 57896 237434 57905
rect 237378 57831 237434 57840
rect 239126 57896 239182 57905
rect 239126 57831 239182 57840
rect 240138 57896 240194 57905
rect 240138 57831 240194 57840
rect 241610 57896 241666 57905
rect 241610 57831 241666 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 245290 57896 245346 57905
rect 245290 57831 245346 57840
rect 245658 57896 245714 57905
rect 245658 57831 245714 57840
rect 247038 57896 247094 57905
rect 247038 57831 247094 57840
rect 248602 57896 248658 57905
rect 248602 57831 248658 57840
rect 249798 57896 249854 57905
rect 249798 57831 249854 57840
rect 251178 57896 251234 57905
rect 251178 57831 251234 57840
rect 251362 57896 251418 57905
rect 251362 57831 251418 57840
rect 253386 57896 253442 57905
rect 253386 57831 253442 57840
rect 253938 57896 253994 57905
rect 253938 57831 253994 57840
rect 258354 57896 258410 57905
rect 258354 57831 258410 57840
rect 264978 57896 265034 57905
rect 264978 57831 265034 57840
rect 266358 57896 266414 57905
rect 266358 57831 266414 57840
rect 268474 57896 268530 57905
rect 268474 57831 268530 57840
rect 271050 57896 271106 57905
rect 271050 57831 271106 57840
rect 271878 57896 271934 57905
rect 271878 57831 271934 57840
rect 273258 57896 273314 57905
rect 273258 57831 273314 57840
rect 275098 57896 275154 57905
rect 275098 57831 275154 57840
rect 283470 57896 283526 57905
rect 283470 57831 283526 57840
rect 293314 57896 293370 57905
rect 293314 57831 293370 57840
rect 295890 57896 295946 57905
rect 295890 57831 295946 57840
rect 298098 57896 298154 57905
rect 298098 57831 298154 57840
rect 303434 57896 303490 57905
rect 303434 57831 303490 57840
rect 305826 57896 305882 57905
rect 305826 57831 305882 57840
rect 310978 57896 311034 57905
rect 310978 57831 310980 57840
rect 236012 56506 236040 57831
rect 236000 56500 236052 56506
rect 236000 56442 236052 56448
rect 219992 55820 220044 55826
rect 219992 55762 220044 55768
rect 219716 54868 219768 54874
rect 219716 54810 219768 54816
rect 218796 54528 218848 54534
rect 218796 54470 218848 54476
rect 216036 54460 216088 54466
rect 216036 54402 216088 54408
rect 237392 54398 237420 57831
rect 239140 55894 239168 57831
rect 239128 55888 239180 55894
rect 239128 55830 239180 55836
rect 237380 54392 237432 54398
rect 237380 54334 237432 54340
rect 240152 54330 240180 57831
rect 241624 56574 241652 57831
rect 241612 56568 241664 56574
rect 241612 56510 241664 56516
rect 242912 54466 242940 57831
rect 244384 54602 244412 57831
rect 245304 55962 245332 57831
rect 245292 55956 245344 55962
rect 245292 55898 245344 55904
rect 244372 54596 244424 54602
rect 244372 54538 244424 54544
rect 245672 54534 245700 57831
rect 247052 54670 247080 57831
rect 248616 56030 248644 57831
rect 248604 56024 248656 56030
rect 248604 55966 248656 55972
rect 249812 54738 249840 57831
rect 251192 56098 251220 57831
rect 251180 56092 251232 56098
rect 251180 56034 251232 56040
rect 251376 54806 251404 57831
rect 253400 56166 253428 57831
rect 253388 56160 253440 56166
rect 253388 56102 253440 56108
rect 253952 54874 253980 57831
rect 258368 57254 258396 57831
rect 258356 57248 258408 57254
rect 258356 57190 258408 57196
rect 264992 54942 265020 57831
rect 266372 56234 266400 57831
rect 266450 57624 266506 57633
rect 266450 57559 266506 57568
rect 266360 56228 266412 56234
rect 266360 56170 266412 56176
rect 266464 55010 266492 57559
rect 268488 56302 268516 57831
rect 269118 57624 269174 57633
rect 269118 57559 269174 57568
rect 268476 56296 268528 56302
rect 268476 56238 268528 56244
rect 269132 55185 269160 57559
rect 271064 56370 271092 57831
rect 271052 56364 271104 56370
rect 271052 56306 271104 56312
rect 269118 55176 269174 55185
rect 269118 55111 269174 55120
rect 271892 55078 271920 57831
rect 273272 56438 273300 57831
rect 273350 57624 273406 57633
rect 273350 57559 273406 57568
rect 273260 56432 273312 56438
rect 273260 56374 273312 56380
rect 273364 55146 273392 57559
rect 275112 55758 275140 57831
rect 277398 57624 277454 57633
rect 277398 57559 277454 57568
rect 275100 55752 275152 55758
rect 275100 55694 275152 55700
rect 277412 55214 277440 57559
rect 283484 57322 283512 57831
rect 293328 57458 293356 57831
rect 295904 57662 295932 57831
rect 295892 57656 295944 57662
rect 295892 57598 295944 57604
rect 293316 57452 293368 57458
rect 293316 57394 293368 57400
rect 298112 57390 298140 57831
rect 303448 57594 303476 57831
rect 303436 57588 303488 57594
rect 303436 57530 303488 57536
rect 305840 57526 305868 57831
rect 311032 57831 311034 57840
rect 313370 57896 313426 57905
rect 313370 57831 313426 57840
rect 318338 57896 318394 57905
rect 318338 57831 318394 57840
rect 323306 57896 323308 57905
rect 343456 57928 343508 57934
rect 323360 57896 323362 57905
rect 323306 57831 323362 57840
rect 343178 57896 343234 57905
rect 343178 57831 343180 57840
rect 310980 57802 311032 57808
rect 313384 57798 313412 57831
rect 313372 57792 313424 57798
rect 313372 57734 313424 57740
rect 318352 57730 318380 57831
rect 343232 57831 343234 57840
rect 343454 57896 343456 57905
rect 343508 57896 343510 57905
rect 357452 57866 357480 165514
rect 357544 156670 357572 253914
rect 358096 253230 358124 282134
rect 358084 253224 358136 253230
rect 358084 253166 358136 253172
rect 358096 175982 358124 253166
rect 358084 175976 358136 175982
rect 358084 175918 358136 175924
rect 357624 165640 357676 165646
rect 357624 165582 357676 165588
rect 357636 164898 357664 165582
rect 357624 164892 357676 164898
rect 357624 164834 357676 164840
rect 357532 156664 357584 156670
rect 357532 156606 357584 156612
rect 357636 57934 357664 164834
rect 357716 156664 357768 156670
rect 357716 156606 357768 156612
rect 357728 146130 357756 156606
rect 357716 146124 357768 146130
rect 357716 146066 357768 146072
rect 358096 145586 358124 175918
rect 358084 145580 358136 145586
rect 358084 145522 358136 145528
rect 358084 68468 358136 68474
rect 358084 68410 358136 68416
rect 358096 59362 358124 68410
rect 358188 59430 358216 485182
rect 358280 166938 358308 485454
rect 358360 485444 358412 485450
rect 358360 485386 358412 485392
rect 358268 166932 358320 166938
rect 358268 166874 358320 166880
rect 358372 166870 358400 485386
rect 364984 485376 365036 485382
rect 364984 485318 365036 485324
rect 362224 485104 362276 485110
rect 362224 485046 362276 485052
rect 359832 482724 359884 482730
rect 359832 482666 359884 482672
rect 359464 478440 359516 478446
rect 359464 478382 359516 478388
rect 358544 469124 358596 469130
rect 358544 469066 358596 469072
rect 358452 468852 358504 468858
rect 358452 468794 358504 468800
rect 358464 272950 358492 468794
rect 358556 376310 358584 469066
rect 358728 467764 358780 467770
rect 358728 467706 358780 467712
rect 358634 417480 358690 417489
rect 358634 417415 358690 417424
rect 358544 376304 358596 376310
rect 358544 376246 358596 376252
rect 358544 358896 358596 358902
rect 358544 358838 358596 358844
rect 358452 272944 358504 272950
rect 358452 272886 358504 272892
rect 358556 271862 358584 358838
rect 358544 271856 358596 271862
rect 358544 271798 358596 271804
rect 358360 166864 358412 166870
rect 358360 166806 358412 166812
rect 358176 59424 358228 59430
rect 358176 59366 358228 59372
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 358648 57934 358676 417415
rect 358740 374882 358768 467706
rect 358820 465112 358872 465118
rect 358820 465054 358872 465060
rect 358832 460193 358860 465054
rect 358818 460184 358874 460193
rect 358818 460119 358874 460128
rect 358728 374876 358780 374882
rect 358728 374818 358780 374824
rect 358832 354674 358860 460119
rect 359094 398168 359150 398177
rect 359094 398103 359150 398112
rect 359002 396808 359058 396817
rect 359002 396743 359058 396752
rect 358910 394088 358966 394097
rect 358910 394023 358966 394032
rect 358924 362234 358952 394023
rect 359016 366382 359044 396743
rect 359108 370530 359136 398103
rect 359186 395312 359242 395321
rect 359186 395247 359242 395256
rect 359200 371890 359228 395247
rect 359476 380526 359504 478382
rect 359556 471912 359608 471918
rect 359556 471854 359608 471860
rect 359464 380520 359516 380526
rect 359464 380462 359516 380468
rect 359568 378826 359596 471854
rect 359740 470348 359792 470354
rect 359740 470290 359792 470296
rect 359648 468988 359700 468994
rect 359648 468930 359700 468936
rect 359660 389162 359688 468930
rect 359752 391950 359780 470290
rect 359844 414730 359872 482666
rect 361304 482656 361356 482662
rect 361304 482598 361356 482604
rect 360936 482316 360988 482322
rect 360936 482258 360988 482264
rect 360844 481024 360896 481030
rect 360844 480966 360896 480972
rect 359924 470484 359976 470490
rect 359924 470426 359976 470432
rect 359832 414724 359884 414730
rect 359832 414666 359884 414672
rect 359936 409154 359964 470426
rect 360016 470416 360068 470422
rect 360016 470358 360068 470364
rect 360028 410582 360056 470358
rect 360200 466472 360252 466478
rect 360200 466414 360252 466420
rect 360016 410576 360068 410582
rect 360016 410518 360068 410524
rect 359924 409148 359976 409154
rect 359924 409090 359976 409096
rect 359830 400344 359886 400353
rect 359830 400279 359886 400288
rect 359740 391944 359792 391950
rect 359740 391886 359792 391892
rect 359648 389156 359700 389162
rect 359648 389098 359700 389104
rect 359556 378820 359608 378826
rect 359556 378762 359608 378768
rect 359372 378344 359424 378350
rect 359372 378286 359424 378292
rect 359188 371884 359240 371890
rect 359188 371826 359240 371832
rect 359200 371278 359228 371826
rect 359188 371272 359240 371278
rect 359188 371214 359240 371220
rect 359096 370524 359148 370530
rect 359096 370466 359148 370472
rect 359108 369322 359136 370466
rect 359108 369294 359228 369322
rect 359096 369164 359148 369170
rect 359096 369106 359148 369112
rect 359004 366376 359056 366382
rect 359004 366318 359056 366324
rect 358912 362228 358964 362234
rect 358912 362170 358964 362176
rect 358832 354646 358952 354674
rect 358924 353161 358952 354646
rect 358910 353152 358966 353161
rect 358910 353087 358966 353096
rect 358818 289776 358874 289785
rect 358818 289711 358874 289720
rect 358832 288833 358860 289711
rect 358818 288824 358874 288833
rect 358818 288759 358874 288768
rect 358832 182073 358860 288759
rect 358924 246265 358952 353087
rect 359016 291009 359044 366318
rect 359108 292777 359136 369106
rect 359200 365022 359228 369294
rect 359188 365016 359240 365022
rect 359188 364958 359240 364964
rect 359188 362228 359240 362234
rect 359188 362170 359240 362176
rect 359094 292768 359150 292777
rect 359094 292703 359150 292712
rect 359094 291816 359150 291825
rect 359094 291751 359150 291760
rect 359002 291000 359058 291009
rect 359002 290935 359058 290944
rect 359002 288416 359058 288425
rect 359002 288351 359058 288360
rect 359016 287609 359044 288351
rect 359002 287600 359058 287609
rect 359002 287535 359058 287544
rect 358910 246256 358966 246265
rect 358910 246191 358966 246200
rect 358818 182064 358874 182073
rect 358818 181999 358874 182008
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68474 358768 145522
rect 358924 139369 358952 246191
rect 359016 180713 359044 287535
rect 359108 184929 359136 291751
rect 359200 288425 359228 362170
rect 359278 292768 359334 292777
rect 359278 292703 359334 292712
rect 359186 288416 359242 288425
rect 359186 288351 359242 288360
rect 359292 190454 359320 292703
rect 359384 271930 359412 378286
rect 359464 371272 359516 371278
rect 359464 371214 359516 371220
rect 359476 363662 359504 371214
rect 359844 370530 359872 400279
rect 360212 390522 360240 466414
rect 360752 465588 360804 465594
rect 360752 465530 360804 465536
rect 360200 390516 360252 390522
rect 360200 390458 360252 390464
rect 360212 389230 360240 390458
rect 360200 389224 360252 389230
rect 360200 389166 360252 389172
rect 360764 380662 360792 465530
rect 360752 380656 360804 380662
rect 360752 380598 360804 380604
rect 359832 370524 359884 370530
rect 359832 370466 359884 370472
rect 359844 369170 359872 370466
rect 359832 369164 359884 369170
rect 359832 369106 359884 369112
rect 359556 365016 359608 365022
rect 359556 364958 359608 364964
rect 359464 363656 359516 363662
rect 359464 363598 359516 363604
rect 359476 289785 359504 363598
rect 359568 291825 359596 364958
rect 360200 359304 360252 359310
rect 360200 359246 360252 359252
rect 360212 358834 360240 359246
rect 360200 358828 360252 358834
rect 360200 358770 360252 358776
rect 359554 291816 359610 291825
rect 359554 291751 359610 291760
rect 359554 291000 359610 291009
rect 359554 290935 359610 290944
rect 359462 289776 359518 289785
rect 359462 289711 359518 289720
rect 359372 271924 359424 271930
rect 359372 271866 359424 271872
rect 359292 190426 359412 190454
rect 359384 186425 359412 190426
rect 359370 186416 359426 186425
rect 359370 186351 359426 186360
rect 359094 184920 359150 184929
rect 359094 184855 359150 184864
rect 359002 180704 359058 180713
rect 359002 180639 359058 180648
rect 358910 139360 358966 139369
rect 358910 139295 358966 139304
rect 359016 74089 359044 180639
rect 359108 78305 359136 184855
rect 359278 183560 359334 183569
rect 359278 183495 359334 183504
rect 359186 182064 359242 182073
rect 359186 181999 359242 182008
rect 359094 78296 359150 78305
rect 359094 78231 359150 78240
rect 359200 75449 359228 181999
rect 359292 76945 359320 183495
rect 359384 79937 359412 186351
rect 359568 183569 359596 290935
rect 360212 253298 360240 358770
rect 360292 271924 360344 271930
rect 360292 271866 360344 271872
rect 360200 253292 360252 253298
rect 360200 253234 360252 253240
rect 359554 183560 359610 183569
rect 359554 183495 359610 183504
rect 360212 146198 360240 253234
rect 360304 165646 360332 271866
rect 360292 165640 360344 165646
rect 360292 165582 360344 165588
rect 360200 146192 360252 146198
rect 360200 146134 360252 146140
rect 359370 79928 359426 79937
rect 359370 79863 359426 79872
rect 359278 76936 359334 76945
rect 359278 76871 359334 76880
rect 359186 75440 359242 75449
rect 359186 75375 359242 75384
rect 359002 74080 359058 74089
rect 359002 74015 359058 74024
rect 358728 68468 358780 68474
rect 358728 68410 358780 68416
rect 357624 57928 357676 57934
rect 357624 57870 357676 57876
rect 358636 57928 358688 57934
rect 358636 57870 358688 57876
rect 343454 57831 343510 57840
rect 357440 57860 357492 57866
rect 343180 57802 343232 57808
rect 357440 57802 357492 57808
rect 360856 57730 360884 480966
rect 360948 165510 360976 482258
rect 361028 479732 361080 479738
rect 361028 479674 361080 479680
rect 361040 271454 361068 479674
rect 361120 469872 361172 469878
rect 361120 469814 361172 469820
rect 361132 273057 361160 469814
rect 361212 468920 361264 468926
rect 361212 468862 361264 468868
rect 361224 284306 361252 468862
rect 361316 377942 361344 482598
rect 361396 480004 361448 480010
rect 361396 479946 361448 479952
rect 361304 377936 361356 377942
rect 361304 377878 361356 377884
rect 361408 376718 361436 479946
rect 361488 473204 361540 473210
rect 361488 473146 361540 473152
rect 361500 377534 361528 473146
rect 362132 467628 362184 467634
rect 362132 467570 362184 467576
rect 362144 377806 362172 467570
rect 362132 377800 362184 377806
rect 362132 377742 362184 377748
rect 361488 377528 361540 377534
rect 361488 377470 361540 377476
rect 361396 376712 361448 376718
rect 361396 376654 361448 376660
rect 361212 284300 361264 284306
rect 361212 284242 361264 284248
rect 361118 273048 361174 273057
rect 361118 272983 361174 272992
rect 361028 271448 361080 271454
rect 361028 271390 361080 271396
rect 360936 165504 360988 165510
rect 360936 165446 360988 165452
rect 362236 58954 362264 485046
rect 363972 484084 364024 484090
rect 363972 484026 364024 484032
rect 363604 483812 363656 483818
rect 363604 483754 363656 483760
rect 362592 482452 362644 482458
rect 362592 482394 362644 482400
rect 362408 475380 362460 475386
rect 362408 475322 362460 475328
rect 362316 474020 362368 474026
rect 362316 473962 362368 473968
rect 362224 58948 362276 58954
rect 362224 58890 362276 58896
rect 318340 57724 318392 57730
rect 318340 57666 318392 57672
rect 360844 57724 360896 57730
rect 360844 57666 360896 57672
rect 362328 57594 362356 473962
rect 362420 165578 362448 475322
rect 362500 473068 362552 473074
rect 362500 473010 362552 473016
rect 362512 167006 362540 473010
rect 362604 271318 362632 482394
rect 362776 477488 362828 477494
rect 362776 477430 362828 477436
rect 362684 467492 362736 467498
rect 362684 467434 362736 467440
rect 362696 273358 362724 467434
rect 362788 374950 362816 477430
rect 363512 475652 363564 475658
rect 363512 475594 363564 475600
rect 362868 467696 362920 467702
rect 362868 467638 362920 467644
rect 362880 376582 362908 467638
rect 362960 466608 363012 466614
rect 362960 466550 363012 466556
rect 362972 466478 363000 466550
rect 362960 466472 363012 466478
rect 362960 466414 363012 466420
rect 362868 376576 362920 376582
rect 362868 376518 362920 376524
rect 362776 374944 362828 374950
rect 362776 374886 362828 374892
rect 362972 359310 363000 466414
rect 363524 377466 363552 475594
rect 363512 377460 363564 377466
rect 363512 377402 363564 377408
rect 362960 359304 363012 359310
rect 362960 359246 363012 359252
rect 362684 273352 362736 273358
rect 362684 273294 362736 273300
rect 362592 271312 362644 271318
rect 362592 271254 362644 271260
rect 362500 167000 362552 167006
rect 362500 166942 362552 166948
rect 362408 165572 362460 165578
rect 362408 165514 362460 165520
rect 363616 57662 363644 483754
rect 363788 479528 363840 479534
rect 363788 479470 363840 479476
rect 363696 474088 363748 474094
rect 363696 474030 363748 474036
rect 363708 57798 363736 474030
rect 363800 70378 363828 479470
rect 363880 467288 363932 467294
rect 363880 467230 363932 467236
rect 363892 178022 363920 467230
rect 363984 271522 364012 484026
rect 364156 477352 364208 477358
rect 364156 477294 364208 477300
rect 364064 474564 364116 474570
rect 364064 474506 364116 474512
rect 364076 272678 364104 474506
rect 364168 377262 364196 477294
rect 364248 477284 364300 477290
rect 364248 477226 364300 477232
rect 364260 377874 364288 477226
rect 364892 469056 364944 469062
rect 364892 468998 364944 469004
rect 364800 464500 364852 464506
rect 364800 464442 364852 464448
rect 364812 380798 364840 464442
rect 364800 380792 364852 380798
rect 364800 380734 364852 380740
rect 364904 380254 364932 468998
rect 364892 380248 364944 380254
rect 364892 380190 364944 380196
rect 364248 377868 364300 377874
rect 364248 377810 364300 377816
rect 364156 377256 364208 377262
rect 364156 377198 364208 377204
rect 364064 272672 364116 272678
rect 364064 272614 364116 272620
rect 363972 271516 364024 271522
rect 363972 271458 364024 271464
rect 363880 178016 363932 178022
rect 363880 177958 363932 177964
rect 363788 70372 363840 70378
rect 363788 70314 363840 70320
rect 364996 58750 365024 485318
rect 366364 485172 366416 485178
rect 366364 485114 366416 485120
rect 365076 481092 365128 481098
rect 365076 481034 365128 481040
rect 365088 165170 365116 481034
rect 365352 477148 365404 477154
rect 365352 477090 365404 477096
rect 365168 471300 365220 471306
rect 365168 471242 365220 471248
rect 365180 166394 365208 471242
rect 365260 465792 365312 465798
rect 365260 465734 365312 465740
rect 365272 175234 365300 465734
rect 365364 271658 365392 477090
rect 365444 477080 365496 477086
rect 365444 477022 365496 477028
rect 365456 273086 365484 477022
rect 365536 473884 365588 473890
rect 365536 473826 365588 473832
rect 365548 376038 365576 473826
rect 366272 470552 366324 470558
rect 366272 470494 366324 470500
rect 365628 469192 365680 469198
rect 365628 469134 365680 469140
rect 365640 380186 365668 469134
rect 366180 466404 366232 466410
rect 366180 466346 366232 466352
rect 365628 380180 365680 380186
rect 365628 380122 365680 380128
rect 366192 378010 366220 466346
rect 366284 380050 366312 470494
rect 366272 380044 366324 380050
rect 366272 379986 366324 379992
rect 366180 378004 366232 378010
rect 366180 377946 366232 377952
rect 365536 376032 365588 376038
rect 365536 375974 365588 375980
rect 365444 273080 365496 273086
rect 365444 273022 365496 273028
rect 365352 271652 365404 271658
rect 365352 271594 365404 271600
rect 365260 175228 365312 175234
rect 365260 175170 365312 175176
rect 365168 166388 365220 166394
rect 365168 166330 365220 166336
rect 365076 165164 365128 165170
rect 365076 165106 365128 165112
rect 366376 58818 366404 485114
rect 371148 484288 371200 484294
rect 371148 484230 371200 484236
rect 366916 484220 366968 484226
rect 366916 484162 366968 484168
rect 366732 481160 366784 481166
rect 366732 481102 366784 481108
rect 366640 474428 366692 474434
rect 366640 474370 366692 474376
rect 366548 474360 366600 474366
rect 366548 474302 366600 474308
rect 366456 474224 366508 474230
rect 366456 474166 366508 474172
rect 366468 165238 366496 474166
rect 366456 165232 366508 165238
rect 366456 165174 366508 165180
rect 366560 164665 366588 474302
rect 366652 166326 366680 474370
rect 366744 271862 366772 481102
rect 366824 477216 366876 477222
rect 366824 477158 366876 477164
rect 366836 272610 366864 477158
rect 366928 376650 366956 484162
rect 369124 483948 369176 483954
rect 369124 483890 369176 483896
rect 368296 482520 368348 482526
rect 368296 482462 368348 482468
rect 367836 476944 367888 476950
rect 367836 476886 367888 476892
rect 367560 474632 367612 474638
rect 367560 474574 367612 474580
rect 367008 470212 367060 470218
rect 367008 470154 367060 470160
rect 367020 378146 367048 470154
rect 367572 380390 367600 474574
rect 367652 473272 367704 473278
rect 367652 473214 367704 473220
rect 367560 380384 367612 380390
rect 367560 380326 367612 380332
rect 367008 378140 367060 378146
rect 367008 378082 367060 378088
rect 366916 376644 366968 376650
rect 366916 376586 366968 376592
rect 367664 375222 367692 473214
rect 367744 472864 367796 472870
rect 367744 472806 367796 472812
rect 367652 375216 367704 375222
rect 367652 375158 367704 375164
rect 366824 272604 366876 272610
rect 366824 272546 366876 272552
rect 366732 271856 366784 271862
rect 366732 271798 366784 271804
rect 366640 166320 366692 166326
rect 366640 166262 366692 166268
rect 366546 164656 366602 164665
rect 366546 164591 366602 164600
rect 366364 58812 366416 58818
rect 366364 58754 366416 58760
rect 364984 58744 365036 58750
rect 364984 58686 365036 58692
rect 363696 57792 363748 57798
rect 363696 57734 363748 57740
rect 363604 57656 363656 57662
rect 363604 57598 363656 57604
rect 362316 57588 362368 57594
rect 362316 57530 362368 57536
rect 367756 57526 367784 472806
rect 367848 165034 367876 476886
rect 367928 468648 367980 468654
rect 367928 468590 367980 468596
rect 367940 166462 367968 468590
rect 368020 467356 368072 467362
rect 368020 467298 368072 467304
rect 368032 271386 368060 467298
rect 368204 467220 368256 467226
rect 368204 467162 368256 467168
rect 368112 464364 368164 464370
rect 368112 464306 368164 464312
rect 368124 272542 368152 464306
rect 368216 282878 368244 467162
rect 368308 376378 368336 482462
rect 368388 477420 368440 477426
rect 368388 477362 368440 477368
rect 368296 376372 368348 376378
rect 368296 376314 368348 376320
rect 368400 375018 368428 477362
rect 369032 473952 369084 473958
rect 369032 473894 369084 473900
rect 368940 471844 368992 471850
rect 368940 471786 368992 471792
rect 368848 471232 368900 471238
rect 368848 471174 368900 471180
rect 368860 379506 368888 471174
rect 368848 379500 368900 379506
rect 368848 379442 368900 379448
rect 368952 375358 368980 471786
rect 369044 377330 369072 473894
rect 369032 377324 369084 377330
rect 369032 377266 369084 377272
rect 368940 375352 368992 375358
rect 368940 375294 368992 375300
rect 368388 375012 368440 375018
rect 368388 374954 368440 374960
rect 368204 282872 368256 282878
rect 368204 282814 368256 282820
rect 369032 273420 369084 273426
rect 369032 273362 369084 273368
rect 368112 272536 368164 272542
rect 368112 272478 368164 272484
rect 368020 271380 368072 271386
rect 368020 271322 368072 271328
rect 367928 166456 367980 166462
rect 367928 166398 367980 166404
rect 367836 165028 367888 165034
rect 367836 164970 367888 164976
rect 369044 145625 369072 273362
rect 369136 165306 369164 483890
rect 370504 483744 370556 483750
rect 370504 483686 370556 483692
rect 369584 482588 369636 482594
rect 369584 482530 369636 482536
rect 369400 471368 369452 471374
rect 369400 471310 369452 471316
rect 369308 466132 369360 466138
rect 369308 466074 369360 466080
rect 369216 465860 369268 465866
rect 369216 465802 369268 465808
rect 369124 165300 369176 165306
rect 369124 165242 369176 165248
rect 369228 165102 369256 465802
rect 369320 166734 369348 466074
rect 369412 273290 369440 471310
rect 369492 466268 369544 466274
rect 369492 466210 369544 466216
rect 369400 273284 369452 273290
rect 369400 273226 369452 273232
rect 369504 271726 369532 466210
rect 369596 376446 369624 482530
rect 370412 481296 370464 481302
rect 370412 481238 370464 481244
rect 370320 479868 370372 479874
rect 370320 479810 370372 479816
rect 370228 471776 370280 471782
rect 370228 471718 370280 471724
rect 369676 467560 369728 467566
rect 369676 467502 369728 467508
rect 369688 380322 369716 467502
rect 369676 380316 369728 380322
rect 369676 380258 369728 380264
rect 369674 379128 369730 379137
rect 369674 379063 369730 379072
rect 369584 376440 369636 376446
rect 369584 376382 369636 376388
rect 369584 375352 369636 375358
rect 369584 375294 369636 375300
rect 369492 271720 369544 271726
rect 369492 271662 369544 271668
rect 369596 251870 369624 375294
rect 369688 270434 369716 379063
rect 369766 378992 369822 379001
rect 369766 378927 369822 378936
rect 369780 270502 369808 378927
rect 370044 375216 370096 375222
rect 370044 375158 370096 375164
rect 370056 374542 370084 375158
rect 370240 374678 370268 471718
rect 370332 380458 370360 479810
rect 370424 380905 370452 481238
rect 370410 380896 370466 380905
rect 370410 380831 370466 380840
rect 370320 380452 370372 380458
rect 370320 380394 370372 380400
rect 370228 374672 370280 374678
rect 370228 374614 370280 374620
rect 370044 374536 370096 374542
rect 370044 374478 370096 374484
rect 370412 374536 370464 374542
rect 370412 374478 370464 374484
rect 370320 273488 370372 273494
rect 370320 273430 370372 273436
rect 369768 270496 369820 270502
rect 369768 270438 369820 270444
rect 369676 270428 369728 270434
rect 369676 270370 369728 270376
rect 369584 251864 369636 251870
rect 369584 251806 369636 251812
rect 369308 166728 369360 166734
rect 369308 166670 369360 166676
rect 369216 165096 369268 165102
rect 369216 165038 369268 165044
rect 369688 147626 369716 270370
rect 369676 147620 369728 147626
rect 369676 147562 369728 147568
rect 370332 145761 370360 273430
rect 370424 251938 370452 374478
rect 370412 251932 370464 251938
rect 370412 251874 370464 251880
rect 370318 145752 370374 145761
rect 370318 145687 370374 145696
rect 369030 145616 369086 145625
rect 369030 145551 369086 145560
rect 305828 57520 305880 57526
rect 305828 57462 305880 57468
rect 367744 57520 367796 57526
rect 367744 57462 367796 57468
rect 298100 57384 298152 57390
rect 298100 57326 298152 57332
rect 370516 57322 370544 483686
rect 370872 479664 370924 479670
rect 370872 479606 370924 479612
rect 370596 472660 370648 472666
rect 370596 472602 370648 472608
rect 370608 57390 370636 472602
rect 370780 466064 370832 466070
rect 370780 466006 370832 466012
rect 370688 465928 370740 465934
rect 370688 465870 370740 465876
rect 370700 165374 370728 465870
rect 370792 166598 370820 466006
rect 370884 271250 370912 479606
rect 370964 473136 371016 473142
rect 370964 473078 371016 473084
rect 370976 272814 371004 473078
rect 371056 379704 371108 379710
rect 371056 379646 371108 379652
rect 370964 272808 371016 272814
rect 370964 272750 371016 272756
rect 370872 271244 370924 271250
rect 370872 271186 370924 271192
rect 370964 270224 371016 270230
rect 370964 270166 371016 270172
rect 370780 166592 370832 166598
rect 370780 166534 370832 166540
rect 370688 165368 370740 165374
rect 370688 165310 370740 165316
rect 370976 148510 371004 270166
rect 371068 252006 371096 379646
rect 371160 379030 371188 484230
rect 379980 484152 380032 484158
rect 379980 484094 380032 484100
rect 376208 484016 376260 484022
rect 376208 483958 376260 483964
rect 373540 482384 373592 482390
rect 373540 482326 373592 482332
rect 371700 480072 371752 480078
rect 371700 480014 371752 480020
rect 371608 468784 371660 468790
rect 371608 468726 371660 468732
rect 371148 379024 371200 379030
rect 371148 378966 371200 378972
rect 371148 377528 371200 377534
rect 371148 377470 371200 377476
rect 371160 377398 371188 377470
rect 371148 377392 371200 377398
rect 371148 377334 371200 377340
rect 371160 273222 371188 377334
rect 371148 273216 371200 273222
rect 371148 273158 371200 273164
rect 371620 272921 371648 468726
rect 371712 374746 371740 480014
rect 372436 479936 372488 479942
rect 372436 479878 372488 479884
rect 371976 479596 372028 479602
rect 371976 479538 372028 479544
rect 371884 472728 371936 472734
rect 371884 472670 371936 472676
rect 371792 466336 371844 466342
rect 371792 466278 371844 466284
rect 371804 376106 371832 466278
rect 371792 376100 371844 376106
rect 371792 376042 371844 376048
rect 371700 374740 371752 374746
rect 371700 374682 371752 374688
rect 371790 374640 371846 374649
rect 371790 374575 371846 374584
rect 371606 272912 371662 272921
rect 371606 272847 371662 272856
rect 371700 270496 371752 270502
rect 371700 270438 371752 270444
rect 371712 270094 371740 270438
rect 371700 270088 371752 270094
rect 371700 270030 371752 270036
rect 371056 252000 371108 252006
rect 371056 251942 371108 251948
rect 371712 148578 371740 270030
rect 371804 269822 371832 374575
rect 371792 269816 371844 269822
rect 371792 269758 371844 269764
rect 371700 148572 371752 148578
rect 371700 148514 371752 148520
rect 370964 148504 371016 148510
rect 370964 148446 371016 148452
rect 371896 57458 371924 472670
rect 371988 165442 372016 479538
rect 372160 475448 372212 475454
rect 372160 475390 372212 475396
rect 372068 468580 372120 468586
rect 372068 468522 372120 468528
rect 372080 166530 372108 468522
rect 372172 271590 372200 475390
rect 372252 467424 372304 467430
rect 372252 467366 372304 467372
rect 372160 271584 372212 271590
rect 372160 271526 372212 271532
rect 372264 270881 372292 467366
rect 372448 377738 372476 479878
rect 373172 478372 373224 478378
rect 373172 478314 373224 478320
rect 373080 471708 373132 471714
rect 373080 471650 373132 471656
rect 372988 382288 373040 382294
rect 372988 382230 373040 382236
rect 372526 378448 372582 378457
rect 372526 378383 372582 378392
rect 372436 377732 372488 377738
rect 372436 377674 372488 377680
rect 372436 374672 372488 374678
rect 372436 374614 372488 374620
rect 372344 273012 372396 273018
rect 372344 272954 372396 272960
rect 372250 270872 372306 270881
rect 372250 270807 372306 270816
rect 372252 269000 372304 269006
rect 372252 268942 372304 268948
rect 372160 252408 372212 252414
rect 372160 252350 372212 252356
rect 372068 166524 372120 166530
rect 372068 166466 372120 166472
rect 371976 165436 372028 165442
rect 371976 165378 372028 165384
rect 372172 163606 372200 252350
rect 372160 163600 372212 163606
rect 372160 163542 372212 163548
rect 372264 162246 372292 268942
rect 372252 162240 372304 162246
rect 372252 162182 372304 162188
rect 372356 162178 372384 272954
rect 372448 252414 372476 374614
rect 372540 270026 372568 378383
rect 372528 270020 372580 270026
rect 372528 269962 372580 269968
rect 373000 269793 373028 382230
rect 373092 375290 373120 471650
rect 373184 376174 373212 478314
rect 373264 476876 373316 476882
rect 373264 476818 373316 476824
rect 373172 376168 373224 376174
rect 373172 376110 373224 376116
rect 373080 375284 373132 375290
rect 373080 375226 373132 375232
rect 373092 369854 373120 375226
rect 373092 369826 373212 369854
rect 373184 273018 373212 369826
rect 373172 273012 373224 273018
rect 373172 272954 373224 272960
rect 373170 270056 373226 270065
rect 373170 269991 373226 270000
rect 372986 269784 373042 269793
rect 372986 269719 373042 269728
rect 372436 252408 372488 252414
rect 372436 252350 372488 252356
rect 372436 251864 372488 251870
rect 372436 251806 372488 251812
rect 372344 162172 372396 162178
rect 372344 162114 372396 162120
rect 371976 148504 372028 148510
rect 371976 148446 372028 148452
rect 371884 57452 371936 57458
rect 371884 57394 371936 57400
rect 370596 57384 370648 57390
rect 370596 57326 370648 57332
rect 283472 57316 283524 57322
rect 283472 57258 283524 57264
rect 370504 57316 370556 57322
rect 370504 57258 370556 57264
rect 371988 55894 372016 148446
rect 372448 148374 372476 251806
rect 373184 163538 373212 269991
rect 373276 164898 373304 476818
rect 373356 472932 373408 472938
rect 373356 472874 373408 472880
rect 373368 166190 373396 472874
rect 373448 465996 373500 466002
rect 373448 465938 373500 465944
rect 373460 166666 373488 465938
rect 373552 271794 373580 482326
rect 376024 478236 376076 478242
rect 376024 478178 376076 478184
rect 375288 475516 375340 475522
rect 375288 475458 375340 475464
rect 375104 474496 375156 474502
rect 375104 474438 375156 474444
rect 374828 474292 374880 474298
rect 374828 474234 374880 474240
rect 374644 473000 374696 473006
rect 374644 472942 374696 472948
rect 374460 471436 374512 471442
rect 374460 471378 374512 471384
rect 373724 470008 373776 470014
rect 373724 469950 373776 469956
rect 373632 464432 373684 464438
rect 373632 464374 373684 464380
rect 373644 380594 373672 464374
rect 373632 380588 373684 380594
rect 373632 380530 373684 380536
rect 373736 378894 373764 469950
rect 373816 380724 373868 380730
rect 373816 380666 373868 380672
rect 373724 378888 373776 378894
rect 373630 378856 373686 378865
rect 373724 378830 373776 378836
rect 373630 378791 373686 378800
rect 373540 271788 373592 271794
rect 373540 271730 373592 271736
rect 373644 270230 373672 378791
rect 373632 270224 373684 270230
rect 373632 270166 373684 270172
rect 373736 269754 373764 378830
rect 373724 269748 373776 269754
rect 373724 269690 373776 269696
rect 373828 269006 373856 380666
rect 373906 379264 373962 379273
rect 373906 379199 373962 379208
rect 373920 378865 373948 379199
rect 373906 378856 373962 378865
rect 373906 378791 373962 378800
rect 374472 375970 374500 471378
rect 374552 378548 374604 378554
rect 374552 378490 374604 378496
rect 374564 378146 374592 378490
rect 374552 378140 374604 378146
rect 374552 378082 374604 378088
rect 374552 376032 374604 376038
rect 374552 375974 374604 375980
rect 374460 375964 374512 375970
rect 374460 375906 374512 375912
rect 374368 375420 374420 375426
rect 374368 375362 374420 375368
rect 374380 270473 374408 375362
rect 374460 274780 374512 274786
rect 374460 274722 374512 274728
rect 374472 272082 374500 274722
rect 374564 272474 374592 375974
rect 374552 272468 374604 272474
rect 374552 272410 374604 272416
rect 374472 272054 374592 272082
rect 374460 271924 374512 271930
rect 374460 271866 374512 271872
rect 374366 270464 374422 270473
rect 374366 270399 374422 270408
rect 373908 270020 373960 270026
rect 373908 269962 373960 269968
rect 373816 269000 373868 269006
rect 373816 268942 373868 268948
rect 373632 252476 373684 252482
rect 373632 252418 373684 252424
rect 373540 251932 373592 251938
rect 373540 251874 373592 251880
rect 373448 166660 373500 166666
rect 373448 166602 373500 166608
rect 373356 166184 373408 166190
rect 373356 166126 373408 166132
rect 373264 164892 373316 164898
rect 373264 164834 373316 164840
rect 373172 163532 373224 163538
rect 373172 163474 373224 163480
rect 373552 163441 373580 251874
rect 373644 165646 373672 252418
rect 373632 165640 373684 165646
rect 373632 165582 373684 165588
rect 373816 165640 373868 165646
rect 373816 165582 373868 165588
rect 373538 163432 373594 163441
rect 373538 163367 373594 163376
rect 373724 162240 373776 162246
rect 373724 162182 373776 162188
rect 372712 148436 372764 148442
rect 372712 148378 372764 148384
rect 372436 148368 372488 148374
rect 372436 148310 372488 148316
rect 372724 147626 372752 148378
rect 372712 147620 372764 147626
rect 372712 147562 372764 147568
rect 373264 147620 373316 147626
rect 373264 147562 373316 147568
rect 371976 55888 372028 55894
rect 371976 55830 372028 55836
rect 277400 55208 277452 55214
rect 277400 55150 277452 55156
rect 273352 55140 273404 55146
rect 273352 55082 273404 55088
rect 271880 55072 271932 55078
rect 271880 55014 271932 55020
rect 266452 55004 266504 55010
rect 266452 54946 266504 54952
rect 264980 54936 265032 54942
rect 264980 54878 265032 54884
rect 253940 54868 253992 54874
rect 253940 54810 253992 54816
rect 251364 54800 251416 54806
rect 251364 54742 251416 54748
rect 249800 54732 249852 54738
rect 249800 54674 249852 54680
rect 247040 54664 247092 54670
rect 247040 54606 247092 54612
rect 373276 54534 373304 147562
rect 245660 54528 245712 54534
rect 245660 54470 245712 54476
rect 373264 54528 373316 54534
rect 373264 54470 373316 54476
rect 373736 54466 373764 162182
rect 373828 56438 373856 165582
rect 373920 148646 373948 269962
rect 374368 269884 374420 269890
rect 374368 269826 374420 269832
rect 373908 148640 373960 148646
rect 373908 148582 373960 148588
rect 374380 144906 374408 269826
rect 374472 146198 374500 271866
rect 374564 271017 374592 272054
rect 374550 271008 374606 271017
rect 374550 270943 374606 270952
rect 374656 166258 374684 472942
rect 374736 465724 374788 465730
rect 374736 465666 374788 465672
rect 374644 166252 374696 166258
rect 374644 166194 374696 166200
rect 374748 164966 374776 465666
rect 374840 271046 374868 474234
rect 375012 468716 375064 468722
rect 375012 468658 375064 468664
rect 374920 468512 374972 468518
rect 374920 468454 374972 468460
rect 374932 271182 374960 468454
rect 375024 379370 375052 468658
rect 375012 379364 375064 379370
rect 375012 379306 375064 379312
rect 375012 378548 375064 378554
rect 375012 378490 375064 378496
rect 375024 274786 375052 378490
rect 375116 377534 375144 474438
rect 375196 378820 375248 378826
rect 375196 378762 375248 378768
rect 375208 378350 375236 378762
rect 375196 378344 375248 378350
rect 375196 378286 375248 378292
rect 375104 377528 375156 377534
rect 375104 377470 375156 377476
rect 375208 277394 375236 378286
rect 375300 376242 375328 475458
rect 375380 470280 375432 470286
rect 375380 470222 375432 470228
rect 375392 383654 375420 470222
rect 375392 383626 375512 383654
rect 375288 376236 375340 376242
rect 375288 376178 375340 376184
rect 375484 375426 375512 383626
rect 375472 375420 375524 375426
rect 375472 375362 375524 375368
rect 375484 375222 375512 375362
rect 375472 375216 375524 375222
rect 375472 375158 375524 375164
rect 375564 375080 375616 375086
rect 375564 375022 375616 375028
rect 375576 374814 375604 375022
rect 375748 375012 375800 375018
rect 375748 374954 375800 374960
rect 375564 374808 375616 374814
rect 375564 374750 375616 374756
rect 375288 358692 375340 358698
rect 375288 358634 375340 358640
rect 375116 277366 375236 277394
rect 375012 274780 375064 274786
rect 375012 274722 375064 274728
rect 375010 274680 375066 274689
rect 375010 274615 375066 274624
rect 374920 271176 374972 271182
rect 374920 271118 374972 271124
rect 374828 271040 374880 271046
rect 374828 270982 374880 270988
rect 374918 271008 374974 271017
rect 374918 270943 374974 270952
rect 374932 270042 374960 270943
rect 375024 270178 375052 274615
rect 375116 270298 375144 277366
rect 375196 273216 375248 273222
rect 375196 273158 375248 273164
rect 375208 271930 375236 273158
rect 375196 271924 375248 271930
rect 375196 271866 375248 271872
rect 375104 270292 375156 270298
rect 375104 270234 375156 270240
rect 375024 270150 375144 270178
rect 374932 270014 375052 270042
rect 374920 268660 374972 268666
rect 374920 268602 374972 268608
rect 374828 252544 374880 252550
rect 374828 252486 374880 252492
rect 374736 164960 374788 164966
rect 374736 164902 374788 164908
rect 374840 164778 374868 252486
rect 374564 164750 374868 164778
rect 374564 164150 374592 164750
rect 374552 164144 374604 164150
rect 374552 164086 374604 164092
rect 374460 146192 374512 146198
rect 374460 146134 374512 146140
rect 374368 144900 374420 144906
rect 374368 144842 374420 144848
rect 374564 56506 374592 164086
rect 374932 162518 374960 268602
rect 375024 164082 375052 270014
rect 375116 171134 375144 270150
rect 375300 252550 375328 358634
rect 375656 270156 375708 270162
rect 375656 270098 375708 270104
rect 375564 268252 375616 268258
rect 375564 268194 375616 268200
rect 375288 252544 375340 252550
rect 375288 252486 375340 252492
rect 375116 171106 375236 171134
rect 375012 164076 375064 164082
rect 375012 164018 375064 164024
rect 375208 163674 375236 171106
rect 375196 163668 375248 163674
rect 375196 163610 375248 163616
rect 375012 163600 375064 163606
rect 375012 163542 375064 163548
rect 374920 162512 374972 162518
rect 374920 162454 374972 162460
rect 374828 162172 374880 162178
rect 374828 162114 374880 162120
rect 374644 148572 374696 148578
rect 374644 148514 374696 148520
rect 374656 56574 374684 148514
rect 374736 146260 374788 146266
rect 374736 146202 374788 146208
rect 374748 59226 374776 146202
rect 374736 59220 374788 59226
rect 374736 59162 374788 59168
rect 374644 56568 374696 56574
rect 374644 56510 374696 56516
rect 374552 56500 374604 56506
rect 374552 56442 374604 56448
rect 373816 56432 373868 56438
rect 373816 56374 373868 56380
rect 374840 56370 374868 162114
rect 374828 56364 374880 56370
rect 374828 56306 374880 56312
rect 375024 55010 375052 163542
rect 375104 163532 375156 163538
rect 375104 163474 375156 163480
rect 375116 55078 375144 163474
rect 375208 162926 375236 163610
rect 375196 162920 375248 162926
rect 375196 162862 375248 162868
rect 375576 146266 375604 268194
rect 375564 146260 375616 146266
rect 375564 146202 375616 146208
rect 375196 146192 375248 146198
rect 375196 146134 375248 146140
rect 375208 145790 375236 146134
rect 375196 145784 375248 145790
rect 375196 145726 375248 145732
rect 375208 59362 375236 145726
rect 375576 145722 375604 146202
rect 375668 145858 375696 270098
rect 375760 268666 375788 374954
rect 375840 357536 375892 357542
rect 375840 357478 375892 357484
rect 375748 268660 375800 268666
rect 375748 268602 375800 268608
rect 375852 252482 375880 357478
rect 375932 268932 375984 268938
rect 375932 268874 375984 268880
rect 375840 252476 375892 252482
rect 375840 252418 375892 252424
rect 375944 162586 375972 268874
rect 376036 165345 376064 478178
rect 376116 476808 376168 476814
rect 376116 476750 376168 476756
rect 376022 165336 376078 165345
rect 376022 165271 376078 165280
rect 376128 164830 376156 476750
rect 376220 271561 376248 483958
rect 378784 483880 378836 483886
rect 378784 483822 378836 483828
rect 376484 481228 376536 481234
rect 376484 481170 376536 481176
rect 376300 477012 376352 477018
rect 376300 476954 376352 476960
rect 376312 272746 376340 476954
rect 376392 466200 376444 466206
rect 376392 466142 376444 466148
rect 376300 272740 376352 272746
rect 376300 272682 376352 272688
rect 376404 271697 376432 466142
rect 376496 376514 376524 481170
rect 377312 478304 377364 478310
rect 377312 478246 377364 478252
rect 376760 475584 376812 475590
rect 376760 475526 376812 475532
rect 376576 471572 376628 471578
rect 376576 471514 376628 471520
rect 376588 379642 376616 471514
rect 376772 382294 376800 475526
rect 376852 471640 376904 471646
rect 376852 471582 376904 471588
rect 376760 382288 376812 382294
rect 376760 382230 376812 382236
rect 376772 380934 376800 382230
rect 376760 380928 376812 380934
rect 376760 380870 376812 380876
rect 376668 380656 376720 380662
rect 376668 380598 376720 380604
rect 376576 379636 376628 379642
rect 376576 379578 376628 379584
rect 376588 379545 376616 379578
rect 376680 379574 376708 380598
rect 376864 379710 376892 471582
rect 377220 417444 377272 417450
rect 377220 417386 377272 417392
rect 377232 416945 377260 417386
rect 377218 416936 377274 416945
rect 377218 416871 377274 416880
rect 377126 412040 377182 412049
rect 377126 411975 377182 411984
rect 377140 411942 377168 411975
rect 377128 411936 377180 411942
rect 377128 411878 377180 411884
rect 377218 410952 377274 410961
rect 377218 410887 377274 410896
rect 377232 410582 377260 410887
rect 377220 410576 377272 410582
rect 377220 410518 377272 410524
rect 376944 391944 376996 391950
rect 376944 391886 376996 391892
rect 376956 390969 376984 391886
rect 376942 390960 376998 390969
rect 376942 390895 376998 390904
rect 376944 390516 376996 390522
rect 376944 390458 376996 390464
rect 376956 389337 376984 390458
rect 376942 389328 376998 389337
rect 376942 389263 376998 389272
rect 376944 389156 376996 389162
rect 376944 389098 376996 389104
rect 376956 389065 376984 389098
rect 376942 389056 376998 389065
rect 376942 388991 376998 389000
rect 376942 381032 376998 381041
rect 376942 380967 376998 380976
rect 376852 379704 376904 379710
rect 376852 379646 376904 379652
rect 376668 379568 376720 379574
rect 376574 379536 376630 379545
rect 376668 379510 376720 379516
rect 376574 379471 376630 379480
rect 376484 376508 376536 376514
rect 376484 376450 376536 376456
rect 376576 375080 376628 375086
rect 376576 375022 376628 375028
rect 376484 374876 376536 374882
rect 376484 374818 376536 374824
rect 376390 271688 376446 271697
rect 376390 271623 376446 271632
rect 376206 271552 376262 271561
rect 376206 271487 376262 271496
rect 376300 270360 376352 270366
rect 376300 270302 376352 270308
rect 376208 269748 376260 269754
rect 376208 269690 376260 269696
rect 376116 164824 376168 164830
rect 376116 164766 376168 164772
rect 376220 164014 376248 269690
rect 376208 164008 376260 164014
rect 376208 163950 376260 163956
rect 376312 162858 376340 270302
rect 376496 269142 376524 374818
rect 376484 269136 376536 269142
rect 376484 269078 376536 269084
rect 376496 258074 376524 269078
rect 376588 269074 376616 375022
rect 376680 269226 376708 379510
rect 376956 378185 376984 380967
rect 377324 380662 377352 478246
rect 377588 470076 377640 470082
rect 377588 470018 377640 470024
rect 377496 469940 377548 469946
rect 377496 469882 377548 469888
rect 377404 468444 377456 468450
rect 377404 468386 377456 468392
rect 377416 410310 377444 468386
rect 377508 413953 377536 469882
rect 377600 417897 377628 470018
rect 378140 468376 378192 468382
rect 378140 468318 378192 468324
rect 377586 417888 377642 417897
rect 377586 417823 377642 417832
rect 377494 413944 377550 413953
rect 377494 413879 377550 413888
rect 377494 412040 377550 412049
rect 377494 411975 377550 411984
rect 377404 410304 377456 410310
rect 377404 410246 377456 410252
rect 377402 409184 377458 409193
rect 377402 409119 377404 409128
rect 377456 409119 377458 409128
rect 377404 409090 377456 409096
rect 377312 380656 377364 380662
rect 377312 380598 377364 380604
rect 377404 379704 377456 379710
rect 377404 379646 377456 379652
rect 377416 379438 377444 379646
rect 377404 379432 377456 379438
rect 377404 379374 377456 379380
rect 376942 378176 376998 378185
rect 376942 378111 376998 378120
rect 377312 375964 377364 375970
rect 377312 375906 377364 375912
rect 377128 374944 377180 374950
rect 377128 374886 377180 374892
rect 377036 358012 377088 358018
rect 377036 357954 377088 357960
rect 376942 310856 376998 310865
rect 376942 310791 376998 310800
rect 376956 287054 376984 310791
rect 376864 287026 376984 287054
rect 376760 282872 376812 282878
rect 376760 282814 376812 282820
rect 376772 282169 376800 282814
rect 376758 282160 376814 282169
rect 376758 282095 376814 282104
rect 376864 277394 376892 287026
rect 376944 284300 376996 284306
rect 376944 284242 376996 284248
rect 376956 284073 376984 284242
rect 376942 284064 376998 284073
rect 376942 283999 376998 284008
rect 376942 282296 376998 282305
rect 376942 282231 376998 282240
rect 376956 282198 376984 282231
rect 376944 282192 376996 282198
rect 376944 282134 376996 282140
rect 376864 277366 376984 277394
rect 376680 269198 376800 269226
rect 376666 269104 376722 269113
rect 376576 269068 376628 269074
rect 376666 269039 376722 269048
rect 376576 269010 376628 269016
rect 376404 258046 376524 258074
rect 376300 162852 376352 162858
rect 376300 162794 376352 162800
rect 376404 162738 376432 258046
rect 376128 162716 376432 162738
rect 376128 162710 376300 162716
rect 375932 162580 375984 162586
rect 375932 162522 375984 162528
rect 375944 161474 375972 162522
rect 375852 161446 375972 161474
rect 375656 145852 375708 145858
rect 375656 145794 375708 145800
rect 375564 145716 375616 145722
rect 375564 145658 375616 145664
rect 375668 145602 375696 145794
rect 375300 145574 375696 145602
rect 375196 59356 375248 59362
rect 375196 59298 375248 59304
rect 375104 55072 375156 55078
rect 375104 55014 375156 55020
rect 375012 55004 375064 55010
rect 375012 54946 375064 54952
rect 375300 54670 375328 145574
rect 375852 55214 375880 161446
rect 376024 148640 376076 148646
rect 376024 148582 376076 148588
rect 375932 146192 375984 146198
rect 375932 146134 375984 146140
rect 375840 55208 375892 55214
rect 375840 55150 375892 55156
rect 375288 54664 375340 54670
rect 375288 54606 375340 54612
rect 375944 54602 375972 146134
rect 376036 55146 376064 148582
rect 376128 59158 376156 162710
rect 376352 162710 376432 162716
rect 376300 162658 376352 162664
rect 376208 162648 376260 162654
rect 376312 162627 376340 162658
rect 376392 162648 376444 162654
rect 376208 162590 376260 162596
rect 376392 162590 376444 162596
rect 376220 59566 376248 162590
rect 376208 59560 376260 59566
rect 376208 59502 376260 59508
rect 376116 59152 376168 59158
rect 376116 59094 376168 59100
rect 376404 59090 376432 162590
rect 376576 161968 376628 161974
rect 376576 161910 376628 161916
rect 376484 146260 376536 146266
rect 376484 146202 376536 146208
rect 376392 59084 376444 59090
rect 376392 59026 376444 59032
rect 376024 55140 376076 55146
rect 376024 55082 376076 55088
rect 376496 54738 376524 146202
rect 376588 59022 376616 161910
rect 376576 59016 376628 59022
rect 376576 58958 376628 58964
rect 376680 57866 376708 269039
rect 376772 268938 376800 269198
rect 376760 268932 376812 268938
rect 376760 268874 376812 268880
rect 376758 204232 376814 204241
rect 376758 204167 376814 204176
rect 376772 203017 376800 204167
rect 376956 203969 376984 277366
rect 377048 270502 377076 357954
rect 377036 270496 377088 270502
rect 377036 270438 377088 270444
rect 377140 270366 377168 374886
rect 377218 310040 377274 310049
rect 377218 309975 377274 309984
rect 377128 270360 377180 270366
rect 377128 270302 377180 270308
rect 377140 269686 377168 270302
rect 377128 269680 377180 269686
rect 377128 269622 377180 269628
rect 377128 252068 377180 252074
rect 377128 252010 377180 252016
rect 376942 203960 376998 203969
rect 376942 203895 376998 203904
rect 376758 203008 376814 203017
rect 376758 202943 376814 202952
rect 376772 95985 376800 202943
rect 376850 201376 376906 201385
rect 376850 201311 376906 201320
rect 376758 95976 376814 95985
rect 376758 95911 376814 95920
rect 376864 93809 376892 201311
rect 376956 200114 376984 203895
rect 376956 200086 377076 200114
rect 376942 198792 376998 198801
rect 376942 198727 376998 198736
rect 376956 176066 376984 198727
rect 377048 180794 377076 200086
rect 377140 190454 377168 252010
rect 377232 204241 377260 309975
rect 377324 268598 377352 375906
rect 377508 306374 377536 411975
rect 377600 310865 377628 417823
rect 377862 416936 377918 416945
rect 377862 416871 377918 416880
rect 377678 414760 377734 414769
rect 377678 414695 377680 414704
rect 377732 414695 377734 414704
rect 377680 414666 377732 414672
rect 377586 310856 377642 310865
rect 377586 310791 377642 310800
rect 377692 307873 377720 414666
rect 377770 410952 377826 410961
rect 377770 410887 377826 410896
rect 377678 307864 377734 307873
rect 377678 307799 377734 307808
rect 377508 306346 377628 306374
rect 377600 305017 377628 306346
rect 377586 305008 377642 305017
rect 377586 304943 377642 304952
rect 377402 302152 377458 302161
rect 377402 302087 377458 302096
rect 377312 268592 377364 268598
rect 377312 268534 377364 268540
rect 377324 268258 377352 268534
rect 377312 268252 377364 268258
rect 377312 268194 377364 268200
rect 377218 204232 377274 204241
rect 377218 204167 377274 204176
rect 377310 197024 377366 197033
rect 377310 196959 377366 196968
rect 377140 190426 377260 190454
rect 377048 180766 377168 180794
rect 377036 178016 377088 178022
rect 377036 177958 377088 177964
rect 377048 177041 377076 177958
rect 377034 177032 377090 177041
rect 377034 176967 377090 176976
rect 376956 176038 377076 176066
rect 376944 175976 376996 175982
rect 376944 175918 376996 175924
rect 376956 175409 376984 175918
rect 376942 175400 376998 175409
rect 376942 175335 376998 175344
rect 377048 175250 377076 176038
rect 376956 175222 377076 175250
rect 376850 93800 376906 93809
rect 376850 93735 376906 93744
rect 376956 92857 376984 175222
rect 377140 175114 377168 180766
rect 377048 175086 377168 175114
rect 377048 96937 377076 175086
rect 377232 162790 377260 190426
rect 377220 162784 377272 162790
rect 377220 162726 377272 162732
rect 377232 161974 377260 162726
rect 377220 161968 377272 161974
rect 377220 161910 377272 161916
rect 377218 145752 377274 145761
rect 377218 145687 377274 145696
rect 377034 96928 377090 96937
rect 377034 96863 377090 96872
rect 376942 92848 376998 92857
rect 376942 92783 376998 92792
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 377232 59498 377260 145687
rect 377324 90001 377352 196959
rect 377416 195265 377444 302087
rect 377496 270292 377548 270298
rect 377496 270234 377548 270240
rect 377508 269958 377536 270234
rect 377496 269952 377548 269958
rect 377496 269894 377548 269900
rect 377402 195256 377458 195265
rect 377402 195191 377458 195200
rect 377404 175228 377456 175234
rect 377404 175170 377456 175176
rect 377416 175137 377444 175170
rect 377402 175128 377458 175137
rect 377402 175063 377458 175072
rect 377404 164212 377456 164218
rect 377404 164154 377456 164160
rect 377416 163441 377444 164154
rect 377402 163432 377458 163441
rect 377402 163367 377458 163376
rect 377416 163033 377444 163367
rect 377402 163024 377458 163033
rect 377402 162959 377458 162968
rect 377508 146266 377536 269894
rect 377600 198121 377628 304943
rect 377692 201385 377720 307799
rect 377784 306374 377812 410887
rect 377876 310049 377904 416871
rect 377954 413944 378010 413953
rect 377954 413879 378010 413888
rect 377862 310040 377918 310049
rect 377862 309975 377918 309984
rect 377968 306785 377996 413879
rect 378046 409184 378102 409193
rect 378046 409119 378102 409128
rect 377954 306776 378010 306785
rect 377954 306711 378010 306720
rect 377784 306346 377904 306374
rect 377876 303929 377904 306346
rect 377862 303920 377918 303929
rect 377862 303855 377918 303864
rect 377678 201376 377734 201385
rect 377678 201311 377734 201320
rect 377692 200841 377720 201311
rect 377678 200832 377734 200841
rect 377678 200767 377734 200776
rect 377586 198112 377642 198121
rect 377586 198047 377642 198056
rect 377600 190454 377628 198047
rect 377876 197033 377904 303855
rect 377968 199889 377996 306711
rect 378060 302161 378088 409119
rect 378152 380730 378180 468318
rect 378140 380724 378192 380730
rect 378140 380666 378192 380672
rect 378140 374808 378192 374814
rect 378140 374750 378192 374756
rect 378046 302152 378102 302161
rect 378046 302087 378102 302096
rect 378152 273426 378180 374750
rect 378692 357876 378744 357882
rect 378692 357818 378744 357824
rect 378140 273420 378192 273426
rect 378140 273362 378192 273368
rect 378600 273420 378652 273426
rect 378600 273362 378652 273368
rect 378612 273154 378640 273362
rect 378600 273148 378652 273154
rect 378600 273090 378652 273096
rect 378048 270496 378100 270502
rect 378048 270438 378100 270444
rect 377954 199880 378010 199889
rect 377954 199815 378010 199824
rect 377968 198801 377996 199815
rect 377954 198792 378010 198801
rect 377954 198727 378010 198736
rect 377862 197024 377918 197033
rect 377862 196959 377918 196968
rect 377954 195256 378010 195265
rect 377954 195191 378010 195200
rect 377600 190426 377812 190454
rect 377496 146260 377548 146266
rect 377496 146202 377548 146208
rect 377508 145926 377536 146202
rect 377496 145920 377548 145926
rect 377496 145862 377548 145868
rect 377784 91089 377812 190426
rect 377864 145988 377916 145994
rect 377864 145930 377916 145936
rect 377770 91080 377826 91089
rect 377770 91015 377826 91024
rect 377310 89992 377366 90001
rect 377310 89927 377366 89936
rect 377220 59492 377272 59498
rect 377220 59434 377272 59440
rect 376668 57860 376720 57866
rect 376668 57802 376720 57808
rect 377876 54806 377904 145930
rect 377968 88233 377996 195191
rect 378060 145314 378088 270438
rect 378704 270337 378732 357818
rect 378690 270328 378746 270337
rect 378600 270292 378652 270298
rect 378690 270263 378746 270272
rect 378600 270234 378652 270240
rect 378612 146062 378640 270234
rect 378704 146169 378732 270263
rect 378796 165481 378824 483822
rect 378876 478168 378928 478174
rect 378876 478110 378928 478116
rect 378782 165472 378838 165481
rect 378782 165407 378838 165416
rect 378888 164762 378916 478110
rect 379060 474156 379112 474162
rect 379060 474098 379112 474104
rect 378968 472796 379020 472802
rect 378968 472738 379020 472744
rect 378876 164756 378928 164762
rect 378876 164698 378928 164704
rect 378980 164694 379008 472738
rect 379072 271114 379100 474098
rect 379336 471504 379388 471510
rect 379336 471446 379388 471452
rect 379152 467152 379204 467158
rect 379152 467094 379204 467100
rect 379060 271108 379112 271114
rect 379060 271050 379112 271056
rect 379164 270978 379192 467094
rect 379244 410304 379296 410310
rect 379244 410246 379296 410252
rect 379256 379710 379284 410246
rect 379244 379704 379296 379710
rect 379244 379646 379296 379652
rect 379244 377324 379296 377330
rect 379244 377266 379296 377272
rect 379152 270972 379204 270978
rect 379152 270914 379204 270920
rect 379152 269816 379204 269822
rect 379152 269758 379204 269764
rect 379164 269210 379192 269758
rect 379152 269204 379204 269210
rect 379152 269146 379204 269152
rect 379060 269068 379112 269074
rect 379060 269010 379112 269016
rect 379072 268394 379100 269010
rect 379060 268388 379112 268394
rect 379060 268330 379112 268336
rect 378968 164688 379020 164694
rect 378968 164630 379020 164636
rect 379072 151814 379100 268330
rect 379164 162654 379192 269146
rect 379256 268802 379284 377266
rect 379348 375154 379376 471446
rect 379520 380792 379572 380798
rect 379520 380734 379572 380740
rect 379532 379846 379560 380734
rect 379520 379840 379572 379846
rect 379520 379782 379572 379788
rect 379888 379840 379940 379846
rect 379888 379782 379940 379788
rect 379520 378956 379572 378962
rect 379520 378898 379572 378904
rect 379532 378418 379560 378898
rect 379704 378820 379756 378826
rect 379704 378762 379756 378768
rect 379520 378412 379572 378418
rect 379520 378354 379572 378360
rect 379336 375148 379388 375154
rect 379336 375090 379388 375096
rect 379348 273494 379376 375090
rect 379428 358760 379480 358766
rect 379428 358702 379480 358708
rect 379336 273488 379388 273494
rect 379336 273430 379388 273436
rect 379348 273222 379376 273430
rect 379336 273216 379388 273222
rect 379336 273158 379388 273164
rect 379440 270450 379468 358702
rect 379440 270422 379652 270450
rect 379624 269822 379652 270422
rect 379716 270162 379744 378762
rect 379796 378412 379848 378418
rect 379796 378354 379848 378360
rect 379808 270298 379836 378354
rect 379900 270298 379928 379782
rect 379992 378826 380020 484094
rect 429304 480962 429332 591223
rect 429396 538257 429424 647838
rect 430580 645176 430632 645182
rect 430580 645118 430632 645124
rect 429844 639464 429896 639470
rect 429844 639406 429896 639412
rect 429856 627910 429884 639406
rect 430592 634137 430620 645118
rect 430764 643204 430816 643210
rect 430764 643146 430816 643152
rect 430672 643136 430724 643142
rect 430672 643078 430724 643084
rect 430578 634128 430634 634137
rect 430578 634063 430634 634072
rect 429844 627904 429896 627910
rect 429844 627846 429896 627852
rect 430684 624617 430712 643078
rect 430776 629377 430804 643146
rect 494072 642394 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 649330 542400 702406
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 542360 649324 542412 649330
rect 542360 649266 542412 649272
rect 494060 642388 494112 642394
rect 494060 642330 494112 642336
rect 435364 641776 435416 641782
rect 435364 641718 435416 641724
rect 430854 640384 430910 640393
rect 430854 640319 430910 640328
rect 430762 629368 430818 629377
rect 430762 629303 430818 629312
rect 430670 624608 430726 624617
rect 430670 624543 430726 624552
rect 430868 619857 430896 640319
rect 432604 639532 432656 639538
rect 432604 639474 432656 639480
rect 432616 630018 432644 639474
rect 435376 630086 435404 641718
rect 457444 640348 457496 640354
rect 457444 640290 457496 640296
rect 435364 630080 435416 630086
rect 435364 630022 435416 630028
rect 432604 630012 432656 630018
rect 432604 629954 432656 629960
rect 456800 627904 456852 627910
rect 456800 627846 456852 627852
rect 456812 627745 456840 627846
rect 456798 627736 456854 627745
rect 456798 627671 456854 627680
rect 430854 619848 430910 619857
rect 430854 619783 430910 619792
rect 430578 610328 430634 610337
rect 430578 610263 430634 610272
rect 429474 596048 429530 596057
rect 429474 595983 429530 595992
rect 429382 538248 429438 538257
rect 429382 538183 429438 538192
rect 429488 526590 429516 595983
rect 429566 586664 429622 586673
rect 429566 586599 429622 586608
rect 429580 527882 429608 586599
rect 429658 557288 429714 557297
rect 429658 557223 429714 557232
rect 429568 527876 429620 527882
rect 429568 527818 429620 527824
rect 429476 526584 429528 526590
rect 429476 526526 429528 526532
rect 429672 522850 429700 557223
rect 430592 528358 430620 610263
rect 430670 605568 430726 605577
rect 430670 605503 430726 605512
rect 430580 528352 430632 528358
rect 430580 528294 430632 528300
rect 430684 528086 430712 605503
rect 457456 590345 457484 640290
rect 457536 639396 457588 639402
rect 457536 639338 457588 639344
rect 457548 621625 457576 639338
rect 470600 639328 470652 639334
rect 470600 639270 470652 639276
rect 470612 634814 470640 639270
rect 512000 639260 512052 639266
rect 512000 639202 512052 639208
rect 510620 639192 510672 639198
rect 510620 639134 510672 639140
rect 470612 634786 471192 634814
rect 471164 627994 471192 634786
rect 483204 630080 483256 630086
rect 483204 630022 483256 630028
rect 465448 627972 465500 627978
rect 465198 627920 465448 627926
rect 471164 627966 471638 627994
rect 483216 627980 483244 630022
rect 494796 630012 494848 630018
rect 494796 629954 494848 629960
rect 494808 627980 494836 629954
rect 501236 629944 501288 629950
rect 501236 629886 501288 629892
rect 501248 627980 501276 629886
rect 465198 627914 465500 627920
rect 465198 627898 465488 627914
rect 477130 627872 477186 627881
rect 488722 627872 488778 627881
rect 477186 627830 477434 627858
rect 477130 627807 477186 627816
rect 506754 627872 506810 627881
rect 488778 627830 489026 627858
rect 488722 627807 488778 627816
rect 506810 627830 507058 627858
rect 506754 627807 506810 627816
rect 457534 621616 457590 621625
rect 457534 621551 457590 621560
rect 510632 618905 510660 639134
rect 510618 618896 510674 618905
rect 510618 618831 510674 618840
rect 457626 615496 457682 615505
rect 457626 615431 457682 615440
rect 457534 596456 457590 596465
rect 457534 596391 457590 596400
rect 457442 590336 457498 590345
rect 457442 590271 457498 590280
rect 457442 584216 457498 584225
rect 457442 584151 457498 584160
rect 430762 581088 430818 581097
rect 430762 581023 430818 581032
rect 430672 528080 430724 528086
rect 430672 528022 430724 528028
rect 430776 526726 430804 581023
rect 430854 576328 430910 576337
rect 430854 576263 430910 576272
rect 430868 527950 430896 576263
rect 430946 571568 431002 571577
rect 430946 571503 431002 571512
rect 430856 527944 430908 527950
rect 430856 527886 430908 527892
rect 430960 526794 430988 571503
rect 431038 562048 431094 562057
rect 431038 561983 431094 561992
rect 430948 526788 431000 526794
rect 430948 526730 431000 526736
rect 430764 526720 430816 526726
rect 430764 526662 430816 526668
rect 431052 526658 431080 561983
rect 431130 552528 431186 552537
rect 431130 552463 431186 552472
rect 431144 528018 431172 552463
rect 431222 547768 431278 547777
rect 431222 547703 431278 547712
rect 431236 528290 431264 547703
rect 431314 543008 431370 543017
rect 431314 542943 431370 542952
rect 431224 528284 431276 528290
rect 431224 528226 431276 528232
rect 431328 528222 431356 542943
rect 431406 533488 431462 533497
rect 431406 533423 431462 533432
rect 431316 528216 431368 528222
rect 431316 528158 431368 528164
rect 431420 528154 431448 533423
rect 457456 528426 457484 584151
rect 457444 528420 457496 528426
rect 457444 528362 457496 528368
rect 431408 528148 431460 528154
rect 431408 528090 431460 528096
rect 431132 528012 431184 528018
rect 431132 527954 431184 527960
rect 431040 526652 431092 526658
rect 431040 526594 431092 526600
rect 429660 522844 429712 522850
rect 429660 522786 429712 522792
rect 429292 480956 429344 480962
rect 429292 480898 429344 480904
rect 457548 478145 457576 596391
rect 457640 526862 457668 615431
rect 512012 612105 512040 639202
rect 580264 639124 580316 639130
rect 580264 639066 580316 639072
rect 512092 637628 512144 637634
rect 512092 637570 512144 637576
rect 512104 625025 512132 637570
rect 580276 630873 580304 639066
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580264 627972 580316 627978
rect 580264 627914 580316 627920
rect 512090 625016 512146 625025
rect 512090 624951 512146 624960
rect 511998 612096 512054 612105
rect 511998 612031 512054 612040
rect 457718 609376 457774 609385
rect 457718 609311 457774 609320
rect 457628 526856 457680 526862
rect 457628 526798 457680 526804
rect 457732 522918 457760 609311
rect 511998 605976 512054 605985
rect 511998 605911 512054 605920
rect 457810 602576 457866 602585
rect 457810 602511 457866 602520
rect 457824 526998 457852 602511
rect 459572 578054 460046 578082
rect 465092 578054 465842 578082
rect 470612 578054 471638 578082
rect 476132 578054 477434 578082
rect 483032 578054 483230 578082
rect 488552 578054 489670 578082
rect 457812 526992 457864 526998
rect 457812 526934 457864 526940
rect 459572 526930 459600 578054
rect 459560 526924 459612 526930
rect 459560 526866 459612 526872
rect 465092 522986 465120 578054
rect 470612 524278 470640 578054
rect 476132 528494 476160 578054
rect 476120 528488 476172 528494
rect 476120 528430 476172 528436
rect 470600 524272 470652 524278
rect 470600 524214 470652 524220
rect 465080 522980 465132 522986
rect 465080 522922 465132 522928
rect 457720 522912 457772 522918
rect 457720 522854 457772 522860
rect 457534 478136 457590 478145
rect 457534 478071 457590 478080
rect 483032 475425 483060 578054
rect 488552 524346 488580 578054
rect 495452 528562 495480 578068
rect 500972 578054 501262 578082
rect 506492 578054 507058 578082
rect 495440 528556 495492 528562
rect 495440 528498 495492 528504
rect 500972 527066 501000 578054
rect 500960 527060 501012 527066
rect 500960 527002 501012 527008
rect 488540 524340 488592 524346
rect 488540 524282 488592 524288
rect 506492 487801 506520 578054
rect 506478 487792 506534 487801
rect 506478 487727 506534 487736
rect 512012 485217 512040 605911
rect 512182 599856 512238 599865
rect 512182 599791 512238 599800
rect 512090 593736 512146 593745
rect 512090 593671 512146 593680
rect 511998 485208 512054 485217
rect 511998 485143 512054 485152
rect 512104 479505 512132 593671
rect 512196 524414 512224 599791
rect 512274 587616 512330 587625
rect 512274 587551 512330 587560
rect 512288 527134 512316 587551
rect 513010 580816 513066 580825
rect 513010 580751 513066 580760
rect 513024 579698 513052 580751
rect 513012 579692 513064 579698
rect 513012 579634 513064 579640
rect 560944 579692 560996 579698
rect 560944 579634 560996 579640
rect 512276 527128 512328 527134
rect 512276 527070 512328 527076
rect 512184 524408 512236 524414
rect 512184 524350 512236 524356
rect 560956 511970 560984 579634
rect 580276 577697 580304 627914
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 578884 523728 578936 523734
rect 578884 523670 578936 523676
rect 560944 511964 560996 511970
rect 560944 511906 560996 511912
rect 520924 495508 520976 495514
rect 520924 495450 520976 495456
rect 512090 479496 512146 479505
rect 512090 479431 512146 479440
rect 483018 475416 483074 475425
rect 483018 475351 483074 475360
rect 498200 466608 498252 466614
rect 498198 466576 498200 466585
rect 517796 466608 517848 466614
rect 498252 466576 498254 466585
rect 498198 466511 498254 466520
rect 499762 466576 499818 466585
rect 499762 466511 499764 466520
rect 498212 466478 498240 466511
rect 499816 466511 499818 466520
rect 510894 466576 510950 466585
rect 517796 466550 517848 466556
rect 510894 466511 510896 466520
rect 499764 466482 499816 466488
rect 510948 466511 510950 466520
rect 517520 466540 517572 466546
rect 510896 466482 510948 466488
rect 517520 466482 517572 466488
rect 498200 466472 498252 466478
rect 498200 466414 498252 466420
rect 421748 380928 421800 380934
rect 421748 380870 421800 380876
rect 421760 380769 421788 380870
rect 421102 380760 421158 380769
rect 421102 380695 421158 380704
rect 421746 380760 421802 380769
rect 421746 380695 421802 380704
rect 425978 380760 426034 380769
rect 425978 380695 426034 380704
rect 433614 380760 433670 380769
rect 433614 380695 433670 380704
rect 434350 380760 434406 380769
rect 434350 380695 434352 380704
rect 408682 380624 408738 380633
rect 408682 380559 408738 380568
rect 413466 380624 413522 380633
rect 413466 380559 413522 380568
rect 408696 379846 408724 380559
rect 408684 379840 408736 379846
rect 408684 379782 408736 379788
rect 413480 379778 413508 380559
rect 421116 380526 421144 380695
rect 425992 380662 426020 380695
rect 425980 380656 426032 380662
rect 422850 380624 422906 380633
rect 422850 380559 422906 380568
rect 425242 380624 425298 380633
rect 425980 380598 426032 380604
rect 433628 380594 433656 380695
rect 434404 380695 434406 380704
rect 436006 380760 436062 380769
rect 436006 380695 436062 380704
rect 438490 380760 438546 380769
rect 438490 380695 438546 380704
rect 440882 380760 440938 380769
rect 440882 380695 440938 380704
rect 443458 380760 443514 380769
rect 443458 380695 443514 380704
rect 434352 380666 434404 380672
rect 425242 380559 425298 380568
rect 433616 380588 433668 380594
rect 421104 380520 421156 380526
rect 421104 380462 421156 380468
rect 381084 379772 381136 379778
rect 381084 379714 381136 379720
rect 413468 379772 413520 379778
rect 413468 379714 413520 379720
rect 380900 379704 380952 379710
rect 380900 379646 380952 379652
rect 379980 378820 380032 378826
rect 379980 378762 380032 378768
rect 379980 377460 380032 377466
rect 379980 377402 380032 377408
rect 379796 270292 379848 270298
rect 379796 270234 379848 270240
rect 379888 270292 379940 270298
rect 379888 270234 379940 270240
rect 379704 270156 379756 270162
rect 379704 270098 379756 270104
rect 379900 269890 379928 270234
rect 379888 269884 379940 269890
rect 379888 269826 379940 269832
rect 379612 269816 379664 269822
rect 379612 269758 379664 269764
rect 379244 268796 379296 268802
rect 379244 268738 379296 268744
rect 379152 162648 379204 162654
rect 379152 162590 379204 162596
rect 379152 162512 379204 162518
rect 379152 162454 379204 162460
rect 379164 161498 379192 162454
rect 379152 161492 379204 161498
rect 379152 161434 379204 161440
rect 378980 151786 379100 151814
rect 378980 146198 379008 151786
rect 379058 146296 379114 146305
rect 379058 146231 379114 146240
rect 378968 146192 379020 146198
rect 378690 146160 378746 146169
rect 378968 146134 379020 146140
rect 378690 146095 378746 146104
rect 378600 146056 378652 146062
rect 378600 145998 378652 146004
rect 378048 145308 378100 145314
rect 378048 145250 378100 145256
rect 377954 88224 378010 88233
rect 377954 88159 378010 88168
rect 378060 54874 378088 145250
rect 378612 56030 378640 145998
rect 379072 145897 379100 146231
rect 379058 145888 379114 145897
rect 379058 145823 379114 145832
rect 378784 145648 378836 145654
rect 378784 145590 378836 145596
rect 378796 144906 378824 145590
rect 378968 145512 379020 145518
rect 378968 145454 379020 145460
rect 378876 145444 378928 145450
rect 378876 145386 378928 145392
rect 378784 144900 378836 144906
rect 378784 144842 378836 144848
rect 378600 56024 378652 56030
rect 378600 55966 378652 55972
rect 378796 55962 378824 144842
rect 378888 59702 378916 145386
rect 378980 59770 379008 145454
rect 378968 59764 379020 59770
rect 378968 59706 379020 59712
rect 378876 59696 378928 59702
rect 378876 59638 378928 59644
rect 379072 57254 379100 145823
rect 379164 59634 379192 161434
rect 379256 145994 379284 268738
rect 379428 147688 379480 147694
rect 379428 147630 379480 147636
rect 379336 146260 379388 146266
rect 379336 146202 379388 146208
rect 379244 145988 379296 145994
rect 379244 145930 379296 145936
rect 379152 59628 379204 59634
rect 379152 59570 379204 59576
rect 379060 57248 379112 57254
rect 379060 57190 379112 57196
rect 379348 56098 379376 146202
rect 379440 56302 379468 147630
rect 379624 146266 379652 269758
rect 379992 268870 380020 377402
rect 380912 357882 380940 379646
rect 380990 379400 381046 379409
rect 380990 379335 381046 379344
rect 381004 378865 381032 379335
rect 380990 378856 381046 378865
rect 380990 378791 381046 378800
rect 381096 378706 381124 379714
rect 422864 379642 422892 380559
rect 425256 379710 425284 380559
rect 433616 380530 433668 380536
rect 436020 380458 436048 380695
rect 436926 380624 436982 380633
rect 436926 380559 436982 380568
rect 436008 380452 436060 380458
rect 436008 380394 436060 380400
rect 425244 379704 425296 379710
rect 425244 379646 425296 379652
rect 422852 379636 422904 379642
rect 422852 379578 422904 379584
rect 436940 379574 436968 380559
rect 438504 380390 438532 380695
rect 438492 380384 438544 380390
rect 438492 380326 438544 380332
rect 440896 380322 440924 380695
rect 440884 380316 440936 380322
rect 440884 380258 440936 380264
rect 443472 380254 443500 380695
rect 465906 380624 465962 380633
rect 465906 380559 465962 380568
rect 443460 380248 443512 380254
rect 443460 380190 443512 380196
rect 465920 380186 465948 380559
rect 465908 380180 465960 380186
rect 465908 380122 465960 380128
rect 436928 379568 436980 379574
rect 436928 379510 436980 379516
rect 439044 379500 439096 379506
rect 439044 379442 439096 379448
rect 427452 379432 427504 379438
rect 396170 379400 396226 379409
rect 396170 379335 396226 379344
rect 405738 379400 405794 379409
rect 405738 379335 405794 379344
rect 407578 379400 407634 379409
rect 407578 379335 407634 379344
rect 408314 379400 408370 379409
rect 408314 379335 408316 379344
rect 381268 379024 381320 379030
rect 381268 378966 381320 378972
rect 381174 378856 381230 378865
rect 381174 378791 381230 378800
rect 381004 378678 381124 378706
rect 381004 358766 381032 378678
rect 381082 378584 381138 378593
rect 381082 378519 381138 378528
rect 380992 358760 381044 358766
rect 380992 358702 381044 358708
rect 381096 358698 381124 378519
rect 381084 358692 381136 358698
rect 381084 358634 381136 358640
rect 380900 357876 380952 357882
rect 380900 357818 380952 357824
rect 381188 357542 381216 378791
rect 381280 378486 381308 378966
rect 396184 378894 396212 379335
rect 402978 379264 403034 379273
rect 402978 379199 403034 379208
rect 405370 379264 405426 379273
rect 405370 379199 405426 379208
rect 396172 378888 396224 378894
rect 396172 378830 396224 378836
rect 396078 378584 396134 378593
rect 396078 378519 396080 378528
rect 396132 378519 396134 378528
rect 396080 378490 396132 378496
rect 381268 378480 381320 378486
rect 381268 378422 381320 378428
rect 381280 358018 381308 378422
rect 402992 377398 403020 379199
rect 403622 378584 403678 378593
rect 403622 378519 403678 378528
rect 402980 377392 403032 377398
rect 402980 377334 403032 377340
rect 403636 375970 403664 378519
rect 403624 375964 403676 375970
rect 403624 375906 403676 375912
rect 405384 375086 405412 379199
rect 405752 378826 405780 379335
rect 405740 378820 405792 378826
rect 405740 378762 405792 378768
rect 407592 378350 407620 379335
rect 408368 379335 408370 379344
rect 410614 379400 410670 379409
rect 410614 379335 410670 379344
rect 411258 379400 411314 379409
rect 411258 379335 411314 379344
rect 412362 379400 412418 379409
rect 412362 379335 412418 379344
rect 413098 379400 413154 379409
rect 413098 379335 413154 379344
rect 423402 379400 423458 379409
rect 423402 379335 423458 379344
rect 427450 379400 427452 379409
rect 439056 379409 439084 379442
rect 427504 379400 427506 379409
rect 427450 379335 427506 379344
rect 439042 379400 439098 379409
rect 439042 379335 439098 379344
rect 445850 379400 445906 379409
rect 445850 379335 445906 379344
rect 448150 379400 448206 379409
rect 448150 379335 448206 379344
rect 451002 379400 451058 379409
rect 451002 379335 451058 379344
rect 452750 379400 452806 379409
rect 452750 379335 452806 379344
rect 455510 379400 455566 379409
rect 455510 379335 455566 379344
rect 458362 379400 458418 379409
rect 458362 379335 458418 379344
rect 408316 379306 408368 379312
rect 409970 379264 410026 379273
rect 409970 379199 410026 379208
rect 407580 378344 407632 378350
rect 407580 378286 407632 378292
rect 409984 377330 410012 379199
rect 410628 377602 410656 379335
rect 411272 378418 411300 379335
rect 412376 378486 412404 379335
rect 412364 378480 412416 378486
rect 412364 378422 412416 378428
rect 411260 378412 411312 378418
rect 411260 378354 411312 378360
rect 410616 377596 410668 377602
rect 410616 377538 410668 377544
rect 413112 377534 413140 379335
rect 414570 379264 414626 379273
rect 414570 379199 414626 379208
rect 415398 379264 415454 379273
rect 415398 379199 415454 379208
rect 416042 379264 416098 379273
rect 416042 379199 416098 379208
rect 418342 379264 418398 379273
rect 418342 379199 418398 379208
rect 413100 377528 413152 377534
rect 413100 377470 413152 377476
rect 414584 377466 414612 379199
rect 414572 377460 414624 377466
rect 414572 377402 414624 377408
rect 409972 377324 410024 377330
rect 409972 377266 410024 377272
rect 415412 376038 415440 379199
rect 416056 376106 416084 379199
rect 418250 378856 418306 378865
rect 418250 378791 418306 378800
rect 416962 378176 417018 378185
rect 416962 378111 417018 378120
rect 418158 378176 418214 378185
rect 418158 378111 418214 378120
rect 416044 376100 416096 376106
rect 416044 376042 416096 376048
rect 415400 376032 415452 376038
rect 415400 375974 415452 375980
rect 405372 375080 405424 375086
rect 405372 375022 405424 375028
rect 416976 375018 417004 378111
rect 416964 375012 417016 375018
rect 416964 374954 417016 374960
rect 418172 374950 418200 378111
rect 418264 376310 418292 378791
rect 418252 376304 418304 376310
rect 418252 376246 418304 376252
rect 418160 374944 418212 374950
rect 418160 374886 418212 374892
rect 418356 374882 418384 379199
rect 419814 378176 419870 378185
rect 419814 378111 419870 378120
rect 418344 374876 418396 374882
rect 418344 374818 418396 374824
rect 419828 374649 419856 378111
rect 423416 377670 423444 379335
rect 437754 379264 437810 379273
rect 437754 379199 437810 379208
rect 428186 378584 428242 378593
rect 428186 378519 428242 378528
rect 430670 378584 430726 378593
rect 430670 378519 430726 378528
rect 423954 378176 424010 378185
rect 423954 378111 424010 378120
rect 426438 378176 426494 378185
rect 426438 378111 426494 378120
rect 423404 377664 423456 377670
rect 423404 377606 423456 377612
rect 423968 375154 423996 378111
rect 423956 375148 424008 375154
rect 423956 375090 424008 375096
rect 426452 374814 426480 378111
rect 428200 376174 428228 378519
rect 428278 378312 428334 378321
rect 428278 378247 428334 378256
rect 428188 376168 428240 376174
rect 428188 376110 428240 376116
rect 428292 375358 428320 378247
rect 429382 378176 429438 378185
rect 429382 378111 429438 378120
rect 428280 375352 428332 375358
rect 428280 375294 428332 375300
rect 426440 374808 426492 374814
rect 426440 374750 426492 374756
rect 429396 374746 429424 378111
rect 430684 376242 430712 378519
rect 431130 378176 431186 378185
rect 431130 378111 431186 378120
rect 432234 378176 432290 378185
rect 432234 378111 432290 378120
rect 430672 376236 430724 376242
rect 430672 376178 430724 376184
rect 431144 375290 431172 378111
rect 431132 375284 431184 375290
rect 431132 375226 431184 375232
rect 432248 375222 432276 378111
rect 432236 375216 432288 375222
rect 432236 375158 432288 375164
rect 429384 374740 429436 374746
rect 429384 374682 429436 374688
rect 437768 374678 437796 379199
rect 439056 378350 439084 379335
rect 439044 378344 439096 378350
rect 439044 378286 439096 378292
rect 445864 377806 445892 379335
rect 448164 377942 448192 379335
rect 448152 377936 448204 377942
rect 448152 377878 448204 377884
rect 451016 377874 451044 379335
rect 452764 378010 452792 379335
rect 452752 378004 452804 378010
rect 452752 377946 452804 377952
rect 451004 377868 451056 377874
rect 451004 377810 451056 377816
rect 445852 377800 445904 377806
rect 445852 377742 445904 377748
rect 455524 377738 455552 379335
rect 458376 378078 458404 379335
rect 463514 379264 463570 379273
rect 463514 379199 463570 379208
rect 473450 379264 473506 379273
rect 473450 379199 473506 379208
rect 474738 379264 474794 379273
rect 474738 379199 474794 379208
rect 480810 379264 480866 379273
rect 480810 379199 480866 379208
rect 503074 379264 503130 379273
rect 503074 379199 503130 379208
rect 503534 379264 503590 379273
rect 503534 379199 503590 379208
rect 458364 378072 458416 378078
rect 458364 378014 458416 378020
rect 455512 377732 455564 377738
rect 455512 377674 455564 377680
rect 463528 376378 463556 379199
rect 467930 378856 467986 378865
rect 467930 378791 467986 378800
rect 470874 378856 470930 378865
rect 470874 378791 470930 378800
rect 467944 376446 467972 378791
rect 470888 376582 470916 378791
rect 473464 376718 473492 379199
rect 474752 377262 474780 379199
rect 477590 378856 477646 378865
rect 477590 378791 477646 378800
rect 474740 377256 474792 377262
rect 474740 377198 474792 377204
rect 473452 376712 473504 376718
rect 473452 376654 473504 376660
rect 477604 376650 477632 378791
rect 480824 376689 480852 379199
rect 483386 378856 483442 378865
rect 483386 378791 483442 378800
rect 480810 376680 480866 376689
rect 477592 376644 477644 376650
rect 480810 376615 480866 376624
rect 477592 376586 477644 376592
rect 470876 376576 470928 376582
rect 470876 376518 470928 376524
rect 483400 376514 483428 378791
rect 503088 378282 503116 379199
rect 503076 378276 503128 378282
rect 503076 378218 503128 378224
rect 503548 378214 503576 379199
rect 516600 378344 516652 378350
rect 516600 378286 516652 378292
rect 503536 378208 503588 378214
rect 503536 378150 503588 378156
rect 483388 376508 483440 376514
rect 483388 376450 483440 376456
rect 467932 376440 467984 376446
rect 467932 376382 467984 376388
rect 463516 376372 463568 376378
rect 463516 376314 463568 376320
rect 437756 374672 437808 374678
rect 419814 374640 419870 374649
rect 437756 374614 437808 374620
rect 419814 374575 419870 374584
rect 500776 359712 500828 359718
rect 500776 359654 500828 359660
rect 498936 359576 498988 359582
rect 498936 359518 498988 359524
rect 498948 358873 498976 359518
rect 500788 358873 500816 359654
rect 498934 358864 498990 358873
rect 498934 358799 498990 358808
rect 500774 358864 500830 358873
rect 500774 358799 500830 358808
rect 510894 358864 510950 358873
rect 510894 358799 510896 358808
rect 510948 358799 510950 358808
rect 510896 358770 510948 358776
rect 381268 358012 381320 358018
rect 381268 357954 381320 357960
rect 381176 357536 381228 357542
rect 381176 357478 381228 357484
rect 421102 273592 421158 273601
rect 421102 273527 421158 273536
rect 451002 273592 451058 273601
rect 451002 273527 451058 273536
rect 421116 273358 421144 273527
rect 421104 273352 421156 273358
rect 421104 273294 421156 273300
rect 423402 273320 423458 273329
rect 423402 273255 423458 273264
rect 423770 273320 423826 273329
rect 423770 273255 423826 273264
rect 426438 273320 426494 273329
rect 451016 273290 451044 273527
rect 426438 273255 426494 273264
rect 451004 273284 451056 273290
rect 423416 273086 423444 273255
rect 423784 273222 423812 273255
rect 423772 273216 423824 273222
rect 423772 273158 423824 273164
rect 426452 273154 426480 273255
rect 451004 273226 451056 273232
rect 426440 273148 426492 273154
rect 426440 273090 426492 273096
rect 423404 273080 423456 273086
rect 423404 273022 423456 273028
rect 431132 273012 431184 273018
rect 431132 272954 431184 272960
rect 425980 272944 426032 272950
rect 425980 272886 426032 272892
rect 425992 272785 426020 272886
rect 428188 272876 428240 272882
rect 428188 272818 428240 272824
rect 428200 272785 428228 272818
rect 431144 272785 431172 272954
rect 468484 272808 468536 272814
rect 425978 272776 426034 272785
rect 425978 272711 426034 272720
rect 428186 272776 428242 272785
rect 428186 272711 428242 272720
rect 431130 272776 431186 272785
rect 431130 272711 431186 272720
rect 468482 272776 468484 272785
rect 468536 272776 468538 272785
rect 468482 272711 468538 272720
rect 470874 272776 470930 272785
rect 470874 272711 470930 272720
rect 473450 272776 473506 272785
rect 473450 272711 473452 272720
rect 470888 272678 470916 272711
rect 473504 272711 473506 272720
rect 473452 272682 473504 272688
rect 470876 272672 470928 272678
rect 470876 272614 470928 272620
rect 475842 272640 475898 272649
rect 475842 272575 475844 272584
rect 475896 272575 475898 272584
rect 478418 272640 478474 272649
rect 478418 272575 478474 272584
rect 475844 272546 475896 272552
rect 478432 272542 478460 272575
rect 478420 272536 478472 272542
rect 478420 272478 478472 272484
rect 396724 272468 396776 272474
rect 396724 272410 396776 272416
rect 396736 271289 396764 272410
rect 401690 272232 401746 272241
rect 401690 272167 401746 272176
rect 416042 272232 416098 272241
rect 416042 272167 416098 272176
rect 437938 272232 437994 272241
rect 437938 272167 437994 272176
rect 455786 272232 455842 272241
rect 455786 272167 455842 272176
rect 396722 271280 396778 271289
rect 396722 271215 396778 271224
rect 396078 270600 396134 270609
rect 396078 270535 396134 270544
rect 389272 269884 389324 269890
rect 389272 269826 389324 269832
rect 389284 269793 389312 269826
rect 389270 269784 389326 269793
rect 396092 269754 396120 270535
rect 389270 269719 389326 269728
rect 396080 269748 396132 269754
rect 389180 269204 389232 269210
rect 389180 269146 389232 269152
rect 383396 269074 383608 269090
rect 383396 269068 383620 269074
rect 383396 269062 383568 269068
rect 383396 268938 383424 269062
rect 383568 269010 383620 269016
rect 383384 268932 383436 268938
rect 383384 268874 383436 268880
rect 383476 268932 383528 268938
rect 383476 268874 383528 268880
rect 379980 268864 380032 268870
rect 379980 268806 380032 268812
rect 379992 258074 380020 268806
rect 383488 268666 383516 268874
rect 389192 268734 389220 269146
rect 389180 268728 389232 268734
rect 389180 268670 389232 268676
rect 383476 268660 383528 268666
rect 383476 268602 383528 268608
rect 389284 258074 389312 269719
rect 396080 269690 396132 269696
rect 391940 269680 391992 269686
rect 391940 269622 391992 269628
rect 390560 269136 390612 269142
rect 390560 269078 390612 269084
rect 390572 268666 390600 269078
rect 390560 268660 390612 268666
rect 390560 268602 390612 268608
rect 391952 268530 391980 269622
rect 391940 268524 391992 268530
rect 391940 268466 391992 268472
rect 379900 258046 380020 258074
rect 389192 258046 389312 258074
rect 379704 252000 379756 252006
rect 379704 251942 379756 251948
rect 379716 149054 379744 251942
rect 379796 162852 379848 162858
rect 379796 162794 379848 162800
rect 379808 162314 379836 162794
rect 379796 162308 379848 162314
rect 379796 162250 379848 162256
rect 379704 149048 379756 149054
rect 379704 148990 379756 148996
rect 379716 147694 379744 148990
rect 379704 147688 379756 147694
rect 379704 147630 379756 147636
rect 379612 146260 379664 146266
rect 379612 146202 379664 146208
rect 379702 145616 379758 145625
rect 379702 145551 379758 145560
rect 379428 56296 379480 56302
rect 379428 56238 379480 56244
rect 379716 56234 379744 145551
rect 379808 59294 379836 162250
rect 379900 145382 379928 258046
rect 389192 252074 389220 258046
rect 389180 252068 389232 252074
rect 389180 252010 389232 252016
rect 396736 251841 396764 271215
rect 397458 270600 397514 270609
rect 397458 270535 397514 270544
rect 398838 270600 398894 270609
rect 398838 270535 398894 270544
rect 400218 270600 400274 270609
rect 400218 270535 400274 270544
rect 397472 270094 397500 270535
rect 397460 270088 397512 270094
rect 397460 270030 397512 270036
rect 398852 270026 398880 270535
rect 400232 270230 400260 270535
rect 401704 270434 401732 272167
rect 402980 271924 403032 271930
rect 402980 271866 403032 271872
rect 402992 271833 403020 271866
rect 402978 271824 403034 271833
rect 402978 271759 403034 271768
rect 412822 271824 412878 271833
rect 412822 271759 412878 271768
rect 412836 271425 412864 271759
rect 412822 271416 412878 271425
rect 412822 271351 412878 271360
rect 413098 271280 413154 271289
rect 413098 271215 413154 271224
rect 413112 271182 413140 271215
rect 413100 271176 413152 271182
rect 409878 271144 409934 271153
rect 413100 271118 413152 271124
rect 414018 271144 414074 271153
rect 409878 271079 409934 271088
rect 416056 271114 416084 272167
rect 437952 271998 437980 272167
rect 421564 271992 421616 271998
rect 421564 271934 421616 271940
rect 437940 271992 437992 271998
rect 437940 271934 437992 271940
rect 416778 271144 416834 271153
rect 414018 271079 414074 271088
rect 416044 271108 416096 271114
rect 409892 271046 409920 271079
rect 409880 271040 409932 271046
rect 404358 271008 404414 271017
rect 404358 270943 404414 270952
rect 407118 271008 407174 271017
rect 409880 270982 409932 270988
rect 411258 271008 411314 271017
rect 407118 270943 407120 270952
rect 403530 270600 403586 270609
rect 403530 270535 403586 270544
rect 401692 270428 401744 270434
rect 401692 270370 401744 270376
rect 400220 270224 400272 270230
rect 400220 270166 400272 270172
rect 398840 270020 398892 270026
rect 398840 269962 398892 269968
rect 403544 268598 403572 270535
rect 403532 268592 403584 268598
rect 403532 268534 403584 268540
rect 404372 268394 404400 270943
rect 407172 270943 407174 270952
rect 411258 270943 411314 270952
rect 407120 270914 407172 270920
rect 405738 270600 405794 270609
rect 405738 270535 405794 270544
rect 407118 270600 407174 270609
rect 407118 270535 407174 270544
rect 408498 270600 408554 270609
rect 408498 270535 408554 270544
rect 409878 270600 409934 270609
rect 409878 270535 409934 270544
rect 405752 270162 405780 270535
rect 405740 270156 405792 270162
rect 405740 270098 405792 270104
rect 407132 269958 407160 270535
rect 408512 270298 408540 270535
rect 408500 270292 408552 270298
rect 408500 270234 408552 270240
rect 407120 269952 407172 269958
rect 407120 269894 407172 269900
rect 409892 268802 409920 270535
rect 411272 270502 411300 270943
rect 412914 270736 412970 270745
rect 412914 270671 412970 270680
rect 411350 270600 411406 270609
rect 411350 270535 411406 270544
rect 411260 270496 411312 270502
rect 411260 270438 411312 270444
rect 411364 270366 411392 270535
rect 411352 270360 411404 270366
rect 411352 270302 411404 270308
rect 412928 269822 412956 270671
rect 412916 269816 412968 269822
rect 412916 269758 412968 269764
rect 414032 268870 414060 271079
rect 416778 271079 416834 271088
rect 416044 271050 416096 271056
rect 416792 268938 416820 271079
rect 418250 270736 418306 270745
rect 418250 270671 418306 270680
rect 418158 270600 418214 270609
rect 418158 270535 418214 270544
rect 416780 268932 416832 268938
rect 416780 268874 416832 268880
rect 414020 268864 414072 268870
rect 414020 268806 414072 268812
rect 409880 268796 409932 268802
rect 409880 268738 409932 268744
rect 418172 268530 418200 270535
rect 418264 268666 418292 270671
rect 419538 270600 419594 270609
rect 419538 270535 419594 270544
rect 420918 270600 420974 270609
rect 420918 270535 420974 270544
rect 419552 268734 419580 270535
rect 420932 269890 420960 270535
rect 420920 269884 420972 269890
rect 420920 269826 420972 269832
rect 419540 268728 419592 268734
rect 419540 268670 419592 268676
rect 418252 268660 418304 268666
rect 418252 268602 418304 268608
rect 418160 268524 418212 268530
rect 418160 268466 418212 268472
rect 404360 268388 404412 268394
rect 404360 268330 404412 268336
rect 421576 251938 421604 271934
rect 455800 271862 455828 272167
rect 455788 271856 455840 271862
rect 433338 271824 433394 271833
rect 433338 271759 433394 271768
rect 434718 271824 434774 271833
rect 434718 271759 434774 271768
rect 437478 271824 437534 271833
rect 437478 271759 437534 271768
rect 445758 271824 445814 271833
rect 445758 271759 445814 271768
rect 447138 271824 447194 271833
rect 447138 271759 447194 271768
rect 452658 271824 452714 271833
rect 455788 271798 455840 271804
rect 458178 271824 458234 271833
rect 452658 271759 452714 271768
rect 458178 271759 458180 271768
rect 433352 271454 433380 271759
rect 433340 271448 433392 271454
rect 433340 271390 433392 271396
rect 434732 271318 434760 271759
rect 437492 271522 437520 271759
rect 445772 271658 445800 271759
rect 445760 271652 445812 271658
rect 445760 271594 445812 271600
rect 447152 271590 447180 271759
rect 452672 271726 452700 271759
rect 458232 271759 458234 271768
rect 458180 271730 458232 271736
rect 452660 271720 452712 271726
rect 452660 271662 452712 271668
rect 503626 271688 503682 271697
rect 503626 271623 503682 271632
rect 447140 271584 447192 271590
rect 447140 271526 447192 271532
rect 437480 271516 437532 271522
rect 437480 271458 437532 271464
rect 440238 271416 440294 271425
rect 503640 271386 503668 271623
rect 440238 271351 440240 271360
rect 440292 271351 440294 271360
rect 503628 271380 503680 271386
rect 440240 271322 440292 271328
rect 503628 271322 503680 271328
rect 434720 271312 434772 271318
rect 434720 271254 434772 271260
rect 440146 271280 440202 271289
rect 440146 271215 440202 271224
rect 442998 271280 443054 271289
rect 442998 271215 443000 271224
rect 440160 271182 440188 271215
rect 443052 271215 443054 271224
rect 503626 271280 503682 271289
rect 503626 271215 503628 271224
rect 443000 271186 443052 271192
rect 503680 271215 503682 271224
rect 503628 271186 503680 271192
rect 516612 271182 516640 378286
rect 517532 358834 517560 466482
rect 517612 378276 517664 378282
rect 517612 378218 517664 378224
rect 517520 358828 517572 358834
rect 517520 358770 517572 358776
rect 440148 271176 440200 271182
rect 433338 271144 433394 271153
rect 440148 271118 440200 271124
rect 516600 271176 516652 271182
rect 516600 271118 516652 271124
rect 433338 271079 433394 271088
rect 427082 271008 427138 271017
rect 427082 270943 427138 270952
rect 429198 271008 429254 271017
rect 429198 270943 429254 270952
rect 425702 270736 425758 270745
rect 425702 270671 425758 270680
rect 425716 252006 425744 270671
rect 425704 252000 425756 252006
rect 425704 251942 425756 251948
rect 421564 251932 421616 251938
rect 421564 251874 421616 251880
rect 427096 251870 427124 270943
rect 429212 252414 429240 270943
rect 433352 269006 433380 271079
rect 434718 271008 434774 271017
rect 434718 270943 434774 270952
rect 436098 271008 436154 271017
rect 436098 270943 436154 270952
rect 433340 269000 433392 269006
rect 433340 268942 433392 268948
rect 434732 252482 434760 270943
rect 436112 252550 436140 270943
rect 436190 270600 436246 270609
rect 436190 270535 436246 270544
rect 436204 269074 436232 270535
rect 436192 269068 436244 269074
rect 436192 269010 436244 269016
rect 500868 253360 500920 253366
rect 500866 253328 500868 253337
rect 500920 253328 500922 253337
rect 499212 253292 499264 253298
rect 500866 253263 500922 253272
rect 499212 253234 499264 253240
rect 499224 252793 499252 253234
rect 499210 252784 499266 252793
rect 499210 252719 499266 252728
rect 510894 252648 510950 252657
rect 510894 252583 510896 252592
rect 510948 252583 510950 252592
rect 510896 252554 510948 252560
rect 436100 252544 436152 252550
rect 436100 252486 436152 252492
rect 434720 252476 434772 252482
rect 434720 252418 434772 252424
rect 429200 252408 429252 252414
rect 429200 252350 429252 252356
rect 427084 251864 427136 251870
rect 396722 251832 396778 251841
rect 427084 251806 427136 251812
rect 396722 251767 396778 251776
rect 423404 167000 423456 167006
rect 423404 166942 423456 166948
rect 418436 166932 418488 166938
rect 418436 166874 418488 166880
rect 418448 166841 418476 166874
rect 421012 166864 421064 166870
rect 418434 166832 418490 166841
rect 418434 166767 418490 166776
rect 421010 166832 421012 166841
rect 423416 166841 423444 166942
rect 421064 166832 421066 166841
rect 421010 166767 421066 166776
rect 423402 166832 423458 166841
rect 423402 166767 423458 166776
rect 445850 166832 445906 166841
rect 445850 166767 445852 166776
rect 445904 166767 445906 166776
rect 470966 166832 471022 166841
rect 470966 166767 471022 166776
rect 473450 166832 473506 166841
rect 473450 166767 473506 166776
rect 475842 166832 475898 166841
rect 475842 166767 475898 166776
rect 478418 166832 478474 166841
rect 478418 166767 478474 166776
rect 480902 166832 480958 166841
rect 480902 166767 480958 166776
rect 445852 166738 445904 166744
rect 470980 166734 471008 166767
rect 470968 166728 471020 166734
rect 470968 166670 471020 166676
rect 473464 166598 473492 166767
rect 475856 166666 475884 166767
rect 475844 166660 475896 166666
rect 475844 166602 475896 166608
rect 473452 166592 473504 166598
rect 473452 166534 473504 166540
rect 478432 166462 478460 166767
rect 480916 166530 480944 166767
rect 483386 166696 483442 166705
rect 483386 166631 483442 166640
rect 485962 166696 486018 166705
rect 485962 166631 486018 166640
rect 480904 166524 480956 166530
rect 480904 166466 480956 166472
rect 478420 166456 478472 166462
rect 478420 166398 478472 166404
rect 483400 166394 483428 166631
rect 483388 166388 483440 166394
rect 483388 166330 483440 166336
rect 485976 166326 486004 166631
rect 503258 166560 503314 166569
rect 503258 166495 503314 166504
rect 485964 166320 486016 166326
rect 428186 166288 428242 166297
rect 428186 166223 428242 166232
rect 430946 166288 431002 166297
rect 485964 166262 486016 166268
rect 430946 166223 430948 166232
rect 428200 166190 428228 166223
rect 431000 166223 431002 166232
rect 430948 166194 431000 166200
rect 428188 166184 428240 166190
rect 428188 166126 428240 166132
rect 433340 165640 433392 165646
rect 397458 165608 397514 165617
rect 397458 165543 397514 165552
rect 401598 165608 401654 165617
rect 401598 165543 401654 165552
rect 404358 165608 404414 165617
rect 404358 165543 404414 165552
rect 407118 165608 407174 165617
rect 407118 165543 407174 165552
rect 409878 165608 409934 165617
rect 409878 165543 409934 165552
rect 415398 165608 415454 165617
rect 415398 165543 415454 165552
rect 416042 165608 416098 165617
rect 416042 165543 416098 165552
rect 418618 165608 418674 165617
rect 418618 165543 418674 165552
rect 423678 165608 423734 165617
rect 423678 165543 423734 165552
rect 427634 165608 427690 165617
rect 427634 165543 427690 165552
rect 433338 165608 433340 165617
rect 433392 165608 433394 165617
rect 433338 165543 433394 165552
rect 433522 165608 433578 165617
rect 433522 165543 433578 165552
rect 434718 165608 434774 165617
rect 434718 165543 434774 165552
rect 437754 165608 437810 165617
rect 437754 165543 437810 165552
rect 438030 165608 438086 165617
rect 438030 165543 438086 165552
rect 442998 165608 443054 165617
rect 442998 165543 443054 165552
rect 447322 165608 447378 165617
rect 447322 165543 447378 165552
rect 449898 165608 449954 165617
rect 449898 165543 449954 165552
rect 452658 165608 452714 165617
rect 452658 165543 452714 165552
rect 455418 165608 455474 165617
rect 455418 165543 455474 165552
rect 458362 165608 458418 165617
rect 458362 165543 458364 165552
rect 396078 164384 396134 164393
rect 396078 164319 396134 164328
rect 396092 164014 396120 164319
rect 396170 164248 396226 164257
rect 396170 164183 396226 164192
rect 396184 164082 396212 164183
rect 396172 164076 396224 164082
rect 396172 164018 396224 164024
rect 396080 164008 396132 164014
rect 396080 163950 396132 163956
rect 379980 162852 380032 162858
rect 379980 162794 380032 162800
rect 379992 162586 380020 162794
rect 379980 162580 380032 162586
rect 379980 162522 380032 162528
rect 379980 148368 380032 148374
rect 379980 148310 380032 148316
rect 379888 145376 379940 145382
rect 379888 145318 379940 145324
rect 379796 59288 379848 59294
rect 379796 59230 379848 59236
rect 379704 56228 379756 56234
rect 379704 56170 379756 56176
rect 379900 56166 379928 145318
rect 379888 56160 379940 56166
rect 379888 56102 379940 56108
rect 379336 56092 379388 56098
rect 379336 56034 379388 56040
rect 378784 55956 378836 55962
rect 378784 55898 378836 55904
rect 379992 54942 380020 148310
rect 396092 145450 396120 163950
rect 396184 145518 396212 164018
rect 396724 161492 396776 161498
rect 396724 161434 396776 161440
rect 396736 146198 396764 161434
rect 397472 148578 397500 165543
rect 398838 164248 398894 164257
rect 398838 164183 398894 164192
rect 400218 164248 400274 164257
rect 400218 164183 400274 164192
rect 398852 148646 398880 164183
rect 398840 148640 398892 148646
rect 398840 148582 398892 148588
rect 397460 148572 397512 148578
rect 397460 148514 397512 148520
rect 400232 148510 400260 164183
rect 400220 148504 400272 148510
rect 400220 148446 400272 148452
rect 401612 148442 401640 165543
rect 402978 164384 403034 164393
rect 402978 164319 403034 164328
rect 401600 148436 401652 148442
rect 401600 148378 401652 148384
rect 396724 146192 396776 146198
rect 396724 146134 396776 146140
rect 402992 145722 403020 164319
rect 403070 164248 403126 164257
rect 403070 164183 403126 164192
rect 403084 145790 403112 164183
rect 404372 146266 404400 165543
rect 407132 164694 407160 165543
rect 409892 164830 409920 165543
rect 409880 164824 409932 164830
rect 409880 164766 409932 164772
rect 412638 164792 412694 164801
rect 412638 164727 412640 164736
rect 412692 164727 412694 164736
rect 412640 164698 412692 164704
rect 407120 164688 407172 164694
rect 407120 164630 407172 164636
rect 411350 164384 411406 164393
rect 411350 164319 411406 164328
rect 405738 164248 405794 164257
rect 405738 164183 405794 164192
rect 407210 164248 407266 164257
rect 407210 164183 407266 164192
rect 408498 164248 408554 164257
rect 408498 164183 408554 164192
rect 409970 164248 410026 164257
rect 409970 164183 410026 164192
rect 411258 164248 411314 164257
rect 411258 164183 411314 164192
rect 404360 146260 404412 146266
rect 404360 146202 404412 146208
rect 405752 145858 405780 164183
rect 407224 145926 407252 164183
rect 407212 145920 407264 145926
rect 407212 145862 407264 145868
rect 405740 145852 405792 145858
rect 405740 145794 405792 145800
rect 403072 145784 403124 145790
rect 403072 145726 403124 145732
rect 402980 145716 403032 145722
rect 402980 145658 403032 145664
rect 408512 145654 408540 164183
rect 409984 145994 410012 164183
rect 411272 146062 411300 164183
rect 411260 146056 411312 146062
rect 411260 145998 411312 146004
rect 409972 145988 410024 145994
rect 409972 145930 410024 145936
rect 408500 145648 408552 145654
rect 408500 145590 408552 145596
rect 396172 145512 396224 145518
rect 396172 145454 396224 145460
rect 396080 145444 396132 145450
rect 396080 145386 396132 145392
rect 411364 145314 411392 164319
rect 412730 164248 412786 164257
rect 412730 164183 412786 164192
rect 414018 164248 414074 164257
rect 414018 164183 414074 164192
rect 412744 146130 412772 164183
rect 412732 146124 412784 146130
rect 412732 146066 412784 146072
rect 414032 145382 414060 164183
rect 415412 145897 415440 165543
rect 416056 164898 416084 165543
rect 416044 164892 416096 164898
rect 416044 164834 416096 164840
rect 416778 164248 416834 164257
rect 416778 164183 416834 164192
rect 418158 164248 418214 164257
rect 418158 164183 418214 164192
rect 416792 146198 416820 164183
rect 418172 162314 418200 164183
rect 418632 162722 418660 165543
rect 420918 164792 420974 164801
rect 420918 164727 420974 164736
rect 419538 164248 419594 164257
rect 419538 164183 419594 164192
rect 418620 162716 418672 162722
rect 418620 162658 418672 162664
rect 419552 162654 419580 164183
rect 420932 162790 420960 164727
rect 422298 164248 422354 164257
rect 422298 164183 422354 164192
rect 422312 163674 422340 164183
rect 422300 163668 422352 163674
rect 422300 163610 422352 163616
rect 420920 162784 420972 162790
rect 420920 162726 420972 162732
rect 419540 162648 419592 162654
rect 419540 162590 419592 162596
rect 418160 162308 418212 162314
rect 418160 162250 418212 162256
rect 416780 146192 416832 146198
rect 416780 146134 416832 146140
rect 415398 145888 415454 145897
rect 415398 145823 415454 145832
rect 423692 145761 423720 165543
rect 426346 164248 426402 164257
rect 426402 164206 426480 164234
rect 426346 164183 426402 164192
rect 426452 146305 426480 164206
rect 427648 164098 427676 165543
rect 433338 165064 433394 165073
rect 433338 164999 433340 165008
rect 433392 164999 433394 165008
rect 433340 164970 433392 164976
rect 433536 164626 433564 165543
rect 434732 165102 434760 165543
rect 434720 165096 434772 165102
rect 434720 165038 434772 165044
rect 428924 164620 428976 164626
rect 428924 164562 428976 164568
rect 433524 164620 433576 164626
rect 433524 164562 433576 164568
rect 427726 164248 427782 164257
rect 427782 164206 427952 164234
rect 427726 164183 427782 164192
rect 427648 164070 427860 164098
rect 426438 146296 426494 146305
rect 426438 146231 426494 146240
rect 423678 145752 423734 145761
rect 423678 145687 423734 145696
rect 427832 145625 427860 164070
rect 427924 149054 427952 164206
rect 428936 162246 428964 164562
rect 436098 164520 436154 164529
rect 436098 164455 436154 164464
rect 429290 164384 429346 164393
rect 429290 164319 429346 164328
rect 429106 164248 429162 164257
rect 429162 164206 429240 164234
rect 429106 164183 429162 164192
rect 428924 162240 428976 162246
rect 428924 162182 428976 162188
rect 427912 149048 427964 149054
rect 427912 148990 427964 148996
rect 429212 148374 429240 164206
rect 429304 163606 429332 164319
rect 430578 164248 430634 164257
rect 430578 164183 430634 164192
rect 431958 164248 432014 164257
rect 431958 164183 432014 164192
rect 434718 164248 434774 164257
rect 434718 164183 434774 164192
rect 429292 163600 429344 163606
rect 429292 163542 429344 163548
rect 430592 162178 430620 164183
rect 431972 163538 432000 164183
rect 434732 164150 434760 164183
rect 434720 164144 434772 164150
rect 434720 164086 434772 164092
rect 431960 163532 432012 163538
rect 431960 163474 432012 163480
rect 436112 162858 436140 164455
rect 437768 164218 437796 165543
rect 438044 165170 438072 165543
rect 443012 165238 443040 165543
rect 447336 165510 447364 165543
rect 447324 165504 447376 165510
rect 447324 165446 447376 165452
rect 449912 165306 449940 165543
rect 452672 165374 452700 165543
rect 455432 165442 455460 165543
rect 458416 165543 458418 165552
rect 458364 165514 458416 165520
rect 455420 165436 455472 165442
rect 455420 165378 455472 165384
rect 452660 165368 452712 165374
rect 452660 165310 452712 165316
rect 449900 165300 449952 165306
rect 449900 165242 449952 165248
rect 443000 165232 443052 165238
rect 443000 165174 443052 165180
rect 503272 165170 503300 166495
rect 503350 165608 503406 165617
rect 503350 165543 503406 165552
rect 438032 165164 438084 165170
rect 438032 165106 438084 165112
rect 503260 165164 503312 165170
rect 503260 165106 503312 165112
rect 440240 165096 440292 165102
rect 440240 165038 440292 165044
rect 440146 164248 440202 164257
rect 437756 164212 437808 164218
rect 440252 164234 440280 165038
rect 503364 165034 503392 165543
rect 516612 165102 516640 271118
rect 517532 252618 517560 358770
rect 517624 271386 517652 378218
rect 517704 378208 517756 378214
rect 517704 378150 517756 378156
rect 517612 271380 517664 271386
rect 517612 271322 517664 271328
rect 517520 252612 517572 252618
rect 517520 252554 517572 252560
rect 516600 165096 516652 165102
rect 516600 165038 516652 165044
rect 503352 165028 503404 165034
rect 503352 164970 503404 164976
rect 517532 164966 517560 252554
rect 517624 165170 517652 271322
rect 517716 271250 517744 378150
rect 517808 364334 517836 466550
rect 517888 466472 517940 466478
rect 517888 466414 517940 466420
rect 517900 383654 517928 466414
rect 518900 465112 518952 465118
rect 518900 465054 518952 465060
rect 518912 459649 518940 465054
rect 518898 459640 518954 459649
rect 518898 459575 518954 459584
rect 519542 459640 519598 459649
rect 519542 459575 519598 459584
rect 518990 400344 519046 400353
rect 518990 400279 519046 400288
rect 517900 383626 518112 383654
rect 517808 364306 518020 364334
rect 517992 359582 518020 364306
rect 518084 359718 518112 383626
rect 519004 370530 519032 400279
rect 519082 398168 519138 398177
rect 519082 398103 519138 398112
rect 518992 370524 519044 370530
rect 518992 370466 519044 370472
rect 518900 365016 518952 365022
rect 518900 364958 518952 364964
rect 518072 359712 518124 359718
rect 518072 359654 518124 359660
rect 517980 359576 518032 359582
rect 517980 359518 518032 359524
rect 517704 271244 517756 271250
rect 517704 271186 517756 271192
rect 517716 267734 517744 271186
rect 517716 267706 517928 267734
rect 517796 253360 517848 253366
rect 517796 253302 517848 253308
rect 517704 253292 517756 253298
rect 517704 253234 517756 253240
rect 517612 165164 517664 165170
rect 517612 165106 517664 165112
rect 510528 164960 510580 164966
rect 440330 164928 440386 164937
rect 510528 164902 510580 164908
rect 517520 164960 517572 164966
rect 517520 164902 517572 164908
rect 440330 164863 440386 164872
rect 440344 164830 440372 164863
rect 440332 164824 440384 164830
rect 440332 164766 440384 164772
rect 440202 164206 440280 164234
rect 440146 164183 440202 164192
rect 437756 164154 437808 164160
rect 436100 162852 436152 162858
rect 436100 162794 436152 162800
rect 430580 162172 430632 162178
rect 430580 162114 430632 162120
rect 429200 148368 429252 148374
rect 429200 148310 429252 148316
rect 427818 145616 427874 145625
rect 427818 145551 427874 145560
rect 414020 145376 414072 145382
rect 414020 145318 414072 145324
rect 411352 145308 411404 145314
rect 411352 145250 411404 145256
rect 440252 144129 440280 164206
rect 500224 146192 500276 146198
rect 500224 146134 500276 146140
rect 498660 146124 498712 146130
rect 498660 146066 498712 146072
rect 498672 144945 498700 146066
rect 500236 144945 500264 146134
rect 510540 145586 510568 164902
rect 517520 146192 517572 146198
rect 517520 146134 517572 146140
rect 517532 145654 517560 146134
rect 517520 145648 517572 145654
rect 517520 145590 517572 145596
rect 510528 145580 510580 145586
rect 510528 145522 510580 145528
rect 510540 145466 510568 145522
rect 510618 145480 510674 145489
rect 510540 145438 510618 145466
rect 510618 145415 510674 145424
rect 498658 144936 498714 144945
rect 498658 144871 498714 144880
rect 500222 144936 500278 144945
rect 500222 144871 500278 144880
rect 440238 144120 440294 144129
rect 440238 144055 440294 144064
rect 396078 59800 396134 59809
rect 396078 59735 396080 59744
rect 396132 59735 396134 59744
rect 397090 59800 397146 59809
rect 397090 59735 397146 59744
rect 416042 59800 416098 59809
rect 416042 59735 416098 59744
rect 416962 59800 417018 59809
rect 416962 59735 417018 59744
rect 422850 59800 422906 59809
rect 422850 59735 422906 59744
rect 423954 59800 424010 59809
rect 423954 59735 424010 59744
rect 396080 59706 396132 59712
rect 397104 59702 397132 59735
rect 397092 59696 397144 59702
rect 397092 59638 397144 59644
rect 403070 59664 403126 59673
rect 403070 59599 403126 59608
rect 404174 59664 404230 59673
rect 404174 59599 404230 59608
rect 412546 59664 412602 59673
rect 412546 59599 412602 59608
rect 403084 59362 403112 59599
rect 403072 59356 403124 59362
rect 403072 59298 403124 59304
rect 404188 59226 404216 59599
rect 404176 59220 404228 59226
rect 404176 59162 404228 59168
rect 398194 57896 398250 57905
rect 398194 57831 398250 57840
rect 398838 57896 398894 57905
rect 398838 57831 398894 57840
rect 400402 57896 400458 57905
rect 400402 57831 400458 57840
rect 401598 57896 401654 57905
rect 401598 57831 401654 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407210 57896 407266 57905
rect 407210 57831 407266 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 398208 56574 398236 57831
rect 398196 56568 398248 56574
rect 398196 56510 398248 56516
rect 398852 55146 398880 57831
rect 400416 55894 400444 57831
rect 400404 55888 400456 55894
rect 400404 55830 400456 55836
rect 398840 55140 398892 55146
rect 398840 55082 398892 55088
rect 379980 54936 380032 54942
rect 379980 54878 380032 54884
rect 378048 54868 378100 54874
rect 378048 54810 378100 54816
rect 377864 54800 377916 54806
rect 377864 54742 377916 54748
rect 376484 54732 376536 54738
rect 376484 54674 376536 54680
rect 375932 54596 375984 54602
rect 375932 54538 375984 54544
rect 401612 54534 401640 57831
rect 404372 54602 404400 57831
rect 405844 54670 405872 57831
rect 407224 54738 407252 57831
rect 408328 55826 408356 57831
rect 408696 55962 408724 57831
rect 408684 55956 408736 55962
rect 408684 55898 408736 55904
rect 408316 55820 408368 55826
rect 408316 55762 408368 55768
rect 409892 54806 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 56030 411300 56879
rect 411260 56024 411312 56030
rect 411260 55966 411312 55972
rect 411364 54874 411392 57831
rect 412560 56953 412588 59599
rect 416056 59430 416084 59735
rect 416976 59634 417004 59735
rect 416964 59628 417016 59634
rect 416964 59570 417016 59576
rect 422864 59566 422892 59735
rect 423494 59664 423550 59673
rect 423494 59599 423550 59608
rect 422852 59560 422904 59566
rect 422852 59502 422904 59508
rect 416044 59424 416096 59430
rect 416044 59366 416096 59372
rect 418158 59392 418214 59401
rect 418158 59327 418214 59336
rect 419354 59392 419410 59401
rect 419354 59327 419410 59336
rect 420642 59392 420698 59401
rect 420642 59327 420698 59336
rect 421746 59392 421802 59401
rect 421746 59327 421802 59336
rect 418172 59294 418200 59327
rect 418160 59288 418212 59294
rect 418160 59230 418212 59236
rect 419368 59158 419396 59327
rect 419356 59152 419408 59158
rect 419356 59094 419408 59100
rect 420656 59090 420684 59327
rect 420644 59084 420696 59090
rect 420644 59026 420696 59032
rect 421760 59022 421788 59327
rect 421748 59016 421800 59022
rect 421748 58958 421800 58964
rect 423508 58954 423536 59599
rect 423968 59498 423996 59735
rect 423956 59492 424008 59498
rect 423956 59434 424008 59440
rect 425978 59392 426034 59401
rect 425978 59327 426034 59336
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 453394 59392 453450 59401
rect 453394 59327 453450 59336
rect 423496 58948 423548 58954
rect 423496 58890 423548 58896
rect 425992 58886 426020 59327
rect 425980 58880 426032 58886
rect 425980 58822 426032 58828
rect 428200 58682 428228 59327
rect 453408 58818 453436 59327
rect 475842 58984 475898 58993
rect 475842 58919 475898 58928
rect 453396 58812 453448 58818
rect 453396 58754 453448 58760
rect 475856 58750 475884 58919
rect 475844 58744 475896 58750
rect 475844 58686 475896 58692
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 517624 57934 517652 165106
rect 517716 146130 517744 253234
rect 517808 253230 517836 253302
rect 517796 253224 517848 253230
rect 517796 253166 517848 253172
rect 517808 146198 517836 253166
rect 517900 165034 517928 267706
rect 517992 253298 518020 359518
rect 517980 253292 518032 253298
rect 517980 253234 518032 253240
rect 518084 253230 518112 359654
rect 518912 292505 518940 364958
rect 519004 293865 519032 370466
rect 519096 365022 519124 398103
rect 519266 396808 519322 396817
rect 519266 396743 519322 396752
rect 519174 395312 519230 395321
rect 519174 395247 519230 395256
rect 519084 365016 519136 365022
rect 519084 364958 519136 364964
rect 519188 363662 519216 395247
rect 519280 366382 519308 396743
rect 519358 394088 519414 394097
rect 519358 394023 519414 394032
rect 519372 383654 519400 394023
rect 519372 383626 519492 383654
rect 519268 366376 519320 366382
rect 519268 366318 519320 366324
rect 519176 363656 519228 363662
rect 519176 363598 519228 363604
rect 518990 293856 519046 293865
rect 518990 293791 519046 293800
rect 518898 292496 518954 292505
rect 518898 292431 518954 292440
rect 519082 290320 519138 290329
rect 519082 290255 519138 290264
rect 518990 287600 519046 287609
rect 518990 287535 519046 287544
rect 519004 287094 519032 287535
rect 518992 287088 519044 287094
rect 518992 287030 519044 287036
rect 518072 253224 518124 253230
rect 518072 253166 518124 253172
rect 518898 186416 518954 186425
rect 518898 186351 518954 186360
rect 517888 165028 517940 165034
rect 517888 164970 517940 164976
rect 517796 146192 517848 146198
rect 517796 146134 517848 146140
rect 517704 146124 517756 146130
rect 517704 146066 517756 146072
rect 517716 145586 517744 146066
rect 517704 145580 517756 145586
rect 517704 145522 517756 145528
rect 478420 57928 478472 57934
rect 414570 57896 414626 57905
rect 414570 57831 414626 57840
rect 415490 57896 415546 57905
rect 415490 57831 415546 57840
rect 418434 57896 418490 57905
rect 418434 57831 418490 57840
rect 425058 57896 425114 57905
rect 425058 57831 425114 57840
rect 426438 57896 426494 57905
rect 426438 57831 426494 57840
rect 427634 57896 427690 57905
rect 427634 57831 427690 57840
rect 427818 57896 427874 57905
rect 427818 57831 427874 57840
rect 429198 57896 429254 57905
rect 429198 57831 429254 57840
rect 431130 57896 431186 57905
rect 431130 57831 431186 57840
rect 431958 57896 432014 57905
rect 431958 57831 432014 57840
rect 433338 57896 433394 57905
rect 433338 57831 433394 57840
rect 433522 57896 433578 57905
rect 433522 57831 433578 57840
rect 435730 57896 435786 57905
rect 435730 57831 435786 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 443458 57896 443514 57905
rect 443458 57831 443514 57840
rect 445850 57896 445906 57905
rect 445850 57831 445906 57840
rect 448242 57896 448298 57905
rect 448242 57831 448298 57840
rect 465906 57896 465962 57905
rect 465906 57831 465962 57840
rect 478418 57896 478420 57905
rect 503260 57928 503312 57934
rect 478472 57896 478474 57905
rect 478418 57831 478474 57840
rect 485962 57896 486018 57905
rect 485962 57831 485964 57840
rect 412546 56944 412602 56953
rect 412546 56879 412602 56888
rect 412638 56808 412694 56817
rect 412638 56743 412694 56752
rect 412652 56098 412680 56743
rect 414584 56166 414612 57831
rect 415504 57254 415532 57831
rect 418448 57322 418476 57831
rect 418436 57316 418488 57322
rect 418436 57258 418488 57264
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 414572 56160 414624 56166
rect 414572 56102 414624 56108
rect 412640 56092 412692 56098
rect 412640 56034 412692 56040
rect 425072 55049 425100 57831
rect 426452 56234 426480 57831
rect 427648 56302 427676 57831
rect 427636 56296 427688 56302
rect 427636 56238 427688 56244
rect 426440 56228 426492 56234
rect 426440 56170 426492 56176
rect 425058 55040 425114 55049
rect 425058 54975 425114 54984
rect 427832 54942 427860 57831
rect 429212 55010 429240 57831
rect 431144 56370 431172 57831
rect 431132 56364 431184 56370
rect 431132 56306 431184 56312
rect 431972 55078 432000 57831
rect 433246 57624 433302 57633
rect 433246 57559 433302 57568
rect 433260 57225 433288 57559
rect 433246 57216 433302 57225
rect 433246 57151 433302 57160
rect 433352 56438 433380 57831
rect 433430 57624 433486 57633
rect 433430 57559 433486 57568
rect 433340 56432 433392 56438
rect 433340 56374 433392 56380
rect 431960 55072 432012 55078
rect 431960 55014 432012 55020
rect 429200 55004 429252 55010
rect 429200 54946 429252 54952
rect 427820 54936 427872 54942
rect 427820 54878 427872 54884
rect 411352 54868 411404 54874
rect 411352 54810 411404 54816
rect 409880 54800 409932 54806
rect 409880 54742 409932 54748
rect 407212 54732 407264 54738
rect 407212 54674 407264 54680
rect 405832 54664 405884 54670
rect 405832 54606 405884 54612
rect 404360 54596 404412 54602
rect 404360 54538 404412 54544
rect 401600 54528 401652 54534
rect 401600 54470 401652 54476
rect 433444 54466 433472 57559
rect 433536 57390 433564 57831
rect 433524 57384 433576 57390
rect 433524 57326 433576 57332
rect 435744 56506 435772 57831
rect 435928 57526 435956 57831
rect 436098 57624 436154 57633
rect 436098 57559 436154 57568
rect 435916 57520 435968 57526
rect 435916 57462 435968 57468
rect 435732 56500 435784 56506
rect 435732 56442 435784 56448
rect 436112 55214 436140 57559
rect 438504 57458 438532 57831
rect 438858 57624 438914 57633
rect 443472 57594 443500 57831
rect 445864 57730 445892 57831
rect 445852 57724 445904 57730
rect 445852 57666 445904 57672
rect 448256 57662 448284 57831
rect 465920 57798 465948 57831
rect 486016 57831 486018 57840
rect 503258 57896 503260 57905
rect 517612 57928 517664 57934
rect 503312 57896 503314 57905
rect 503258 57831 503314 57840
rect 503534 57896 503590 57905
rect 517612 57870 517664 57876
rect 517900 57866 517928 164970
rect 518912 79937 518940 186351
rect 519004 180713 519032 287030
rect 519096 183433 519124 290255
rect 519188 288833 519216 363598
rect 519464 362234 519492 383626
rect 519452 362228 519504 362234
rect 519452 362170 519504 362176
rect 519266 352880 519322 352889
rect 519266 352815 519322 352824
rect 519174 288824 519230 288833
rect 519174 288759 519230 288768
rect 519082 183424 519138 183433
rect 519082 183359 519138 183368
rect 518990 180704 519046 180713
rect 518990 180639 519046 180648
rect 518898 79928 518954 79937
rect 518898 79863 518954 79872
rect 519004 74225 519032 180639
rect 519096 76809 519124 183359
rect 519188 181937 519216 288759
rect 519280 246265 519308 352815
rect 519358 293856 519414 293865
rect 519358 293791 519414 293800
rect 519266 246256 519322 246265
rect 519266 246191 519322 246200
rect 519174 181928 519230 181937
rect 519174 181863 519230 181872
rect 519280 139369 519308 246191
rect 519372 186425 519400 293791
rect 519464 287094 519492 362170
rect 519556 352889 519584 459575
rect 520936 396778 520964 495450
rect 578896 404977 578924 523670
rect 580264 515432 580316 515438
rect 580264 515374 580316 515380
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580276 458153 580304 515374
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 578882 404968 578938 404977
rect 578882 404903 578938 404912
rect 520924 396772 520976 396778
rect 520924 396714 520976 396720
rect 580356 396772 580408 396778
rect 580356 396714 580408 396720
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580264 378276 580316 378282
rect 580264 378218 580316 378224
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 519636 366376 519688 366382
rect 519636 366318 519688 366324
rect 519542 352880 519598 352889
rect 519542 352815 519598 352824
rect 519542 292496 519598 292505
rect 519542 292431 519598 292440
rect 519452 287088 519504 287094
rect 519452 287030 519504 287036
rect 519358 186416 519414 186425
rect 519358 186351 519414 186360
rect 519556 184793 519584 292431
rect 519648 290329 519676 366318
rect 580276 325281 580304 378218
rect 580368 351937 580396 396714
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 519634 290320 519690 290329
rect 519634 290255 519690 290264
rect 520186 288824 520242 288833
rect 520186 288759 520242 288768
rect 520200 288454 520228 288759
rect 520188 288448 520240 288454
rect 520188 288390 520240 288396
rect 580264 288448 580316 288454
rect 580264 288390 580316 288396
rect 580276 232393 580304 288390
rect 580356 287088 580408 287094
rect 580356 287030 580408 287036
rect 580368 272241 580396 287030
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 519542 184784 519598 184793
rect 519542 184719 519598 184728
rect 520186 184784 520242 184793
rect 520186 184719 520242 184728
rect 520200 183598 520228 184719
rect 519452 183592 519504 183598
rect 519452 183534 519504 183540
rect 520188 183592 520240 183598
rect 520188 183534 520240 183540
rect 580264 183592 580316 183598
rect 580264 183534 580316 183540
rect 519358 181928 519414 181937
rect 519358 181863 519414 181872
rect 519266 139360 519322 139369
rect 519266 139295 519322 139304
rect 519082 76800 519138 76809
rect 519082 76735 519138 76744
rect 519372 75449 519400 181863
rect 519464 78305 519492 183534
rect 520096 183524 520148 183530
rect 520096 183466 520148 183472
rect 520108 183433 520136 183466
rect 520094 183424 520150 183433
rect 520094 183359 520150 183368
rect 580276 152697 580304 183534
rect 580368 183530 580396 192471
rect 580356 183524 580408 183530
rect 580356 183466 580408 183472
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580264 145648 580316 145654
rect 580264 145590 580316 145596
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519450 78296 519506 78305
rect 519450 78231 519506 78240
rect 519358 75440 519414 75449
rect 519358 75375 519414 75384
rect 518990 74216 519046 74225
rect 518990 74151 519046 74160
rect 503534 57831 503536 57840
rect 485964 57802 486016 57808
rect 503588 57831 503590 57840
rect 517888 57860 517940 57866
rect 503536 57802 503588 57808
rect 517888 57802 517940 57808
rect 465908 57792 465960 57798
rect 465908 57734 465960 57740
rect 448244 57656 448296 57662
rect 448244 57598 448296 57604
rect 438858 57559 438914 57568
rect 443460 57588 443512 57594
rect 438492 57452 438544 57458
rect 438492 57394 438544 57400
rect 436100 55208 436152 55214
rect 438872 55185 438900 57559
rect 443460 57530 443512 57536
rect 436100 55150 436152 55156
rect 438858 55176 438914 55185
rect 438858 55111 438914 55120
rect 242900 54460 242952 54466
rect 242900 54402 242952 54408
rect 373724 54460 373776 54466
rect 373724 54402 373776 54408
rect 433432 54460 433484 54466
rect 433432 54402 433484 54408
rect 213644 54324 213696 54330
rect 213644 54266 213696 54272
rect 240140 54324 240192 54330
rect 240140 54266 240192 54272
rect 580276 33153 580304 145590
rect 580356 145580 580408 145586
rect 580356 145522 580408 145528
rect 580368 73001 580396 145522
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 140042 4040 140098 4049
rect 140042 3975 140098 3984
rect 129370 3904 129426 3913
rect 129370 3839 129426 3848
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 584 480 612 3402
rect 125876 2848 125928 2854
rect 125876 2790 125928 2796
rect 125888 480 125916 2790
rect 129384 480 129412 3839
rect 132958 3360 133014 3369
rect 132958 3295 133014 3304
rect 132972 480 133000 3295
rect 136454 3224 136510 3233
rect 136454 3159 136510 3168
rect 136468 480 136496 3159
rect 140056 480 140084 3975
rect 147126 3768 147182 3777
rect 147126 3703 147182 3712
rect 143538 3632 143594 3641
rect 143538 3567 143594 3576
rect 143552 480 143580 3567
rect 147140 480 147168 3703
rect 150622 3496 150678 3505
rect 150622 3431 150678 3440
rect 150636 480 150664 3431
rect 367098 2952 367154 2961
rect 367098 2887 367154 2896
rect 367112 2854 367140 2887
rect 367100 2848 367152 2854
rect 367100 2790 367152 2796
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 579944 3478 580000
rect 3422 547848 3478 547904
rect 3422 514800 3478 514856
rect 2962 410488 3018 410544
rect 3330 358400 3386 358456
rect 3238 97552 3294 97608
rect 3514 482160 3570 482216
rect 3606 462576 3662 462632
rect 57702 622376 57758 622432
rect 57518 619656 57574 619712
rect 57242 595176 57298 595232
rect 57150 589056 57206 589112
rect 57058 576816 57114 576872
rect 57426 591776 57482 591832
rect 57334 579672 57390 579728
rect 57610 613536 57666 613592
rect 58990 628632 59046 628688
rect 58622 616256 58678 616312
rect 57886 604016 57942 604072
rect 58530 585656 58586 585712
rect 58438 573416 58494 573472
rect 58898 610136 58954 610192
rect 58806 601296 58862 601352
rect 58714 597896 58770 597952
rect 59174 625776 59230 625832
rect 59082 607552 59138 607608
rect 59082 582936 59138 582992
rect 59542 570732 59598 570788
rect 120814 608912 120870 608968
rect 121090 591164 121146 591220
rect 121182 572804 121238 572860
rect 121550 625232 121606 625288
rect 121826 621152 121882 621208
rect 121734 615576 121790 615632
rect 121918 618432 121974 618488
rect 122010 600344 122066 600400
rect 122102 587968 122158 588024
rect 122194 581712 122250 581768
rect 122286 578312 122342 578368
rect 122930 627952 122986 628008
rect 123114 612720 123170 612776
rect 123298 606192 123354 606248
rect 123206 603064 123262 603120
rect 124126 596672 124182 596728
rect 123390 593952 123446 594008
rect 123482 584432 123538 584488
rect 123666 575592 123722 575648
rect 123574 570016 123630 570072
rect 137282 628632 137338 628688
rect 136730 616256 136786 616312
rect 136730 597896 136786 597952
rect 136730 585656 136786 585712
rect 136730 582936 136786 582992
rect 137190 573416 137246 573472
rect 137558 619656 137614 619712
rect 137374 595176 137430 595232
rect 137466 579672 137522 579728
rect 280986 640328 281042 640384
rect 137742 607552 137798 607608
rect 137742 591776 137798 591832
rect 139030 625776 139086 625832
rect 138938 613536 138994 613592
rect 138846 610136 138902 610192
rect 137926 604016 137982 604072
rect 137926 601296 137982 601352
rect 138754 589056 138810 589112
rect 138662 576816 138718 576872
rect 139306 622376 139362 622432
rect 139214 570696 139270 570752
rect 200762 618432 200818 618488
rect 201038 594564 201094 594620
rect 201498 584432 201554 584488
rect 201130 576204 201186 576260
rect 201222 570084 201278 570140
rect 201774 627952 201830 628008
rect 202970 625232 203026 625288
rect 202234 621152 202290 621208
rect 201866 612720 201922 612776
rect 201958 608912 202014 608968
rect 202050 600344 202106 600400
rect 202142 590688 202198 590744
rect 202878 615576 202934 615632
rect 202326 578312 202382 578368
rect 203154 606328 203210 606384
rect 203062 603064 203118 603120
rect 203246 596692 203302 596728
rect 203246 596672 203248 596692
rect 203248 596672 203300 596692
rect 203300 596672 203302 596692
rect 203246 587968 203302 588024
rect 203338 581712 203394 581768
rect 203430 572736 203486 572792
rect 215942 628632 215998 628688
rect 216678 625776 216734 625832
rect 216678 619676 216734 619712
rect 216678 619656 216680 619676
rect 216680 619656 216732 619676
rect 216732 619656 216734 619676
rect 216678 616256 216734 616312
rect 216678 597896 216734 597952
rect 216678 595176 216734 595232
rect 216678 591776 216734 591832
rect 216034 585656 216090 585712
rect 216678 582936 216734 582992
rect 216678 579692 216734 579728
rect 216678 579672 216680 579692
rect 216680 579672 216732 579692
rect 216732 579672 216734 579692
rect 216678 570696 216734 570752
rect 217690 622376 217746 622432
rect 217414 601296 217470 601352
rect 217598 589056 217654 589112
rect 217506 573416 217562 573472
rect 217782 610136 217838 610192
rect 218702 604152 218758 604208
rect 219254 613536 219310 613592
rect 219162 607552 219218 607608
rect 219162 576816 219218 576872
rect 241518 550024 241574 550080
rect 248694 549888 248750 549944
rect 255134 549616 255190 549672
rect 258722 549752 258778 549808
rect 280894 600344 280950 600400
rect 281538 627952 281594 628008
rect 281170 572804 281226 572860
rect 281078 570016 281134 570072
rect 282918 625232 282974 625288
rect 281630 618432 281686 618488
rect 281722 615576 281778 615632
rect 281814 612720 281870 612776
rect 281906 593952 281962 594008
rect 281998 584432 282054 584488
rect 282090 581712 282146 581768
rect 282182 575592 282238 575648
rect 283010 621152 283066 621208
rect 283102 608912 283158 608968
rect 283286 606328 283342 606384
rect 283194 603064 283250 603120
rect 283654 596672 283710 596728
rect 283378 590688 283434 590744
rect 283470 587968 283526 588024
rect 283562 578312 283618 578368
rect 286690 549344 286746 549400
rect 290922 549480 290978 549536
rect 294510 548120 294566 548176
rect 300306 550024 300362 550080
rect 300306 527040 300362 527096
rect 300582 549616 300638 549672
rect 301502 549480 301558 549536
rect 301594 547848 301650 547904
rect 3514 58520 3570 58576
rect 43442 377440 43498 377496
rect 57886 517928 57942 517984
rect 302790 540368 302846 540424
rect 302330 525408 302386 525464
rect 303066 549752 303122 549808
rect 303066 526904 303122 526960
rect 304354 549344 304410 549400
rect 302238 510448 302294 510504
rect 302238 495508 302294 495544
rect 302238 495488 302240 495508
rect 302240 495488 302292 495508
rect 302292 495488 302294 495508
rect 46110 379344 46166 379400
rect 45926 271224 45982 271280
rect 46570 268368 46626 268424
rect 47490 379208 47546 379264
rect 46938 271496 46994 271552
rect 48134 482568 48190 482624
rect 48042 482432 48098 482488
rect 48226 467880 48282 467936
rect 49054 271768 49110 271824
rect 49238 271768 49294 271824
rect 50526 479440 50582 479496
rect 49422 164736 49478 164792
rect 50710 467880 50766 467936
rect 50618 165416 50674 165472
rect 53470 485016 53526 485072
rect 51630 378936 51686 378992
rect 51906 271396 51908 271416
rect 51908 271396 51960 271416
rect 51960 271396 51962 271416
rect 51906 271360 51962 271396
rect 51906 270272 51962 270328
rect 52366 465160 52422 465216
rect 52366 380840 52422 380896
rect 52274 379480 52330 379536
rect 52366 271360 52422 271416
rect 53286 471144 53342 471200
rect 52458 271088 52514 271144
rect 52826 271088 52882 271144
rect 53102 267688 53158 267744
rect 53654 465976 53710 466032
rect 53562 378800 53618 378856
rect 53470 165280 53526 165336
rect 54206 471416 54262 471472
rect 55034 471552 55090 471608
rect 56138 471280 56194 471336
rect 56138 165144 56194 165200
rect 56690 388592 56746 388648
rect 56966 410352 57022 410408
rect 57242 417288 57298 417344
rect 57610 389680 57666 389736
rect 57610 389000 57666 389056
rect 56874 309848 56930 309904
rect 56690 252456 56746 252512
rect 56598 202952 56654 203008
rect 56046 146240 56102 146296
rect 56782 201320 56838 201376
rect 56598 96464 56654 96520
rect 57518 311072 57574 311128
rect 57426 301552 57482 301608
rect 56966 195200 57022 195256
rect 56874 164056 56930 164112
rect 57150 204176 57206 204232
rect 56782 93744 56838 93800
rect 57334 198736 57390 198792
rect 57242 175344 57298 175400
rect 57150 97416 57206 97472
rect 57886 417152 57942 417208
rect 57886 414160 57942 414216
rect 57886 413208 57942 413264
rect 57886 411440 57942 411496
rect 57886 408584 57942 408640
rect 57886 391448 57942 391504
rect 58530 388456 58586 388512
rect 57794 307808 57850 307864
rect 57702 306720 57758 306776
rect 57610 304952 57666 305008
rect 57610 303612 57666 303648
rect 57610 303592 57612 303612
rect 57612 303592 57664 303612
rect 57664 303592 57666 303612
rect 57518 282240 57574 282296
rect 57518 204176 57574 204232
rect 57794 304952 57850 305008
rect 57702 199824 57758 199880
rect 57702 198736 57758 198792
rect 58714 284144 58770 284200
rect 59082 479848 59138 479904
rect 58806 281968 58862 282024
rect 58806 273128 58862 273184
rect 57886 201320 57942 201376
rect 57794 198056 57850 198112
rect 57426 196288 57482 196344
rect 57334 93336 57390 93392
rect 57794 195200 57850 195256
rect 57518 163920 57574 163976
rect 57702 164076 57758 164112
rect 57702 164056 57704 164076
rect 57704 164056 57756 164076
rect 57756 164056 57758 164076
rect 57610 91024 57666 91080
rect 57426 90480 57482 90536
rect 57886 175344 57942 175400
rect 57794 88168 57850 88224
rect 58622 251096 58678 251152
rect 59174 471688 59230 471744
rect 59082 177520 59138 177576
rect 58806 146240 58862 146296
rect 59082 146240 59138 146296
rect 58714 145696 58770 145752
rect 57886 68856 57942 68912
rect 3422 19352 3478 19408
rect 58898 145560 58954 145616
rect 59818 479576 59874 479632
rect 59634 271224 59690 271280
rect 59634 270544 59690 270600
rect 59358 164192 59414 164248
rect 66350 485288 66406 485344
rect 68466 485696 68522 485752
rect 68926 484880 68982 484936
rect 67822 469784 67878 469840
rect 67730 468288 67786 468344
rect 69202 469104 69258 469160
rect 70582 468968 70638 469024
rect 71778 466384 71834 466440
rect 70398 465976 70454 466032
rect 72514 484744 72570 484800
rect 73802 485560 73858 485616
rect 73894 485288 73950 485344
rect 73342 467064 73398 467120
rect 76010 485424 76066 485480
rect 74630 466112 74686 466168
rect 74538 465840 74594 465896
rect 77298 485696 77354 485752
rect 76654 484472 76710 484528
rect 77390 468560 77446 468616
rect 78862 468832 78918 468888
rect 80794 484472 80850 484528
rect 78954 468696 79010 468752
rect 78770 468424 78826 468480
rect 88522 471552 88578 471608
rect 88430 471416 88486 471472
rect 89810 471280 89866 471336
rect 87510 471144 87566 471200
rect 91374 485152 91430 485208
rect 91926 471688 91982 471744
rect 76562 466248 76618 466304
rect 76010 465704 76066 465760
rect 69110 465568 69166 465624
rect 94042 485016 94098 485072
rect 95330 485288 95386 485344
rect 95514 479848 95570 479904
rect 120078 482568 120134 482624
rect 120446 482432 120502 482488
rect 118790 479712 118846 479768
rect 121366 482704 121422 482760
rect 121918 479440 121974 479496
rect 124402 482296 124458 482352
rect 124494 479576 124550 479632
rect 123666 476856 123722 476912
rect 126334 476720 126390 476776
rect 127346 474136 127402 474192
rect 145654 485288 145710 485344
rect 145470 485016 145526 485072
rect 144826 483656 144882 483712
rect 145746 478352 145802 478408
rect 143538 474000 143594 474056
rect 147586 485152 147642 485208
rect 148230 485424 148286 485480
rect 148046 482296 148102 482352
rect 147218 480800 147274 480856
rect 148322 479440 148378 479496
rect 151358 478216 151414 478272
rect 154486 482432 154542 482488
rect 153198 474272 153254 474328
rect 152738 472504 152794 472560
rect 156510 483792 156566 483848
rect 154670 479576 154726 479632
rect 157522 476720 157578 476776
rect 156786 475496 156842 475552
rect 154578 467200 154634 467256
rect 151818 467064 151874 467120
rect 160098 469784 160154 469840
rect 164514 484200 164570 484256
rect 163778 476856 163834 476912
rect 161662 475632 161718 475688
rect 161570 471280 161626 471336
rect 162858 471416 162914 471472
rect 161754 471144 161810 471200
rect 167274 468832 167330 468888
rect 168378 468696 168434 468752
rect 167090 468560 167146 468616
rect 171138 485560 171194 485616
rect 169850 469920 169906 469976
rect 169758 468968 169814 469024
rect 168562 468424 168618 468480
rect 166998 465976 167054 466032
rect 165802 465840 165858 465896
rect 165618 465704 165674 465760
rect 172058 479712 172114 479768
rect 171230 472640 171286 472696
rect 172610 471552 172666 471608
rect 179326 480936 179382 480992
rect 178038 466556 178040 466576
rect 178040 466556 178092 466576
rect 178092 466556 178094 466576
rect 178038 466520 178094 466556
rect 180154 466928 180210 466984
rect 180062 466112 180118 466168
rect 182730 471824 182786 471880
rect 183650 471688 183706 471744
rect 185766 484880 185822 484936
rect 187054 485696 187110 485752
rect 190918 466520 190974 466576
rect 171138 464344 171194 464400
rect 105818 380296 105874 380352
rect 110970 380316 111026 380352
rect 110970 380296 110972 380316
rect 110972 380296 111024 380316
rect 111024 380296 111026 380316
rect 113546 380332 113548 380352
rect 113548 380332 113600 380352
rect 113600 380332 113602 380352
rect 113546 380296 113602 380332
rect 115938 380296 115994 380352
rect 118330 380296 118386 380352
rect 120906 380296 120962 380352
rect 123574 380332 123576 380352
rect 123576 380332 123628 380352
rect 123628 380332 123630 380352
rect 123574 380296 123630 380332
rect 128358 380296 128414 380352
rect 133510 380296 133566 380352
rect 135902 380296 135958 380352
rect 138478 380296 138534 380352
rect 148598 380316 148654 380352
rect 148598 380296 148600 380316
rect 148600 380296 148652 380316
rect 148652 380296 148654 380316
rect 155958 380296 156014 380352
rect 158534 380296 158590 380352
rect 160926 380296 160982 380352
rect 163502 380296 163558 380352
rect 166078 380296 166134 380352
rect 80334 379344 80390 379400
rect 85486 379344 85542 379400
rect 86590 379344 86646 379400
rect 87694 379344 87750 379400
rect 88338 379380 88340 379400
rect 88340 379380 88392 379400
rect 88392 379380 88394 379400
rect 88338 379344 88394 379380
rect 88798 379364 88854 379400
rect 88798 379344 88800 379364
rect 88800 379344 88852 379364
rect 88852 379344 88854 379364
rect 77206 378936 77262 378992
rect 81438 378800 81494 378856
rect 80334 378664 80390 378720
rect 90638 379344 90694 379400
rect 91374 379344 91430 379400
rect 92386 379380 92388 379400
rect 92388 379380 92440 379400
rect 92440 379380 92442 379400
rect 92386 379344 92442 379380
rect 93582 379344 93638 379400
rect 96066 379344 96122 379400
rect 98182 379344 98238 379400
rect 101034 379344 101090 379400
rect 103518 379344 103574 379400
rect 105358 379344 105414 379400
rect 108210 379344 108266 379400
rect 108854 379344 108910 379400
rect 111246 379344 111302 379400
rect 112350 379344 112406 379400
rect 113454 379344 113510 379400
rect 114466 379344 114522 379400
rect 115846 379344 115902 379400
rect 141054 379344 141110 379400
rect 143630 379344 143686 379400
rect 146022 379344 146078 379400
rect 150990 379344 151046 379400
rect 153566 379344 153622 379400
rect 90730 379244 90732 379264
rect 90732 379244 90784 379264
rect 90784 379244 90786 379264
rect 90730 379208 90786 379244
rect 93490 379208 93546 379264
rect 95974 379208 96030 379264
rect 94686 378528 94742 378584
rect 98366 379208 98422 379264
rect 99470 379208 99526 379264
rect 97722 378528 97778 378584
rect 95974 377848 96030 377904
rect 98366 377576 98422 377632
rect 102966 379208 103022 379264
rect 100758 378392 100814 378448
rect 101954 378256 102010 378312
rect 104070 378392 104126 378448
rect 125966 378392 126022 378448
rect 131026 378392 131082 378448
rect 106462 378120 106518 378176
rect 107566 378120 107622 378176
rect 105358 377712 105414 377768
rect 183466 378392 183522 378448
rect 182270 378120 182326 378176
rect 182822 378120 182878 378176
rect 178590 358828 178646 358864
rect 178590 358808 178592 358828
rect 178592 358808 178644 358828
rect 178644 358808 178646 358828
rect 179694 358844 179696 358864
rect 179696 358844 179748 358864
rect 179748 358844 179750 358864
rect 179694 358808 179750 358844
rect 190918 358808 190974 358864
rect 95974 273808 96030 273864
rect 60830 272720 60886 272776
rect 61014 272720 61070 272776
rect 60830 270544 60886 270600
rect 76010 272856 76066 272912
rect 90730 272856 90786 272912
rect 93674 272856 93730 272912
rect 95882 272856 95938 272912
rect 61750 272584 61806 272640
rect 61474 272448 61530 272504
rect 110970 273556 111026 273592
rect 110970 273536 110972 273556
rect 110972 273536 111024 273556
rect 111024 273536 111026 273556
rect 133418 273536 133474 273592
rect 135902 273536 135958 273592
rect 138478 273536 138534 273592
rect 140870 273536 140926 273592
rect 100758 273148 100814 273184
rect 100758 273128 100760 273148
rect 100760 273128 100812 273148
rect 100812 273128 100814 273148
rect 98458 272856 98514 272912
rect 99378 272856 99434 272912
rect 143538 272584 143594 272640
rect 96986 272312 97042 272368
rect 65338 271360 65394 271416
rect 113546 272176 113602 272232
rect 75918 271768 75974 271824
rect 82818 271768 82874 271824
rect 67362 271088 67418 271144
rect 77298 271088 77354 271144
rect 78678 270972 78734 271008
rect 78678 270952 78680 270972
rect 78680 270952 78732 270972
rect 78732 270952 78734 270972
rect 77850 268368 77906 268424
rect 60922 252320 60978 252376
rect 84198 271768 84254 271824
rect 86958 271768 87014 271824
rect 94226 271768 94282 271824
rect 97998 271768 98054 271824
rect 84658 271632 84714 271688
rect 88338 271108 88394 271144
rect 88338 271088 88340 271108
rect 88340 271088 88392 271108
rect 88392 271088 88394 271108
rect 88338 270952 88394 271008
rect 89718 270952 89774 271008
rect 85578 270816 85634 270872
rect 92478 270816 92534 270872
rect 91098 270544 91154 270600
rect 100758 271768 100814 271824
rect 103518 271632 103574 271688
rect 100758 271360 100814 271416
rect 104898 271360 104954 271416
rect 114466 271768 114522 271824
rect 123206 271788 123262 271824
rect 123206 271768 123208 271788
rect 123208 271768 123260 271788
rect 123260 271768 123262 271788
rect 120078 271632 120134 271688
rect 125598 271652 125654 271688
rect 125598 271632 125600 271652
rect 125600 271632 125652 271652
rect 125652 271632 125654 271652
rect 115938 271496 115994 271552
rect 117318 271516 117374 271552
rect 128358 271768 128414 271824
rect 129738 271804 129740 271824
rect 129740 271804 129792 271824
rect 129792 271804 129794 271824
rect 129738 271768 129794 271804
rect 151358 271804 151360 271824
rect 151360 271804 151412 271824
rect 151412 271804 151414 271824
rect 151358 271768 151414 271804
rect 154486 271768 154542 271824
rect 157246 271788 157302 271824
rect 157246 271768 157248 271788
rect 157248 271768 157300 271788
rect 157300 271768 157302 271788
rect 196622 271768 196678 271824
rect 158626 271652 158682 271688
rect 158626 271632 158628 271652
rect 158628 271632 158680 271652
rect 158680 271632 158682 271652
rect 161294 271632 161350 271688
rect 164146 271632 164202 271688
rect 117318 271496 117320 271516
rect 117320 271496 117372 271516
rect 117372 271496 117374 271516
rect 127622 271496 127678 271552
rect 196622 271496 196678 271552
rect 183466 271360 183522 271416
rect 183466 271124 183468 271144
rect 183468 271124 183520 271144
rect 183520 271124 183522 271144
rect 183466 271088 183522 271124
rect 106370 270952 106426 271008
rect 107658 270952 107714 271008
rect 111798 270952 111854 271008
rect 104898 270816 104954 270872
rect 106278 270816 106334 270872
rect 110418 270680 110474 270736
rect 107750 270544 107806 270600
rect 109038 270544 109094 270600
rect 113178 270544 113234 270600
rect 115846 270544 115902 270600
rect 117226 270544 117282 270600
rect 144918 270544 144974 270600
rect 147678 270544 147734 270600
rect 191746 253680 191802 253736
rect 179326 253172 179328 253192
rect 179328 253172 179380 253192
rect 179380 253172 179382 253192
rect 179326 253136 179382 253172
rect 180522 253136 180578 253192
rect 101034 166776 101090 166832
rect 103518 166776 103574 166832
rect 108302 166812 108304 166832
rect 108304 166812 108356 166832
rect 108356 166812 108358 166832
rect 108302 166776 108358 166812
rect 138478 166776 138534 166832
rect 140870 166796 140926 166832
rect 140870 166776 140872 166796
rect 140872 166776 140924 166796
rect 140924 166776 140926 166796
rect 145930 166776 145986 166832
rect 148506 166640 148562 166696
rect 163318 166640 163374 166696
rect 165894 166640 165950 166696
rect 107658 166504 107714 166560
rect 150898 166524 150954 166560
rect 150898 166504 150900 166524
rect 150900 166504 150952 166524
rect 150952 166504 150954 166524
rect 96066 166232 96122 166288
rect 98458 166252 98514 166288
rect 98458 166232 98460 166252
rect 98460 166232 98512 166252
rect 98512 166232 98514 166252
rect 81438 165552 81494 165608
rect 84290 165552 84346 165608
rect 91190 165552 91246 165608
rect 95238 165552 95294 165608
rect 99378 165552 99434 165608
rect 100850 165552 100906 165608
rect 105174 165552 105230 165608
rect 105726 165552 105782 165608
rect 106370 165552 106426 165608
rect 78678 164872 78734 164928
rect 76010 164328 76066 164384
rect 59358 140800 59414 140856
rect 75918 164192 75974 164248
rect 73802 145968 73858 146024
rect 77298 164192 77354 164248
rect 80058 164192 80114 164248
rect 82818 164192 82874 164248
rect 84198 164192 84254 164248
rect 90270 165008 90326 165064
rect 88338 164872 88394 164928
rect 85578 164192 85634 164248
rect 86958 164192 87014 164248
rect 88430 164192 88486 164248
rect 89902 164192 89958 164248
rect 91098 164192 91154 164248
rect 92478 164892 92534 164928
rect 92478 164872 92480 164892
rect 92480 164872 92532 164892
rect 92532 164872 92534 164892
rect 92570 164192 92626 164248
rect 93858 164192 93914 164248
rect 92570 145696 92626 145752
rect 96618 164192 96674 164248
rect 97998 164192 98054 164248
rect 100758 164192 100814 164248
rect 102138 164192 102194 164248
rect 103518 164192 103574 164248
rect 103518 146240 103574 146296
rect 102138 146104 102194 146160
rect 100758 145968 100814 146024
rect 153290 166504 153346 166560
rect 183282 166504 183338 166560
rect 108302 165552 108358 165608
rect 109682 165552 109738 165608
rect 110970 165552 111026 165608
rect 111890 165552 111946 165608
rect 113546 165552 113602 165608
rect 115938 165552 115994 165608
rect 117870 165552 117926 165608
rect 118330 165552 118386 165608
rect 119066 165552 119122 165608
rect 120906 165552 120962 165608
rect 123482 165552 123538 165608
rect 125874 165552 125930 165608
rect 128358 165552 128414 165608
rect 129738 165552 129794 165608
rect 132498 165572 132554 165608
rect 132498 165552 132500 165572
rect 132500 165552 132552 165572
rect 132552 165552 132554 165572
rect 111154 164600 111210 164656
rect 113178 165008 113234 165064
rect 114466 164872 114522 164928
rect 115938 164464 115994 164520
rect 117318 164464 117374 164520
rect 183374 165552 183430 165608
rect 197450 484916 197452 484936
rect 197452 484916 197504 484936
rect 197504 484916 197506 484936
rect 197450 484880 197506 484916
rect 198646 380976 198702 381032
rect 107658 145560 107714 145616
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 191286 144880 191342 144936
rect 77114 59744 77170 59800
rect 83094 59744 83150 59800
rect 94502 59744 94558 59800
rect 99470 59744 99526 59800
rect 102782 59744 102838 59800
rect 105910 59744 105966 59800
rect 89994 59472 90050 59528
rect 95882 59472 95938 59528
rect 96986 59472 97042 59528
rect 100758 59472 100814 59528
rect 101770 59472 101826 59528
rect 107566 59608 107622 59664
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 138386 58928 138442 58984
rect 84198 57976 84254 58032
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 78678 57840 78734 57896
rect 80426 57840 80482 57896
rect 81438 57840 81494 57896
rect 85394 57840 85450 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88338 57840 88394 57896
rect 88706 57840 88762 57896
rect 89718 57840 89774 57896
rect 91098 57840 91154 57896
rect 91466 57840 91522 57896
rect 93306 57840 93362 57896
rect 93674 57840 93730 57896
rect 98090 57840 98146 57896
rect 103794 57840 103850 57896
rect 108578 57840 108634 57896
rect 109498 57840 109554 57896
rect 112074 57840 112130 57896
rect 113178 57840 113234 57896
rect 114098 57840 114154 57896
rect 115938 57840 115994 57896
rect 117870 57840 117926 57896
rect 119066 57840 119122 57896
rect 123482 57840 123538 57896
rect 130842 57840 130898 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 77850 54712 77906 54768
rect 106278 57432 106334 57488
rect 110418 57432 110474 57488
rect 114558 57432 114614 57488
rect 116122 57432 116178 57488
rect 153290 57840 153346 57896
rect 183466 57860 183522 57896
rect 183466 57840 183468 57860
rect 183468 57840 183520 57860
rect 183520 57840 183522 57860
rect 198738 377984 198794 378040
rect 198922 460128 198978 460184
rect 200486 484744 200542 484800
rect 200302 484472 200358 484528
rect 199014 397432 199070 397488
rect 199290 395936 199346 395992
rect 199474 400288 199530 400344
rect 199842 400288 199898 400344
rect 199658 396752 199714 396808
rect 199382 394576 199438 394632
rect 199014 379344 199070 379400
rect 199750 394576 199806 394632
rect 199474 377440 199530 377496
rect 198830 353096 198886 353152
rect 198738 291624 198794 291680
rect 199198 292712 199254 292768
rect 199106 290944 199162 291000
rect 198922 288768 198978 288824
rect 198830 246200 198886 246256
rect 198738 184864 198794 184920
rect 198738 182008 198794 182064
rect 199014 288360 199070 288416
rect 199014 287544 199070 287600
rect 198922 182008 198978 182064
rect 199474 291624 199530 291680
rect 199934 395936 199990 395992
rect 199658 292712 199714 292768
rect 199566 290944 199622 291000
rect 199750 288360 199806 288416
rect 201498 484880 201554 484936
rect 201314 379480 201370 379536
rect 199382 186360 199438 186416
rect 199290 184864 199346 184920
rect 199106 183368 199162 183424
rect 199014 180648 199070 180704
rect 199014 179424 199070 179480
rect 198830 139168 198886 139224
rect 199198 179424 199254 179480
rect 199106 76336 199162 76392
rect 198738 74840 198794 74896
rect 199382 79328 199438 79384
rect 199290 77696 199346 77752
rect 199198 73616 199254 73672
rect 202326 468968 202382 469024
rect 202878 380704 202934 380760
rect 203614 485016 203670 485072
rect 202786 379480 202842 379536
rect 203706 471416 203762 471472
rect 203522 471280 203578 471336
rect 203614 465976 203670 466032
rect 203890 380296 203946 380352
rect 204810 378528 204866 378584
rect 204810 378120 204866 378176
rect 205638 485596 205640 485616
rect 205640 485596 205692 485616
rect 205692 485596 205694 485616
rect 205638 485560 205694 485596
rect 205638 485152 205694 485208
rect 205730 484472 205786 484528
rect 205546 413888 205602 413944
rect 205454 378120 205510 378176
rect 183190 57740 183192 57760
rect 183192 57740 183244 57760
rect 183244 57740 183246 57760
rect 183190 57704 183246 57740
rect 206190 379480 206246 379536
rect 206466 468832 206522 468888
rect 206650 270408 206706 270464
rect 207018 380588 207074 380624
rect 207018 380568 207020 380588
rect 207020 380568 207072 380588
rect 207072 380568 207074 380588
rect 207018 380160 207074 380216
rect 207938 380568 207994 380624
rect 208030 378936 208086 378992
rect 207938 377576 207994 377632
rect 207754 270952 207810 271008
rect 208398 485596 208400 485616
rect 208400 485596 208452 485616
rect 208452 485596 208454 485616
rect 208398 485560 208454 485596
rect 208398 380432 208454 380488
rect 208490 379072 208546 379128
rect 208490 378392 208546 378448
rect 208030 269728 208086 269784
rect 209134 468696 209190 468752
rect 209686 390632 209742 390688
rect 209502 379072 209558 379128
rect 209410 378392 209466 378448
rect 209318 269728 209374 269784
rect 211158 484880 211214 484936
rect 211250 484744 211306 484800
rect 210606 468560 210662 468616
rect 210974 379208 211030 379264
rect 210882 145696 210938 145752
rect 211066 378528 211122 378584
rect 157338 57568 157394 57624
rect 160098 57568 160154 57624
rect 165618 57568 165674 57624
rect 153290 56344 153346 56400
rect 119066 56072 119122 56128
rect 157338 54984 157394 55040
rect 211434 377848 211490 377904
rect 211434 377576 211490 377632
rect 211986 471552 212042 471608
rect 212630 380568 212686 380624
rect 212446 378528 212502 378584
rect 212446 378256 212502 378312
rect 212446 377848 212502 377904
rect 212354 376624 212410 376680
rect 212262 270000 212318 270056
rect 212906 380976 212962 381032
rect 212722 377576 212778 377632
rect 213274 377576 213330 377632
rect 213826 377848 213882 377904
rect 213274 145832 213330 145888
rect 165618 55120 165674 55176
rect 160098 54848 160154 54904
rect 214838 484472 214894 484528
rect 214378 270272 214434 270328
rect 214746 471144 214802 471200
rect 215482 380704 215538 380760
rect 215206 376624 215262 376680
rect 214930 270272 214986 270328
rect 214930 145560 214986 145616
rect 214930 55120 214986 55176
rect 215574 377848 215630 377904
rect 215666 377712 215722 377768
rect 215574 270000 215630 270056
rect 216034 271632 216090 271688
rect 216678 417832 216734 417888
rect 217046 414724 217102 414760
rect 217046 414704 217048 414724
rect 217048 414704 217100 414724
rect 217100 414704 217102 414724
rect 216862 413752 216918 413808
rect 216678 410896 216734 410952
rect 216678 390904 216734 390960
rect 216678 389272 216734 389328
rect 216678 389000 216734 389056
rect 216586 380704 216642 380760
rect 216494 376624 216550 376680
rect 216402 271360 216458 271416
rect 215850 145016 215906 145072
rect 216678 309032 216734 309088
rect 217322 409128 217378 409184
rect 217138 379480 217194 379536
rect 216954 309848 217010 309904
rect 216862 307672 216918 307728
rect 216678 284008 216734 284064
rect 216678 282376 216734 282432
rect 216770 282104 216826 282160
rect 216586 271360 216642 271416
rect 216862 270272 216918 270328
rect 216862 270000 216918 270056
rect 216862 203904 216918 203960
rect 216678 175344 216734 175400
rect 216402 146104 216458 146160
rect 216402 145016 216458 145072
rect 217690 411984 217746 412040
rect 217138 302096 217194 302152
rect 216954 202952 217010 203008
rect 216862 96872 216918 96928
rect 217506 374992 217562 375048
rect 217322 310936 217378 310992
rect 217506 310936 217562 310992
rect 217414 307672 217470 307728
rect 217414 306720 217470 306776
rect 217966 416880 218022 416936
rect 217874 409128 217930 409184
rect 217874 380840 217930 380896
rect 217874 379480 217930 379536
rect 217690 309032 217746 309088
rect 217690 307808 217746 307864
rect 217598 303864 217654 303920
rect 217506 203904 217562 203960
rect 217414 199824 217470 199880
rect 217230 196968 217286 197024
rect 217138 195200 217194 195256
rect 217046 176976 217102 177032
rect 217138 175072 217194 175128
rect 216954 95920 217010 95976
rect 216678 69944 216734 70000
rect 216678 68312 216734 68368
rect 217506 197376 217562 197432
rect 217414 92792 217470 92848
rect 217782 304952 217838 305008
rect 217690 200776 217746 200832
rect 217598 196968 217654 197024
rect 217598 195200 217654 195256
rect 217506 91024 217562 91080
rect 217230 89936 217286 89992
rect 218702 485288 218758 485344
rect 218058 379480 218114 379536
rect 218518 380296 218574 380352
rect 217966 309848 218022 309904
rect 217782 198056 217838 198112
rect 217782 197376 217838 197432
rect 217874 162716 217930 162752
rect 217874 162696 217876 162716
rect 217876 162696 217928 162716
rect 217928 162696 217930 162716
rect 218426 273264 218482 273320
rect 217690 93744 217746 93800
rect 217598 88168 217654 88224
rect 217966 68312 218022 68368
rect 218978 465704 219034 465760
rect 218702 60560 218758 60616
rect 219162 144880 219218 144936
rect 219254 60560 219310 60616
rect 219898 146240 219954 146296
rect 219898 144880 219954 144936
rect 223486 485016 223542 485072
rect 222566 482296 222622 482352
rect 226154 485152 226210 485208
rect 224866 484472 224922 484528
rect 223578 478216 223634 478272
rect 226522 475496 226578 475552
rect 229834 479576 229890 479632
rect 227994 476856 228050 476912
rect 231766 485288 231822 485344
rect 230754 476720 230810 476776
rect 232318 485424 232374 485480
rect 233606 485696 233662 485752
rect 234342 485152 234398 485208
rect 233974 480800 234030 480856
rect 235814 485560 235870 485616
rect 235906 484880 235962 484936
rect 234618 478352 234674 478408
rect 231950 475768 232006 475824
rect 236366 482432 236422 482488
rect 240322 475632 240378 475688
rect 247314 480936 247370 480992
rect 254122 475904 254178 475960
rect 256330 479712 256386 479768
rect 265070 468424 265126 468480
rect 277122 482568 277178 482624
rect 280710 481072 280766 481128
rect 297178 478488 297234 478544
rect 292578 465704 292634 465760
rect 316774 575592 316830 575648
rect 316774 570832 316830 570888
rect 315578 547984 315634 548040
rect 318246 640464 318302 640520
rect 317970 638152 318026 638208
rect 318062 633392 318118 633448
rect 317694 628632 317750 628688
rect 317418 623872 317474 623928
rect 317602 619112 317658 619168
rect 317970 614352 318026 614408
rect 317970 609592 318026 609648
rect 317970 604832 318026 604888
rect 317970 595312 318026 595368
rect 317970 590552 318026 590608
rect 317970 585792 318026 585848
rect 317970 580352 318026 580408
rect 317970 566072 318026 566128
rect 317970 561312 318026 561368
rect 318798 600072 318854 600128
rect 317418 556552 317474 556608
rect 318062 551792 318118 551848
rect 318062 549888 318118 549944
rect 317970 547032 318026 547088
rect 317970 542308 317972 542328
rect 317972 542308 318024 542328
rect 318024 542308 318026 542328
rect 317970 542272 318026 542308
rect 319718 640600 319774 640656
rect 328366 639240 328422 639296
rect 346398 639104 346454 639160
rect 392122 640600 392178 640656
rect 419170 640464 419226 640520
rect 405370 638968 405426 639024
rect 428370 566208 428426 566264
rect 318706 537512 318762 537568
rect 318614 532752 318670 532808
rect 427818 528536 427874 528592
rect 429290 591232 429346 591288
rect 391938 489096 391994 489152
rect 312542 482160 312598 482216
rect 298190 471144 298246 471200
rect 338486 466520 338542 466576
rect 339774 466540 339830 466576
rect 339774 466520 339776 466540
rect 339776 466520 339828 466540
rect 339828 466520 339830 466540
rect 350998 466520 351054 466576
rect 235998 380840 236054 380896
rect 237102 380840 237158 380896
rect 243082 380840 243138 380896
rect 245382 380840 245438 380896
rect 247590 380840 247646 380896
rect 254490 380840 254546 380896
rect 255870 380840 255926 380896
rect 256974 380840 257030 380896
rect 276018 380876 276020 380896
rect 276020 380876 276072 380896
rect 276072 380876 276074 380896
rect 276018 380840 276074 380876
rect 221002 378664 221058 378720
rect 221646 378800 221702 378856
rect 221278 378528 221334 378584
rect 221186 378256 221242 378312
rect 221646 378256 221702 378312
rect 222014 379072 222070 379128
rect 222014 378664 222070 378720
rect 233882 378664 233938 378720
rect 233882 378392 233938 378448
rect 221370 377712 221426 377768
rect 221830 377712 221886 377768
rect 244278 380296 244334 380352
rect 245658 379208 245714 379264
rect 259458 380568 259514 380624
rect 265254 380568 265310 380624
rect 270958 380568 271014 380624
rect 268658 379344 268714 379400
rect 248602 379208 248658 379264
rect 250074 379208 250130 379264
rect 251178 379208 251234 379264
rect 252282 379208 252338 379264
rect 253386 379208 253442 379264
rect 261666 379208 261722 379264
rect 248234 378392 248290 378448
rect 250626 378392 250682 378448
rect 253202 379072 253258 379128
rect 253202 378256 253258 378312
rect 253570 378392 253626 378448
rect 255962 378392 256018 378448
rect 258354 378392 258410 378448
rect 260930 378392 260986 378448
rect 263598 378392 263654 378448
rect 265346 378392 265402 378448
rect 268106 378392 268162 378448
rect 262770 378256 262826 378312
rect 266358 378256 266414 378312
rect 267554 378256 267610 378312
rect 271050 379344 271106 379400
rect 271970 379344 272026 379400
rect 273258 379380 273260 379400
rect 273260 379380 273312 379400
rect 273312 379380 273314 379400
rect 273258 379344 273314 379380
rect 274362 379364 274418 379400
rect 274362 379344 274364 379364
rect 274364 379344 274416 379364
rect 274416 379344 274418 379364
rect 275650 379380 275652 379400
rect 275652 379380 275704 379400
rect 275704 379380 275706 379400
rect 275650 379344 275706 379380
rect 285954 379344 286010 379400
rect 287610 379344 287666 379400
rect 290922 379344 290978 379400
rect 293314 379344 293370 379400
rect 295890 379344 295946 379400
rect 298098 379344 298154 379400
rect 300858 379344 300914 379400
rect 273442 379208 273498 379264
rect 277030 379208 277086 379264
rect 277858 379208 277914 379264
rect 279146 379208 279202 379264
rect 280802 379208 280858 379264
rect 283010 379208 283066 379264
rect 273258 377984 273314 378040
rect 276018 378120 276074 378176
rect 303066 379344 303122 379400
rect 305734 379344 305790 379400
rect 308402 379344 308458 379400
rect 310978 379380 310980 379400
rect 310980 379380 311032 379400
rect 311032 379380 311034 379400
rect 310978 379344 311034 379380
rect 313370 379364 313426 379400
rect 313370 379344 313372 379364
rect 313372 379344 313424 379364
rect 313424 379344 313426 379364
rect 315762 379380 315764 379400
rect 315764 379380 315816 379400
rect 315816 379380 315818 379400
rect 315762 379344 315818 379380
rect 318338 379344 318394 379400
rect 323306 379344 323362 379400
rect 325882 379208 325938 379264
rect 320914 378528 320970 378584
rect 343178 378392 343234 378448
rect 325882 375264 325938 375320
rect 343546 378256 343602 378312
rect 338486 358828 338542 358864
rect 338486 358808 338488 358828
rect 338488 358808 338540 358828
rect 338540 358808 338542 358828
rect 339866 358808 339922 358864
rect 351734 358808 351790 358864
rect 266358 273672 266414 273728
rect 278042 273672 278098 273728
rect 250718 273556 250774 273592
rect 250718 273536 250720 273556
rect 250720 273536 250772 273556
rect 250772 273536 250774 273556
rect 273350 273536 273406 273592
rect 275742 273536 275798 273592
rect 283470 273536 283526 273592
rect 285954 273264 286010 273320
rect 287978 272856 288034 272912
rect 288162 272856 288218 272912
rect 290922 272876 290978 272912
rect 290922 272856 290924 272876
rect 290924 272856 290976 272876
rect 290976 272856 290978 272876
rect 293314 272856 293370 272912
rect 300858 272856 300914 272912
rect 298466 272720 298522 272776
rect 287978 272584 288034 272640
rect 305826 272604 305882 272640
rect 305826 272584 305828 272604
rect 305828 272584 305880 272604
rect 305880 272584 305882 272604
rect 320914 272584 320970 272640
rect 235998 272176 236054 272232
rect 265162 272176 265218 272232
rect 258262 271496 258318 271552
rect 263598 271496 263654 271552
rect 264978 271516 265034 271552
rect 264978 271496 264980 271516
rect 264980 271496 265032 271516
rect 265032 271496 265034 271516
rect 252558 271224 252614 271280
rect 247038 271088 247094 271144
rect 255318 271088 255374 271144
rect 260838 271244 260894 271280
rect 260838 271224 260840 271244
rect 260840 271224 260892 271244
rect 260892 271224 260894 271244
rect 253938 270816 253994 270872
rect 244370 270680 244426 270736
rect 251270 270680 251326 270736
rect 239126 270544 239182 270600
rect 242898 270544 242954 270600
rect 244278 270544 244334 270600
rect 229190 268368 229246 268424
rect 245658 270544 245714 270600
rect 247038 270544 247094 270600
rect 248510 270544 248566 270600
rect 249798 270544 249854 270600
rect 251178 270544 251234 270600
rect 252558 270544 252614 270600
rect 255318 270680 255374 270736
rect 259550 270680 259606 270736
rect 256698 270544 256754 270600
rect 258078 270544 258134 270600
rect 259458 270544 259514 270600
rect 260838 270544 260894 270600
rect 262218 270544 262274 270600
rect 263598 270544 263654 270600
rect 268198 271768 268254 271824
rect 270498 271768 270554 271824
rect 276018 271768 276074 271824
rect 280158 271768 280214 271824
rect 307758 271788 307814 271824
rect 307758 271768 307760 271788
rect 307760 271768 307812 271788
rect 307812 271768 307814 271788
rect 268014 271496 268070 271552
rect 313278 271804 313280 271824
rect 313280 271804 313332 271824
rect 313332 271804 313334 271824
rect 313278 271768 313334 271804
rect 343546 271804 343548 271824
rect 343548 271804 343600 271824
rect 343600 271804 343602 271824
rect 343546 271768 343602 271804
rect 271878 271496 271934 271552
rect 277122 271496 277178 271552
rect 343546 271496 343602 271552
rect 266358 270544 266414 270600
rect 269118 270544 269174 270600
rect 270498 270544 270554 270600
rect 277674 271380 277730 271416
rect 277674 271360 277676 271380
rect 277676 271360 277728 271380
rect 277728 271360 277730 271380
rect 280066 270816 280122 270872
rect 273166 270544 273222 270600
rect 340786 253408 340842 253464
rect 351826 253172 351828 253192
rect 351828 253172 351880 253192
rect 351880 253172 351882 253192
rect 351826 253136 351882 253172
rect 339406 253000 339462 253056
rect 231858 251776 231914 251832
rect 285954 166660 286010 166696
rect 285954 166640 285956 166660
rect 285956 166640 286008 166660
rect 286008 166640 286010 166660
rect 291014 166640 291070 166696
rect 293406 166640 293462 166696
rect 295890 166640 295946 166696
rect 298466 166640 298522 166696
rect 305918 166640 305974 166696
rect 260930 166504 260986 166560
rect 265898 166504 265954 166560
rect 270866 166504 270922 166560
rect 235998 165552 236054 165608
rect 238758 165552 238814 165608
rect 242898 165552 242954 165608
rect 247038 165552 247094 165608
rect 247682 165552 247738 165608
rect 249798 165552 249854 165608
rect 252558 165552 252614 165608
rect 258078 165552 258134 165608
rect 260838 165552 260894 165608
rect 264978 165552 265034 165608
rect 267646 165552 267702 165608
rect 236090 164192 236146 164248
rect 237378 164192 237434 164248
rect 220082 145696 220138 145752
rect 240138 164192 240194 164248
rect 241518 164192 241574 164248
rect 237378 145832 237434 145888
rect 244278 164464 244334 164520
rect 244370 164192 244426 164248
rect 245658 164192 245714 164248
rect 251270 164464 251326 164520
rect 259550 164464 259606 164520
rect 248418 164192 248474 164248
rect 249798 164192 249854 164248
rect 251178 164192 251234 164248
rect 252558 164192 252614 164248
rect 253938 164192 253994 164248
rect 255318 164192 255374 164248
rect 256698 164192 256754 164248
rect 258078 164192 258134 164248
rect 259458 164192 259514 164248
rect 263506 164192 263562 164248
rect 263782 164192 263838 164248
rect 266358 164464 266414 164520
rect 267738 164192 267794 164248
rect 263598 146104 263654 146160
rect 267922 165552 267978 165608
rect 280158 165552 280214 165608
rect 283378 165552 283434 165608
rect 300858 165552 300914 165608
rect 308402 165552 308458 165608
rect 323030 165552 323086 165608
rect 325882 165572 325938 165608
rect 325882 165552 325884 165572
rect 325884 165552 325936 165572
rect 325936 165552 325938 165572
rect 271878 165144 271934 165200
rect 275926 165144 275982 165200
rect 269118 164192 269174 164248
rect 270498 164192 270554 164248
rect 267830 146240 267886 146296
rect 267738 145696 267794 145752
rect 274454 164464 274510 164520
rect 274546 164192 274602 164248
rect 276018 164192 276074 164248
rect 277398 165164 277454 165200
rect 277398 165144 277400 165164
rect 277400 165144 277452 165164
rect 277452 165144 277454 165164
rect 280066 165144 280122 165200
rect 278686 164192 278742 164248
rect 276018 146376 276074 146432
rect 269118 145560 269174 145616
rect 343270 165572 343326 165608
rect 343270 165552 343272 165572
rect 343272 165552 343324 165572
rect 343324 165552 343326 165572
rect 343454 165552 343510 165608
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 237102 59744 237158 59800
rect 255870 59744 255926 59800
rect 256974 59744 257030 59800
rect 262862 59744 262918 59800
rect 263874 59744 263930 59800
rect 258078 59608 258134 59664
rect 260654 59608 260710 59664
rect 261758 59608 261814 59664
rect 308494 59608 308550 59664
rect 315854 59608 315910 59664
rect 279238 59200 279294 59256
rect 290922 59200 290978 59256
rect 300858 59200 300914 59256
rect 320914 59200 320970 59256
rect 325882 59200 325938 59256
rect 235998 57840 236054 57896
rect 237378 57840 237434 57896
rect 239126 57840 239182 57896
rect 240138 57840 240194 57896
rect 241610 57840 241666 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 245290 57840 245346 57896
rect 245658 57840 245714 57896
rect 247038 57840 247094 57896
rect 248602 57840 248658 57896
rect 249798 57840 249854 57896
rect 251178 57840 251234 57896
rect 251362 57840 251418 57896
rect 253386 57840 253442 57896
rect 253938 57840 253994 57896
rect 258354 57840 258410 57896
rect 264978 57840 265034 57896
rect 266358 57840 266414 57896
rect 268474 57840 268530 57896
rect 271050 57840 271106 57896
rect 271878 57840 271934 57896
rect 273258 57840 273314 57896
rect 275098 57840 275154 57896
rect 283470 57840 283526 57896
rect 293314 57840 293370 57896
rect 295890 57840 295946 57896
rect 298098 57840 298154 57896
rect 303434 57840 303490 57896
rect 305826 57840 305882 57896
rect 310978 57860 311034 57896
rect 310978 57840 310980 57860
rect 310980 57840 311032 57860
rect 311032 57840 311034 57860
rect 266450 57568 266506 57624
rect 269118 57568 269174 57624
rect 269118 55120 269174 55176
rect 273350 57568 273406 57624
rect 277398 57568 277454 57624
rect 313370 57840 313426 57896
rect 318338 57840 318394 57896
rect 323306 57876 323308 57896
rect 323308 57876 323360 57896
rect 323360 57876 323362 57896
rect 323306 57840 323362 57876
rect 343178 57860 343234 57896
rect 343178 57840 343180 57860
rect 343180 57840 343232 57860
rect 343232 57840 343234 57860
rect 343454 57876 343456 57896
rect 343456 57876 343508 57896
rect 343508 57876 343510 57896
rect 343454 57840 343510 57876
rect 358634 417424 358690 417480
rect 358818 460128 358874 460184
rect 359094 398112 359150 398168
rect 359002 396752 359058 396808
rect 358910 394032 358966 394088
rect 359186 395256 359242 395312
rect 359830 400288 359886 400344
rect 358910 353096 358966 353152
rect 358818 289720 358874 289776
rect 358818 288768 358874 288824
rect 359094 292712 359150 292768
rect 359094 291760 359150 291816
rect 359002 290944 359058 291000
rect 359002 288360 359058 288416
rect 359002 287544 359058 287600
rect 358910 246200 358966 246256
rect 358818 182008 358874 182064
rect 359278 292712 359334 292768
rect 359186 288360 359242 288416
rect 359554 291760 359610 291816
rect 359554 290944 359610 291000
rect 359462 289720 359518 289776
rect 359370 186360 359426 186416
rect 359094 184864 359150 184920
rect 359002 180648 359058 180704
rect 358910 139304 358966 139360
rect 359278 183504 359334 183560
rect 359186 182008 359242 182064
rect 359094 78240 359150 78296
rect 359554 183504 359610 183560
rect 359370 79872 359426 79928
rect 359278 76880 359334 76936
rect 359186 75384 359242 75440
rect 359002 74024 359058 74080
rect 361118 272992 361174 273048
rect 366546 164600 366602 164656
rect 369674 379072 369730 379128
rect 369766 378936 369822 378992
rect 370410 380840 370466 380896
rect 370318 145696 370374 145752
rect 369030 145560 369086 145616
rect 371790 374584 371846 374640
rect 371606 272856 371662 272912
rect 372526 378392 372582 378448
rect 372250 270816 372306 270872
rect 373170 270000 373226 270056
rect 372986 269728 373042 269784
rect 373630 378800 373686 378856
rect 373906 379208 373962 379264
rect 373906 378800 373962 378856
rect 374366 270408 374422 270464
rect 373538 163376 373594 163432
rect 374550 270952 374606 271008
rect 375010 274624 375066 274680
rect 374918 270952 374974 271008
rect 376022 165280 376078 165336
rect 377218 416880 377274 416936
rect 377126 411984 377182 412040
rect 377218 410896 377274 410952
rect 376942 390904 376998 390960
rect 376942 389272 376998 389328
rect 376942 389000 376998 389056
rect 376942 380976 376998 381032
rect 376574 379480 376630 379536
rect 376390 271632 376446 271688
rect 376206 271496 376262 271552
rect 377586 417832 377642 417888
rect 377494 413888 377550 413944
rect 377494 411984 377550 412040
rect 377402 409148 377458 409184
rect 377402 409128 377404 409148
rect 377404 409128 377456 409148
rect 377456 409128 377458 409148
rect 376942 378120 376998 378176
rect 376942 310800 376998 310856
rect 376758 282104 376814 282160
rect 376942 284008 376998 284064
rect 376942 282240 376998 282296
rect 376666 269048 376722 269104
rect 376758 204176 376814 204232
rect 377218 309984 377274 310040
rect 376942 203904 376998 203960
rect 376758 202952 376814 203008
rect 376850 201320 376906 201376
rect 376758 95920 376814 95976
rect 376942 198736 376998 198792
rect 377862 416880 377918 416936
rect 377678 414724 377734 414760
rect 377678 414704 377680 414724
rect 377680 414704 377732 414724
rect 377732 414704 377734 414724
rect 377586 310800 377642 310856
rect 377770 410896 377826 410952
rect 377678 307808 377734 307864
rect 377586 304952 377642 305008
rect 377402 302096 377458 302152
rect 377218 204176 377274 204232
rect 377310 196968 377366 197024
rect 377034 176976 377090 177032
rect 376942 175344 376998 175400
rect 376850 93744 376906 93800
rect 377218 145696 377274 145752
rect 377034 96872 377090 96928
rect 376942 92792 376998 92848
rect 376942 69944 376998 70000
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 377402 195200 377458 195256
rect 377402 175072 377458 175128
rect 377402 163376 377458 163432
rect 377402 162968 377458 163024
rect 377954 413888 378010 413944
rect 377862 309984 377918 310040
rect 378046 409128 378102 409184
rect 377954 306720 378010 306776
rect 377862 303864 377918 303920
rect 377678 201320 377734 201376
rect 377678 200776 377734 200832
rect 377586 198056 377642 198112
rect 378046 302096 378102 302152
rect 377954 199824 378010 199880
rect 377954 198736 378010 198792
rect 377862 196968 377918 197024
rect 377954 195200 378010 195256
rect 377770 91024 377826 91080
rect 377310 89936 377366 89992
rect 378690 270272 378746 270328
rect 378782 165416 378838 165472
rect 430578 634072 430634 634128
rect 580170 683848 580226 683904
rect 430854 640328 430910 640384
rect 430762 629312 430818 629368
rect 430670 624552 430726 624608
rect 456798 627680 456854 627736
rect 430854 619792 430910 619848
rect 430578 610272 430634 610328
rect 429474 595992 429530 596048
rect 429382 538192 429438 538248
rect 429566 586608 429622 586664
rect 429658 557232 429714 557288
rect 430670 605512 430726 605568
rect 477130 627816 477186 627872
rect 488722 627816 488778 627872
rect 506754 627816 506810 627872
rect 457534 621560 457590 621616
rect 510618 618840 510674 618896
rect 457626 615440 457682 615496
rect 457534 596400 457590 596456
rect 457442 590280 457498 590336
rect 457442 584160 457498 584216
rect 430762 581032 430818 581088
rect 430854 576272 430910 576328
rect 430946 571512 431002 571568
rect 431038 561992 431094 562048
rect 431130 552472 431186 552528
rect 431222 547712 431278 547768
rect 431314 542952 431370 543008
rect 431406 533432 431462 533488
rect 580262 630808 580318 630864
rect 512090 624960 512146 625016
rect 511998 612040 512054 612096
rect 457718 609320 457774 609376
rect 511998 605920 512054 605976
rect 457810 602520 457866 602576
rect 457534 478080 457590 478136
rect 506478 487736 506534 487792
rect 512182 599800 512238 599856
rect 512090 593680 512146 593736
rect 511998 485152 512054 485208
rect 512274 587560 512330 587616
rect 513010 580760 513066 580816
rect 580262 577632 580318 577688
rect 512090 479440 512146 479496
rect 483018 475360 483074 475416
rect 498198 466556 498200 466576
rect 498200 466556 498252 466576
rect 498252 466556 498254 466576
rect 498198 466520 498254 466556
rect 499762 466540 499818 466576
rect 499762 466520 499764 466540
rect 499764 466520 499816 466540
rect 499816 466520 499818 466540
rect 510894 466540 510950 466576
rect 510894 466520 510896 466540
rect 510896 466520 510948 466540
rect 510948 466520 510950 466540
rect 421102 380704 421158 380760
rect 421746 380704 421802 380760
rect 425978 380704 426034 380760
rect 433614 380704 433670 380760
rect 434350 380724 434406 380760
rect 434350 380704 434352 380724
rect 434352 380704 434404 380724
rect 434404 380704 434406 380724
rect 408682 380568 408738 380624
rect 413466 380568 413522 380624
rect 422850 380568 422906 380624
rect 425242 380568 425298 380624
rect 436006 380704 436062 380760
rect 438490 380704 438546 380760
rect 440882 380704 440938 380760
rect 443458 380704 443514 380760
rect 379058 146240 379114 146296
rect 378690 146104 378746 146160
rect 377954 88168 378010 88224
rect 379058 145832 379114 145888
rect 380990 379344 381046 379400
rect 380990 378800 381046 378856
rect 436926 380568 436982 380624
rect 465906 380568 465962 380624
rect 396170 379344 396226 379400
rect 405738 379344 405794 379400
rect 407578 379344 407634 379400
rect 408314 379364 408370 379400
rect 408314 379344 408316 379364
rect 408316 379344 408368 379364
rect 408368 379344 408370 379364
rect 381174 378800 381230 378856
rect 381082 378528 381138 378584
rect 402978 379208 403034 379264
rect 405370 379208 405426 379264
rect 396078 378548 396134 378584
rect 396078 378528 396080 378548
rect 396080 378528 396132 378548
rect 396132 378528 396134 378548
rect 403622 378528 403678 378584
rect 410614 379344 410670 379400
rect 411258 379344 411314 379400
rect 412362 379344 412418 379400
rect 413098 379344 413154 379400
rect 423402 379344 423458 379400
rect 427450 379380 427452 379400
rect 427452 379380 427504 379400
rect 427504 379380 427506 379400
rect 427450 379344 427506 379380
rect 439042 379344 439098 379400
rect 445850 379344 445906 379400
rect 448150 379344 448206 379400
rect 451002 379344 451058 379400
rect 452750 379344 452806 379400
rect 455510 379344 455566 379400
rect 458362 379344 458418 379400
rect 409970 379208 410026 379264
rect 414570 379208 414626 379264
rect 415398 379208 415454 379264
rect 416042 379208 416098 379264
rect 418342 379208 418398 379264
rect 418250 378800 418306 378856
rect 416962 378120 417018 378176
rect 418158 378120 418214 378176
rect 419814 378120 419870 378176
rect 437754 379208 437810 379264
rect 428186 378528 428242 378584
rect 430670 378528 430726 378584
rect 423954 378120 424010 378176
rect 426438 378120 426494 378176
rect 428278 378256 428334 378312
rect 429382 378120 429438 378176
rect 431130 378120 431186 378176
rect 432234 378120 432290 378176
rect 463514 379208 463570 379264
rect 473450 379208 473506 379264
rect 474738 379208 474794 379264
rect 480810 379208 480866 379264
rect 503074 379208 503130 379264
rect 503534 379208 503590 379264
rect 467930 378800 467986 378856
rect 470874 378800 470930 378856
rect 477590 378800 477646 378856
rect 483386 378800 483442 378856
rect 480810 376624 480866 376680
rect 419814 374584 419870 374640
rect 498934 358808 498990 358864
rect 500774 358808 500830 358864
rect 510894 358828 510950 358864
rect 510894 358808 510896 358828
rect 510896 358808 510948 358828
rect 510948 358808 510950 358828
rect 421102 273536 421158 273592
rect 451002 273536 451058 273592
rect 423402 273264 423458 273320
rect 423770 273264 423826 273320
rect 426438 273264 426494 273320
rect 425978 272720 426034 272776
rect 428186 272720 428242 272776
rect 431130 272720 431186 272776
rect 468482 272756 468484 272776
rect 468484 272756 468536 272776
rect 468536 272756 468538 272776
rect 468482 272720 468538 272756
rect 470874 272720 470930 272776
rect 473450 272740 473506 272776
rect 473450 272720 473452 272740
rect 473452 272720 473504 272740
rect 473504 272720 473506 272740
rect 475842 272604 475898 272640
rect 475842 272584 475844 272604
rect 475844 272584 475896 272604
rect 475896 272584 475898 272604
rect 478418 272584 478474 272640
rect 401690 272176 401746 272232
rect 416042 272176 416098 272232
rect 437938 272176 437994 272232
rect 455786 272176 455842 272232
rect 396722 271224 396778 271280
rect 396078 270544 396134 270600
rect 389270 269728 389326 269784
rect 379702 145560 379758 145616
rect 397458 270544 397514 270600
rect 398838 270544 398894 270600
rect 400218 270544 400274 270600
rect 402978 271768 403034 271824
rect 412822 271768 412878 271824
rect 412822 271360 412878 271416
rect 413098 271224 413154 271280
rect 409878 271088 409934 271144
rect 414018 271088 414074 271144
rect 404358 270952 404414 271008
rect 407118 270972 407174 271008
rect 407118 270952 407120 270972
rect 407120 270952 407172 270972
rect 407172 270952 407174 270972
rect 403530 270544 403586 270600
rect 411258 270952 411314 271008
rect 405738 270544 405794 270600
rect 407118 270544 407174 270600
rect 408498 270544 408554 270600
rect 409878 270544 409934 270600
rect 412914 270680 412970 270736
rect 411350 270544 411406 270600
rect 416778 271088 416834 271144
rect 418250 270680 418306 270736
rect 418158 270544 418214 270600
rect 419538 270544 419594 270600
rect 420918 270544 420974 270600
rect 433338 271768 433394 271824
rect 434718 271768 434774 271824
rect 437478 271768 437534 271824
rect 445758 271768 445814 271824
rect 447138 271768 447194 271824
rect 452658 271768 452714 271824
rect 458178 271788 458234 271824
rect 458178 271768 458180 271788
rect 458180 271768 458232 271788
rect 458232 271768 458234 271788
rect 503626 271632 503682 271688
rect 440238 271380 440294 271416
rect 440238 271360 440240 271380
rect 440240 271360 440292 271380
rect 440292 271360 440294 271380
rect 440146 271224 440202 271280
rect 442998 271244 443054 271280
rect 442998 271224 443000 271244
rect 443000 271224 443052 271244
rect 443052 271224 443054 271244
rect 503626 271244 503682 271280
rect 503626 271224 503628 271244
rect 503628 271224 503680 271244
rect 503680 271224 503682 271244
rect 433338 271088 433394 271144
rect 427082 270952 427138 271008
rect 429198 270952 429254 271008
rect 425702 270680 425758 270736
rect 434718 270952 434774 271008
rect 436098 270952 436154 271008
rect 436190 270544 436246 270600
rect 500866 253308 500868 253328
rect 500868 253308 500920 253328
rect 500920 253308 500922 253328
rect 500866 253272 500922 253308
rect 499210 252728 499266 252784
rect 510894 252612 510950 252648
rect 510894 252592 510896 252612
rect 510896 252592 510948 252612
rect 510948 252592 510950 252612
rect 396722 251776 396778 251832
rect 418434 166776 418490 166832
rect 421010 166812 421012 166832
rect 421012 166812 421064 166832
rect 421064 166812 421066 166832
rect 421010 166776 421066 166812
rect 423402 166776 423458 166832
rect 445850 166796 445906 166832
rect 445850 166776 445852 166796
rect 445852 166776 445904 166796
rect 445904 166776 445906 166796
rect 470966 166776 471022 166832
rect 473450 166776 473506 166832
rect 475842 166776 475898 166832
rect 478418 166776 478474 166832
rect 480902 166776 480958 166832
rect 483386 166640 483442 166696
rect 485962 166640 486018 166696
rect 503258 166504 503314 166560
rect 428186 166232 428242 166288
rect 430946 166252 431002 166288
rect 430946 166232 430948 166252
rect 430948 166232 431000 166252
rect 431000 166232 431002 166252
rect 397458 165552 397514 165608
rect 401598 165552 401654 165608
rect 404358 165552 404414 165608
rect 407118 165552 407174 165608
rect 409878 165552 409934 165608
rect 415398 165552 415454 165608
rect 416042 165552 416098 165608
rect 418618 165552 418674 165608
rect 423678 165552 423734 165608
rect 427634 165552 427690 165608
rect 433338 165588 433340 165608
rect 433340 165588 433392 165608
rect 433392 165588 433394 165608
rect 433338 165552 433394 165588
rect 433522 165552 433578 165608
rect 434718 165552 434774 165608
rect 437754 165552 437810 165608
rect 438030 165552 438086 165608
rect 442998 165552 443054 165608
rect 447322 165552 447378 165608
rect 449898 165552 449954 165608
rect 452658 165552 452714 165608
rect 455418 165552 455474 165608
rect 458362 165572 458418 165608
rect 458362 165552 458364 165572
rect 458364 165552 458416 165572
rect 458416 165552 458418 165572
rect 396078 164328 396134 164384
rect 396170 164192 396226 164248
rect 398838 164192 398894 164248
rect 400218 164192 400274 164248
rect 402978 164328 403034 164384
rect 403070 164192 403126 164248
rect 412638 164756 412694 164792
rect 412638 164736 412640 164756
rect 412640 164736 412692 164756
rect 412692 164736 412694 164756
rect 411350 164328 411406 164384
rect 405738 164192 405794 164248
rect 407210 164192 407266 164248
rect 408498 164192 408554 164248
rect 409970 164192 410026 164248
rect 411258 164192 411314 164248
rect 412730 164192 412786 164248
rect 414018 164192 414074 164248
rect 416778 164192 416834 164248
rect 418158 164192 418214 164248
rect 420918 164736 420974 164792
rect 419538 164192 419594 164248
rect 422298 164192 422354 164248
rect 415398 145832 415454 145888
rect 426346 164192 426402 164248
rect 433338 165028 433394 165064
rect 433338 165008 433340 165028
rect 433340 165008 433392 165028
rect 433392 165008 433394 165028
rect 427726 164192 427782 164248
rect 426438 146240 426494 146296
rect 423678 145696 423734 145752
rect 436098 164464 436154 164520
rect 429290 164328 429346 164384
rect 429106 164192 429162 164248
rect 430578 164192 430634 164248
rect 431958 164192 432014 164248
rect 434718 164192 434774 164248
rect 503350 165552 503406 165608
rect 440146 164192 440202 164248
rect 518898 459584 518954 459640
rect 519542 459584 519598 459640
rect 518990 400288 519046 400344
rect 519082 398112 519138 398168
rect 440330 164872 440386 164928
rect 427818 145560 427874 145616
rect 510618 145424 510674 145480
rect 498658 144880 498714 144936
rect 500222 144880 500278 144936
rect 440238 144064 440294 144120
rect 396078 59764 396134 59800
rect 396078 59744 396080 59764
rect 396080 59744 396132 59764
rect 396132 59744 396134 59764
rect 397090 59744 397146 59800
rect 416042 59744 416098 59800
rect 416962 59744 417018 59800
rect 422850 59744 422906 59800
rect 423954 59744 424010 59800
rect 403070 59608 403126 59664
rect 404174 59608 404230 59664
rect 412546 59608 412602 59664
rect 398194 57840 398250 57896
rect 398838 57840 398894 57896
rect 400402 57840 400458 57896
rect 401598 57840 401654 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407210 57840 407266 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 411258 56888 411314 56944
rect 423494 59608 423550 59664
rect 418158 59336 418214 59392
rect 419354 59336 419410 59392
rect 420642 59336 420698 59392
rect 421746 59336 421802 59392
rect 425978 59336 426034 59392
rect 428186 59336 428242 59392
rect 453394 59336 453450 59392
rect 475842 58928 475898 58984
rect 519266 396752 519322 396808
rect 519174 395256 519230 395312
rect 519358 394032 519414 394088
rect 518990 293800 519046 293856
rect 518898 292440 518954 292496
rect 519082 290264 519138 290320
rect 518990 287544 519046 287600
rect 518898 186360 518954 186416
rect 414570 57840 414626 57896
rect 415490 57840 415546 57896
rect 418434 57840 418490 57896
rect 425058 57840 425114 57896
rect 426438 57840 426494 57896
rect 427634 57840 427690 57896
rect 427818 57840 427874 57896
rect 429198 57840 429254 57896
rect 431130 57840 431186 57896
rect 431958 57840 432014 57896
rect 433338 57840 433394 57896
rect 433522 57840 433578 57896
rect 435730 57840 435786 57896
rect 435914 57840 435970 57896
rect 438490 57840 438546 57896
rect 443458 57840 443514 57896
rect 445850 57840 445906 57896
rect 448242 57840 448298 57896
rect 465906 57840 465962 57896
rect 478418 57876 478420 57896
rect 478420 57876 478472 57896
rect 478472 57876 478474 57896
rect 478418 57840 478474 57876
rect 485962 57860 486018 57896
rect 485962 57840 485964 57860
rect 485964 57840 486016 57860
rect 486016 57840 486018 57860
rect 412546 56888 412602 56944
rect 412638 56752 412694 56808
rect 425058 54984 425114 55040
rect 433246 57568 433302 57624
rect 433246 57160 433302 57216
rect 433430 57568 433486 57624
rect 436098 57568 436154 57624
rect 438858 57568 438914 57624
rect 503258 57876 503260 57896
rect 503260 57876 503312 57896
rect 503312 57876 503314 57896
rect 503258 57840 503314 57876
rect 503534 57860 503590 57896
rect 519266 352824 519322 352880
rect 519174 288768 519230 288824
rect 519082 183368 519138 183424
rect 518990 180648 519046 180704
rect 518898 79872 518954 79928
rect 519358 293800 519414 293856
rect 519266 246200 519322 246256
rect 519174 181872 519230 181928
rect 580170 511264 580226 511320
rect 580262 458088 580318 458144
rect 578882 404912 578938 404968
rect 580170 378392 580226 378448
rect 519542 352824 519598 352880
rect 519542 292440 519598 292496
rect 519358 186360 519414 186416
rect 580354 351872 580410 351928
rect 580262 325216 580318 325272
rect 519634 290264 519690 290320
rect 520186 288768 520242 288824
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 519542 184728 519598 184784
rect 520186 184728 520242 184784
rect 519358 181872 519414 181928
rect 519266 139304 519322 139360
rect 519082 76744 519138 76800
rect 520094 183368 520150 183424
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519450 78240 519506 78296
rect 519358 75384 519414 75440
rect 518990 74160 519046 74216
rect 503534 57840 503536 57860
rect 503536 57840 503588 57860
rect 503588 57840 503590 57860
rect 438858 55120 438914 55176
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
rect 140042 3984 140098 4040
rect 129370 3848 129426 3904
rect 132958 3304 133014 3360
rect 136454 3168 136510 3224
rect 147126 3712 147182 3768
rect 143538 3576 143594 3632
rect 150622 3440 150678 3496
rect 367098 2896 367154 2952
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 319713 640658 319779 640661
rect 392117 640658 392183 640661
rect 319713 640656 392183 640658
rect 319713 640600 319718 640656
rect 319774 640600 392122 640656
rect 392178 640600 392183 640656
rect 319713 640598 392183 640600
rect 319713 640595 319779 640598
rect 392117 640595 392183 640598
rect 318241 640522 318307 640525
rect 419165 640522 419231 640525
rect 318241 640520 419231 640522
rect 318241 640464 318246 640520
rect 318302 640464 419170 640520
rect 419226 640464 419231 640520
rect 318241 640462 419231 640464
rect 318241 640459 318307 640462
rect 419165 640459 419231 640462
rect 280981 640386 281047 640389
rect 430849 640386 430915 640389
rect 280981 640384 430915 640386
rect 280981 640328 280986 640384
rect 281042 640328 430854 640384
rect 430910 640328 430915 640384
rect 280981 640326 430915 640328
rect 280981 640323 281047 640326
rect 430849 640323 430915 640326
rect 53046 639236 53052 639300
rect 53116 639298 53122 639300
rect 328361 639298 328427 639301
rect 53116 639296 328427 639298
rect 53116 639240 328366 639296
rect 328422 639240 328427 639296
rect 53116 639238 328427 639240
rect 53116 639236 53122 639238
rect 328361 639235 328427 639238
rect 51574 639100 51580 639164
rect 51644 639162 51650 639164
rect 346393 639162 346459 639165
rect 51644 639160 346459 639162
rect 51644 639104 346398 639160
rect 346454 639104 346459 639160
rect 51644 639102 346459 639104
rect 51644 639100 51650 639102
rect 346393 639099 346459 639102
rect 54334 638964 54340 639028
rect 54404 639026 54410 639028
rect 405365 639026 405431 639029
rect 54404 639024 405431 639026
rect 54404 638968 405370 639024
rect 405426 638968 405431 639024
rect 54404 638966 405431 638968
rect 54404 638964 54410 638966
rect 405365 638963 405431 638966
rect 317965 638210 318031 638213
rect 317965 638208 320068 638210
rect 317965 638152 317970 638208
rect 318026 638152 320068 638208
rect 317965 638150 320068 638152
rect 317965 638147 318031 638150
rect 430573 634130 430639 634133
rect 428812 634128 430639 634130
rect 428812 634072 430578 634128
rect 430634 634072 430639 634128
rect 428812 634070 430639 634072
rect 430573 634067 430639 634070
rect 318057 633450 318123 633453
rect 318057 633448 320068 633450
rect 318057 633392 318062 633448
rect 318118 633392 320068 633448
rect 318057 633390 320068 633392
rect 318057 633387 318123 633390
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect 430757 629370 430823 629373
rect 428812 629368 430823 629370
rect 428812 629312 430762 629368
rect 430818 629312 430823 629368
rect 428812 629310 430823 629312
rect 430757 629307 430823 629310
rect 58985 628690 59051 628693
rect 137277 628690 137343 628693
rect 215937 628690 216003 628693
rect 317689 628690 317755 628693
rect 58985 628688 60106 628690
rect 58985 628632 58990 628688
rect 59046 628632 60106 628688
rect 58985 628630 60106 628632
rect 58985 628627 59051 628630
rect 60046 628592 60106 628630
rect 137277 628688 140146 628690
rect 137277 628632 137282 628688
rect 137338 628632 140146 628688
rect 137277 628630 140146 628632
rect 137277 628627 137343 628630
rect 140086 628592 140146 628630
rect 215937 628688 220186 628690
rect 215937 628632 215942 628688
rect 215998 628632 220186 628688
rect 215937 628630 220186 628632
rect 215937 628627 216003 628630
rect 220126 628592 220186 628630
rect 317689 628688 320068 628690
rect 317689 628632 317694 628688
rect 317750 628632 320068 628688
rect 317689 628630 320068 628632
rect 317689 628627 317755 628630
rect 122925 628010 122991 628013
rect 201769 628010 201835 628013
rect 281533 628010 281599 628013
rect 120766 628008 122991 628010
rect 120766 627952 122930 628008
rect 122986 627952 122991 628008
rect 120766 627950 122991 627952
rect 120766 627912 120826 627950
rect 122925 627947 122991 627950
rect 200806 628008 201835 628010
rect 200806 627952 201774 628008
rect 201830 627952 201835 628008
rect 200806 627950 201835 627952
rect 200806 627912 200866 627950
rect 201769 627947 201835 627950
rect 280846 628008 281599 628010
rect 280846 627952 281538 628008
rect 281594 627952 281599 628008
rect 280846 627950 281599 627952
rect 280846 627912 280906 627950
rect 281533 627947 281599 627950
rect 476062 627812 476068 627876
rect 476132 627874 476138 627876
rect 477125 627874 477191 627877
rect 476132 627872 477191 627874
rect 476132 627816 477130 627872
rect 477186 627816 477191 627872
rect 476132 627814 477191 627816
rect 476132 627812 476138 627814
rect 477125 627811 477191 627814
rect 488574 627812 488580 627876
rect 488644 627874 488650 627876
rect 488717 627874 488783 627877
rect 488644 627872 488783 627874
rect 488644 627816 488722 627872
rect 488778 627816 488783 627872
rect 488644 627814 488783 627816
rect 488644 627812 488650 627814
rect 488717 627811 488783 627814
rect 506606 627812 506612 627876
rect 506676 627874 506682 627876
rect 506749 627874 506815 627877
rect 506676 627872 506815 627874
rect 506676 627816 506754 627872
rect 506810 627816 506815 627872
rect 506676 627814 506815 627816
rect 506676 627812 506682 627814
rect 506749 627811 506815 627814
rect 456793 627738 456859 627741
rect 456793 627736 460092 627738
rect 456793 627680 456798 627736
rect 456854 627680 460092 627736
rect 456793 627678 460092 627680
rect 456793 627675 456859 627678
rect 59169 625834 59235 625837
rect 59494 625834 60076 625870
rect 59169 625832 60076 625834
rect 59169 625776 59174 625832
rect 59230 625810 60076 625832
rect 139025 625834 139091 625837
rect 139534 625834 140116 625870
rect 139025 625832 140116 625834
rect 59230 625776 59554 625810
rect 59169 625774 59554 625776
rect 139025 625776 139030 625832
rect 139086 625810 140116 625832
rect 216673 625834 216739 625837
rect 219758 625834 220156 625870
rect 216673 625832 220156 625834
rect 139086 625776 139594 625810
rect 139025 625774 139594 625776
rect 216673 625776 216678 625832
rect 216734 625810 220156 625832
rect 216734 625776 219818 625810
rect 216673 625774 219818 625776
rect 59169 625771 59235 625774
rect 139025 625771 139091 625774
rect 216673 625771 216739 625774
rect 121545 625290 121611 625293
rect 202965 625290 203031 625293
rect 282913 625290 282979 625293
rect 120766 625288 121611 625290
rect 120766 625232 121550 625288
rect 121606 625232 121611 625288
rect 120766 625230 121611 625232
rect 120766 625192 120826 625230
rect 121545 625227 121611 625230
rect 200806 625288 203031 625290
rect 200806 625232 202970 625288
rect 203026 625232 203031 625288
rect 200806 625230 203031 625232
rect 200806 625192 200866 625230
rect 202965 625227 203031 625230
rect 280846 625288 282979 625290
rect 280846 625232 282918 625288
rect 282974 625232 282979 625288
rect 280846 625230 282979 625232
rect 280846 625192 280906 625230
rect 282913 625227 282979 625230
rect 512085 625018 512151 625021
rect 509956 625016 512151 625018
rect 509956 624960 512090 625016
rect 512146 624960 512151 625016
rect 509956 624958 512151 624960
rect 512085 624955 512151 624958
rect 430665 624610 430731 624613
rect 428812 624608 430731 624610
rect 428812 624552 430670 624608
rect 430726 624552 430731 624608
rect 428812 624550 430731 624552
rect 430665 624547 430731 624550
rect 317413 623930 317479 623933
rect 317413 623928 320068 623930
rect 317413 623872 317418 623928
rect 317474 623872 320068 623928
rect 317413 623870 320068 623872
rect 317413 623867 317479 623870
rect 57697 622434 57763 622437
rect 59494 622434 60076 622470
rect 57697 622432 60076 622434
rect 57697 622376 57702 622432
rect 57758 622410 60076 622432
rect 139301 622434 139367 622437
rect 139534 622434 140116 622470
rect 139301 622432 140116 622434
rect 57758 622376 59554 622410
rect 57697 622374 59554 622376
rect 139301 622376 139306 622432
rect 139362 622410 140116 622432
rect 217685 622434 217751 622437
rect 219758 622434 220156 622470
rect 217685 622432 220156 622434
rect 139362 622376 139594 622410
rect 139301 622374 139594 622376
rect 217685 622376 217690 622432
rect 217746 622410 220156 622432
rect 217746 622376 219818 622410
rect 217685 622374 219818 622376
rect 57697 622371 57763 622374
rect 139301 622371 139367 622374
rect 217685 622371 217751 622374
rect 120766 621210 120826 621792
rect 121821 621210 121887 621213
rect 120766 621208 121887 621210
rect 120766 621152 121826 621208
rect 121882 621152 121887 621208
rect 120766 621150 121887 621152
rect 200806 621210 200866 621792
rect 202229 621210 202295 621213
rect 200806 621208 202295 621210
rect 200806 621152 202234 621208
rect 202290 621152 202295 621208
rect 200806 621150 202295 621152
rect 280846 621210 280906 621792
rect 457529 621618 457595 621621
rect 457529 621616 460092 621618
rect 457529 621560 457534 621616
rect 457590 621560 460092 621616
rect 457529 621558 460092 621560
rect 457529 621555 457595 621558
rect 283005 621210 283071 621213
rect 280846 621208 283071 621210
rect 280846 621152 283010 621208
rect 283066 621152 283071 621208
rect 280846 621150 283071 621152
rect 121821 621147 121887 621150
rect 202229 621147 202295 621150
rect 283005 621147 283071 621150
rect 430849 619850 430915 619853
rect 428812 619848 430915 619850
rect 428812 619792 430854 619848
rect 430910 619792 430915 619848
rect 428812 619790 430915 619792
rect 430849 619787 430915 619790
rect 57513 619714 57579 619717
rect 59494 619714 60076 619750
rect 57513 619712 60076 619714
rect 57513 619656 57518 619712
rect 57574 619690 60076 619712
rect 137553 619714 137619 619717
rect 139534 619714 140116 619750
rect 137553 619712 140116 619714
rect 57574 619656 59554 619690
rect 57513 619654 59554 619656
rect 137553 619656 137558 619712
rect 137614 619690 140116 619712
rect 216673 619714 216739 619717
rect 219758 619714 220156 619750
rect 216673 619712 220156 619714
rect 137614 619656 139594 619690
rect 137553 619654 139594 619656
rect 216673 619656 216678 619712
rect 216734 619690 220156 619712
rect 216734 619656 219818 619690
rect 216673 619654 219818 619656
rect 57513 619651 57579 619654
rect 137553 619651 137619 619654
rect 216673 619651 216739 619654
rect -960 619020 480 619260
rect 317597 619170 317663 619173
rect 317597 619168 320068 619170
rect 317597 619112 317602 619168
rect 317658 619112 320068 619168
rect 317597 619110 320068 619112
rect 317597 619107 317663 619110
rect 120766 618490 120826 619072
rect 200806 618493 200866 619072
rect 121913 618490 121979 618493
rect 120766 618488 121979 618490
rect 120766 618432 121918 618488
rect 121974 618432 121979 618488
rect 120766 618430 121979 618432
rect 121913 618427 121979 618430
rect 200757 618488 200866 618493
rect 200757 618432 200762 618488
rect 200818 618432 200866 618488
rect 200757 618430 200866 618432
rect 280846 618490 280906 619072
rect 510613 618898 510679 618901
rect 509956 618896 510679 618898
rect 509956 618840 510618 618896
rect 510674 618840 510679 618896
rect 509956 618838 510679 618840
rect 510613 618835 510679 618838
rect 281625 618490 281691 618493
rect 280846 618488 281691 618490
rect 280846 618432 281630 618488
rect 281686 618432 281691 618488
rect 280846 618430 281691 618432
rect 200757 618427 200823 618430
rect 281625 618427 281691 618430
rect 583520 617388 584960 617628
rect 58617 616314 58683 616317
rect 59494 616314 60076 616350
rect 58617 616312 60076 616314
rect 58617 616256 58622 616312
rect 58678 616290 60076 616312
rect 136725 616314 136791 616317
rect 139534 616314 140116 616350
rect 136725 616312 140116 616314
rect 58678 616256 59554 616290
rect 58617 616254 59554 616256
rect 136725 616256 136730 616312
rect 136786 616290 140116 616312
rect 216673 616314 216739 616317
rect 219758 616314 220156 616350
rect 216673 616312 220156 616314
rect 136786 616256 139594 616290
rect 136725 616254 139594 616256
rect 216673 616256 216678 616312
rect 216734 616290 220156 616312
rect 216734 616256 219818 616290
rect 216673 616254 219818 616256
rect 58617 616251 58683 616254
rect 136725 616251 136791 616254
rect 216673 616251 216739 616254
rect 120766 615634 120826 615672
rect 121729 615634 121795 615637
rect 120766 615632 121795 615634
rect 120766 615576 121734 615632
rect 121790 615576 121795 615632
rect 120766 615574 121795 615576
rect 200806 615634 200866 615672
rect 202873 615634 202939 615637
rect 200806 615632 202939 615634
rect 200806 615576 202878 615632
rect 202934 615576 202939 615632
rect 200806 615574 202939 615576
rect 280846 615634 280906 615672
rect 281717 615634 281783 615637
rect 280846 615632 281783 615634
rect 280846 615576 281722 615632
rect 281778 615576 281783 615632
rect 280846 615574 281783 615576
rect 121729 615571 121795 615574
rect 202873 615571 202939 615574
rect 281717 615571 281783 615574
rect 457621 615498 457687 615501
rect 457621 615496 460092 615498
rect 457621 615440 457626 615496
rect 457682 615440 460092 615496
rect 457621 615438 460092 615440
rect 457621 615435 457687 615438
rect 430614 615090 430620 615092
rect 428812 615030 430620 615090
rect 430614 615028 430620 615030
rect 430684 615028 430690 615092
rect 317965 614410 318031 614413
rect 317965 614408 320068 614410
rect 317965 614352 317970 614408
rect 318026 614352 320068 614408
rect 317965 614350 320068 614352
rect 317965 614347 318031 614350
rect 57605 613594 57671 613597
rect 59494 613594 60076 613630
rect 57605 613592 60076 613594
rect 57605 613536 57610 613592
rect 57666 613570 60076 613592
rect 138933 613594 138999 613597
rect 139534 613594 140116 613630
rect 138933 613592 140116 613594
rect 57666 613536 59554 613570
rect 57605 613534 59554 613536
rect 138933 613536 138938 613592
rect 138994 613570 140116 613592
rect 219249 613594 219315 613597
rect 219758 613594 220156 613630
rect 219249 613592 220156 613594
rect 138994 613536 139594 613570
rect 138933 613534 139594 613536
rect 219249 613536 219254 613592
rect 219310 613570 220156 613592
rect 219310 613536 219818 613570
rect 219249 613534 219818 613536
rect 57605 613531 57671 613534
rect 138933 613531 138999 613534
rect 219249 613531 219315 613534
rect 120766 612778 120826 612952
rect 123109 612778 123175 612781
rect 120766 612776 123175 612778
rect 120766 612720 123114 612776
rect 123170 612720 123175 612776
rect 120766 612718 123175 612720
rect 200806 612778 200866 612952
rect 201861 612778 201927 612781
rect 200806 612776 201927 612778
rect 200806 612720 201866 612776
rect 201922 612720 201927 612776
rect 200806 612718 201927 612720
rect 280846 612778 280906 612952
rect 281809 612778 281875 612781
rect 280846 612776 281875 612778
rect 280846 612720 281814 612776
rect 281870 612720 281875 612776
rect 280846 612718 281875 612720
rect 123109 612715 123175 612718
rect 201861 612715 201927 612718
rect 281809 612715 281875 612718
rect 511993 612098 512059 612101
rect 509956 612096 512059 612098
rect 509956 612040 511998 612096
rect 512054 612040 512059 612096
rect 509956 612038 512059 612040
rect 511993 612035 512059 612038
rect 430573 610330 430639 610333
rect 428812 610328 430639 610330
rect 428812 610272 430578 610328
rect 430634 610272 430639 610328
rect 428812 610270 430639 610272
rect 430573 610267 430639 610270
rect 58893 610194 58959 610197
rect 59494 610194 60076 610230
rect 58893 610192 60076 610194
rect 58893 610136 58898 610192
rect 58954 610170 60076 610192
rect 138841 610194 138907 610197
rect 139534 610194 140116 610230
rect 138841 610192 140116 610194
rect 58954 610136 59554 610170
rect 58893 610134 59554 610136
rect 138841 610136 138846 610192
rect 138902 610170 140116 610192
rect 217777 610194 217843 610197
rect 219758 610194 220156 610230
rect 217777 610192 220156 610194
rect 138902 610136 139594 610170
rect 138841 610134 139594 610136
rect 217777 610136 217782 610192
rect 217838 610170 220156 610192
rect 217838 610136 219818 610170
rect 217777 610134 219818 610136
rect 58893 610131 58959 610134
rect 138841 610131 138907 610134
rect 217777 610131 217843 610134
rect 317965 609650 318031 609653
rect 317965 609648 320068 609650
rect 317965 609592 317970 609648
rect 318026 609592 320068 609648
rect 317965 609590 320068 609592
rect 317965 609587 318031 609590
rect 120766 608973 120826 609552
rect 120766 608968 120875 608973
rect 120766 608912 120814 608968
rect 120870 608912 120875 608968
rect 120766 608910 120875 608912
rect 200806 608970 200866 609552
rect 201953 608970 202019 608973
rect 200806 608968 202019 608970
rect 200806 608912 201958 608968
rect 202014 608912 202019 608968
rect 200806 608910 202019 608912
rect 280846 608970 280906 609552
rect 457713 609378 457779 609381
rect 457713 609376 460092 609378
rect 457713 609320 457718 609376
rect 457774 609320 460092 609376
rect 457713 609318 460092 609320
rect 457713 609315 457779 609318
rect 283097 608970 283163 608973
rect 280846 608968 283163 608970
rect 280846 608912 283102 608968
rect 283158 608912 283163 608968
rect 280846 608910 283163 608912
rect 120809 608907 120875 608910
rect 201953 608907 202019 608910
rect 283097 608907 283163 608910
rect 59077 607610 59143 607613
rect 137737 607610 137803 607613
rect 219157 607610 219223 607613
rect 59077 607608 59554 607610
rect 59077 607552 59082 607608
rect 59138 607566 59554 607608
rect 137737 607608 139410 607610
rect 59138 607552 60076 607566
rect 59077 607550 60076 607552
rect 59077 607547 59143 607550
rect 59494 607506 60076 607550
rect 137737 607552 137742 607608
rect 137798 607552 139410 607608
rect 137737 607550 139410 607552
rect 137737 607547 137803 607550
rect 139350 607542 139410 607550
rect 219157 607608 219450 607610
rect 219157 607552 219162 607608
rect 219218 607552 219450 607608
rect 219157 607550 219450 607552
rect 219157 607547 219223 607550
rect 219390 607542 219450 607550
rect 139350 607482 140032 607542
rect 219390 607482 220064 607542
rect 120766 606250 120826 606832
rect 200806 606386 200866 606832
rect 203149 606386 203215 606389
rect 200806 606384 203215 606386
rect 200806 606328 203154 606384
rect 203210 606328 203215 606384
rect 200806 606326 203215 606328
rect 280846 606386 280906 606832
rect 283281 606386 283347 606389
rect 280846 606384 283347 606386
rect 280846 606328 283286 606384
rect 283342 606328 283347 606384
rect 280846 606326 283347 606328
rect 203149 606323 203215 606326
rect 283281 606323 283347 606326
rect 123293 606250 123359 606253
rect 120766 606248 123359 606250
rect -960 605964 480 606204
rect 120766 606192 123298 606248
rect 123354 606192 123359 606248
rect 120766 606190 123359 606192
rect 123293 606187 123359 606190
rect 511993 605978 512059 605981
rect 509956 605976 512059 605978
rect 509956 605920 511998 605976
rect 512054 605920 512059 605976
rect 509956 605918 512059 605920
rect 511993 605915 512059 605918
rect 430665 605570 430731 605573
rect 428812 605568 430731 605570
rect 428812 605512 430670 605568
rect 430726 605512 430731 605568
rect 428812 605510 430731 605512
rect 430665 605507 430731 605510
rect 317965 604890 318031 604893
rect 317965 604888 320068 604890
rect 317965 604832 317970 604888
rect 318026 604832 320068 604888
rect 317965 604830 320068 604832
rect 317965 604827 318031 604830
rect 218697 604210 218763 604213
rect 218697 604208 219450 604210
rect 218697 604152 218702 604208
rect 218758 604152 219450 604208
rect 218697 604150 219450 604152
rect 218697 604147 218763 604150
rect 219390 604142 219450 604150
rect 57881 604074 57947 604077
rect 59494 604074 60076 604110
rect 57881 604072 60076 604074
rect 57881 604016 57886 604072
rect 57942 604050 60076 604072
rect 137921 604074 137987 604077
rect 139534 604074 140116 604116
rect 219390 604082 220064 604142
rect 137921 604072 140116 604074
rect 57942 604016 59554 604050
rect 57881 604014 59554 604016
rect 137921 604016 137926 604072
rect 137982 604056 140116 604072
rect 583520 604060 584960 604300
rect 137982 604016 139594 604056
rect 137921 604014 139594 604016
rect 57881 604011 57947 604014
rect 137921 604011 137987 604014
rect 120766 603122 120826 603432
rect 123201 603122 123267 603125
rect 120766 603120 123267 603122
rect 120766 603064 123206 603120
rect 123262 603064 123267 603120
rect 120766 603062 123267 603064
rect 200806 603122 200866 603432
rect 203057 603122 203123 603125
rect 200806 603120 203123 603122
rect 200806 603064 203062 603120
rect 203118 603064 203123 603120
rect 200806 603062 203123 603064
rect 280846 603122 280906 603432
rect 283189 603122 283255 603125
rect 280846 603120 283255 603122
rect 280846 603064 283194 603120
rect 283250 603064 283255 603120
rect 280846 603062 283255 603064
rect 123201 603059 123267 603062
rect 203057 603059 203123 603062
rect 283189 603059 283255 603062
rect 457805 602578 457871 602581
rect 457805 602576 460092 602578
rect 457805 602520 457810 602576
rect 457866 602520 460092 602576
rect 457805 602518 460092 602520
rect 457805 602515 457871 602518
rect 58801 601354 58867 601357
rect 59494 601354 60076 601390
rect 58801 601352 60076 601354
rect 58801 601296 58806 601352
rect 58862 601330 60076 601352
rect 137921 601354 137987 601357
rect 139534 601354 140116 601390
rect 137921 601352 140116 601354
rect 58862 601296 59554 601330
rect 58801 601294 59554 601296
rect 137921 601296 137926 601352
rect 137982 601330 140116 601352
rect 217409 601354 217475 601357
rect 219758 601354 220156 601390
rect 217409 601352 220156 601354
rect 137982 601296 139594 601330
rect 137921 601294 139594 601296
rect 217409 601296 217414 601352
rect 217470 601330 220156 601352
rect 217470 601296 219818 601330
rect 217409 601294 219818 601296
rect 58801 601291 58867 601294
rect 137921 601291 137987 601294
rect 217409 601291 217475 601294
rect 430798 600810 430804 600812
rect 428812 600750 430804 600810
rect 430798 600748 430804 600750
rect 430868 600748 430874 600812
rect 120766 600402 120826 600712
rect 122005 600402 122071 600405
rect 120766 600400 122071 600402
rect 120766 600344 122010 600400
rect 122066 600344 122071 600400
rect 120766 600342 122071 600344
rect 200806 600402 200866 600712
rect 280846 600405 280906 600712
rect 202045 600402 202111 600405
rect 200806 600400 202111 600402
rect 200806 600344 202050 600400
rect 202106 600344 202111 600400
rect 200806 600342 202111 600344
rect 280846 600400 280955 600405
rect 280846 600344 280894 600400
rect 280950 600344 280955 600400
rect 280846 600342 280955 600344
rect 122005 600339 122071 600342
rect 202045 600339 202111 600342
rect 280889 600339 280955 600342
rect 318793 600130 318859 600133
rect 318793 600128 320068 600130
rect 318793 600072 318798 600128
rect 318854 600072 320068 600128
rect 318793 600070 320068 600072
rect 318793 600067 318859 600070
rect 512177 599858 512243 599861
rect 509956 599856 512243 599858
rect 509956 599800 512182 599856
rect 512238 599800 512243 599856
rect 509956 599798 512243 599800
rect 512177 599795 512243 599798
rect 58709 597954 58775 597957
rect 59494 597954 60076 597990
rect 58709 597952 60076 597954
rect 58709 597896 58714 597952
rect 58770 597930 60076 597952
rect 136725 597954 136791 597957
rect 139534 597954 140116 597990
rect 136725 597952 140116 597954
rect 58770 597896 59554 597930
rect 58709 597894 59554 597896
rect 136725 597896 136730 597952
rect 136786 597930 140116 597952
rect 216673 597954 216739 597957
rect 219758 597954 220156 597990
rect 216673 597952 220156 597954
rect 136786 597896 139594 597930
rect 136725 597894 139594 597896
rect 216673 597896 216678 597952
rect 216734 597930 220156 597952
rect 216734 597896 219818 597930
rect 216673 597894 219818 597896
rect 58709 597891 58775 597894
rect 136725 597891 136791 597894
rect 216673 597891 216739 597894
rect 120766 596730 120826 597312
rect 124121 596730 124187 596733
rect 120766 596728 124187 596730
rect 120766 596672 124126 596728
rect 124182 596672 124187 596728
rect 120766 596670 124187 596672
rect 200806 596730 200866 597312
rect 203241 596730 203307 596733
rect 200806 596728 203307 596730
rect 200806 596672 203246 596728
rect 203302 596672 203307 596728
rect 200806 596670 203307 596672
rect 280846 596730 280906 597312
rect 283649 596730 283715 596733
rect 280846 596728 283715 596730
rect 280846 596672 283654 596728
rect 283710 596672 283715 596728
rect 280846 596670 283715 596672
rect 124121 596667 124187 596670
rect 203241 596667 203307 596670
rect 283649 596667 283715 596670
rect 457529 596458 457595 596461
rect 457529 596456 460092 596458
rect 457529 596400 457534 596456
rect 457590 596400 460092 596456
rect 457529 596398 460092 596400
rect 457529 596395 457595 596398
rect 429469 596050 429535 596053
rect 428812 596048 429535 596050
rect 428812 595992 429474 596048
rect 429530 595992 429535 596048
rect 428812 595990 429535 595992
rect 429469 595987 429535 595990
rect 317965 595370 318031 595373
rect 317965 595368 320068 595370
rect 317965 595312 317970 595368
rect 318026 595312 320068 595368
rect 317965 595310 320068 595312
rect 317965 595307 318031 595310
rect 57237 595234 57303 595237
rect 59494 595234 60076 595270
rect 57237 595232 60076 595234
rect 57237 595176 57242 595232
rect 57298 595210 60076 595232
rect 137369 595234 137435 595237
rect 139534 595234 140116 595270
rect 137369 595232 140116 595234
rect 57298 595176 59554 595210
rect 57237 595174 59554 595176
rect 137369 595176 137374 595232
rect 137430 595210 140116 595232
rect 216673 595234 216739 595237
rect 219758 595234 220156 595270
rect 216673 595232 220156 595234
rect 137430 595176 139594 595210
rect 137369 595174 139594 595176
rect 216673 595176 216678 595232
rect 216734 595210 220156 595232
rect 216734 595176 219818 595210
rect 216673 595174 219818 595176
rect 57237 595171 57303 595174
rect 137369 595171 137435 595174
rect 216673 595171 216739 595174
rect 201033 594622 201099 594625
rect 200836 594620 201099 594622
rect 120766 594010 120826 594592
rect 200836 594564 201038 594620
rect 201094 594564 201099 594620
rect 200836 594562 201099 594564
rect 201033 594559 201099 594562
rect 123385 594010 123451 594013
rect 120766 594008 123451 594010
rect 120766 593952 123390 594008
rect 123446 593952 123451 594008
rect 120766 593950 123451 593952
rect 280846 594010 280906 594592
rect 281901 594010 281967 594013
rect 280846 594008 281967 594010
rect 280846 593952 281906 594008
rect 281962 593952 281967 594008
rect 280846 593950 281967 593952
rect 123385 593947 123451 593950
rect 281901 593947 281967 593950
rect 512085 593738 512151 593741
rect 509956 593736 512151 593738
rect 509956 593680 512090 593736
rect 512146 593680 512151 593736
rect 509956 593678 512151 593680
rect 512085 593675 512151 593678
rect -960 592908 480 593148
rect 57421 591834 57487 591837
rect 59494 591834 60076 591870
rect 57421 591832 60076 591834
rect 57421 591776 57426 591832
rect 57482 591810 60076 591832
rect 137737 591834 137803 591837
rect 139534 591834 140116 591870
rect 137737 591832 140116 591834
rect 57482 591776 59554 591810
rect 57421 591774 59554 591776
rect 137737 591776 137742 591832
rect 137798 591810 140116 591832
rect 216673 591834 216739 591837
rect 219758 591834 220156 591870
rect 216673 591832 220156 591834
rect 137798 591776 139594 591810
rect 137737 591774 139594 591776
rect 216673 591776 216678 591832
rect 216734 591810 220156 591832
rect 216734 591776 219818 591810
rect 216673 591774 219818 591776
rect 57421 591771 57487 591774
rect 137737 591771 137803 591774
rect 216673 591771 216739 591774
rect 429285 591290 429351 591293
rect 428812 591288 429351 591290
rect 428812 591232 429290 591288
rect 429346 591232 429351 591288
rect 428812 591230 429351 591232
rect 429285 591227 429351 591230
rect 121085 591222 121151 591225
rect 120796 591220 121151 591222
rect 120796 591164 121090 591220
rect 121146 591164 121151 591220
rect 120796 591162 121151 591164
rect 121085 591159 121151 591162
rect 200806 590746 200866 591192
rect 202137 590746 202203 590749
rect 200806 590744 202203 590746
rect 200806 590688 202142 590744
rect 202198 590688 202203 590744
rect 200806 590686 202203 590688
rect 280846 590746 280906 591192
rect 583520 590868 584960 591108
rect 283373 590746 283439 590749
rect 280846 590744 283439 590746
rect 280846 590688 283378 590744
rect 283434 590688 283439 590744
rect 280846 590686 283439 590688
rect 202137 590683 202203 590686
rect 283373 590683 283439 590686
rect 317965 590610 318031 590613
rect 317965 590608 320068 590610
rect 317965 590552 317970 590608
rect 318026 590552 320068 590608
rect 317965 590550 320068 590552
rect 317965 590547 318031 590550
rect 457437 590338 457503 590341
rect 457437 590336 460092 590338
rect 457437 590280 457442 590336
rect 457498 590280 460092 590336
rect 457437 590278 460092 590280
rect 457437 590275 457503 590278
rect 57145 589114 57211 589117
rect 59494 589114 60076 589150
rect 57145 589112 60076 589114
rect 57145 589056 57150 589112
rect 57206 589090 60076 589112
rect 138749 589114 138815 589117
rect 139534 589114 140116 589150
rect 138749 589112 140116 589114
rect 57206 589056 59554 589090
rect 57145 589054 59554 589056
rect 138749 589056 138754 589112
rect 138810 589090 140116 589112
rect 217593 589114 217659 589117
rect 219758 589114 220156 589150
rect 217593 589112 220156 589114
rect 138810 589056 139594 589090
rect 138749 589054 139594 589056
rect 217593 589056 217598 589112
rect 217654 589090 220156 589112
rect 217654 589056 219818 589090
rect 217593 589054 219818 589056
rect 57145 589051 57211 589054
rect 138749 589051 138815 589054
rect 217593 589051 217659 589054
rect 120766 588026 120826 588472
rect 122097 588026 122163 588029
rect 120766 588024 122163 588026
rect 120766 587968 122102 588024
rect 122158 587968 122163 588024
rect 120766 587966 122163 587968
rect 200806 588026 200866 588472
rect 203241 588026 203307 588029
rect 200806 588024 203307 588026
rect 200806 587968 203246 588024
rect 203302 587968 203307 588024
rect 200806 587966 203307 587968
rect 280846 588026 280906 588472
rect 283465 588026 283531 588029
rect 280846 588024 283531 588026
rect 280846 587968 283470 588024
rect 283526 587968 283531 588024
rect 280846 587966 283531 587968
rect 122097 587963 122163 587966
rect 203241 587963 203307 587966
rect 283465 587963 283531 587966
rect 512269 587618 512335 587621
rect 509956 587616 512335 587618
rect 509956 587560 512274 587616
rect 512330 587560 512335 587616
rect 509956 587558 512335 587560
rect 512269 587555 512335 587558
rect 429561 586666 429627 586669
rect 428782 586664 429627 586666
rect 428782 586608 429566 586664
rect 429622 586608 429627 586664
rect 428782 586606 429627 586608
rect 428782 586500 428842 586606
rect 429561 586603 429627 586606
rect 317965 585850 318031 585853
rect 317965 585848 320068 585850
rect 317965 585792 317970 585848
rect 318026 585792 320068 585848
rect 317965 585790 320068 585792
rect 317965 585787 318031 585790
rect 58525 585714 58591 585717
rect 59494 585714 60076 585750
rect 58525 585712 60076 585714
rect 58525 585656 58530 585712
rect 58586 585690 60076 585712
rect 136725 585714 136791 585717
rect 139534 585714 140116 585750
rect 136725 585712 140116 585714
rect 58586 585656 59554 585690
rect 58525 585654 59554 585656
rect 136725 585656 136730 585712
rect 136786 585690 140116 585712
rect 216029 585714 216095 585717
rect 219758 585714 220156 585750
rect 216029 585712 220156 585714
rect 136786 585656 139594 585690
rect 136725 585654 139594 585656
rect 216029 585656 216034 585712
rect 216090 585690 220156 585712
rect 216090 585656 219818 585690
rect 216029 585654 219818 585656
rect 58525 585651 58591 585654
rect 136725 585651 136791 585654
rect 216029 585651 216095 585654
rect 120766 584490 120826 585072
rect 123477 584490 123543 584493
rect 120766 584488 123543 584490
rect 120766 584432 123482 584488
rect 123538 584432 123543 584488
rect 120766 584430 123543 584432
rect 200806 584490 200866 585072
rect 201493 584490 201559 584493
rect 200806 584488 201559 584490
rect 200806 584432 201498 584488
rect 201554 584432 201559 584488
rect 200806 584430 201559 584432
rect 280846 584490 280906 585072
rect 281993 584490 282059 584493
rect 280846 584488 282059 584490
rect 280846 584432 281998 584488
rect 282054 584432 282059 584488
rect 280846 584430 282059 584432
rect 123477 584427 123543 584430
rect 201493 584427 201559 584430
rect 281993 584427 282059 584430
rect 457437 584218 457503 584221
rect 457437 584216 460092 584218
rect 457437 584160 457442 584216
rect 457498 584160 460092 584216
rect 457437 584158 460092 584160
rect 457437 584155 457503 584158
rect 59077 582994 59143 582997
rect 59494 582994 60076 583030
rect 59077 582992 60076 582994
rect 59077 582936 59082 582992
rect 59138 582970 60076 582992
rect 136725 582994 136791 582997
rect 139534 582994 140116 583030
rect 136725 582992 140116 582994
rect 59138 582936 59554 582970
rect 59077 582934 59554 582936
rect 136725 582936 136730 582992
rect 136786 582970 140116 582992
rect 216673 582994 216739 582997
rect 219758 582994 220156 583030
rect 216673 582992 220156 582994
rect 136786 582936 139594 582970
rect 136725 582934 139594 582936
rect 216673 582936 216678 582992
rect 216734 582970 220156 582992
rect 216734 582936 219818 582970
rect 216673 582934 219818 582936
rect 59077 582931 59143 582934
rect 136725 582931 136791 582934
rect 216673 582931 216739 582934
rect 120766 581770 120826 582352
rect 122189 581770 122255 581773
rect 120766 581768 122255 581770
rect 120766 581712 122194 581768
rect 122250 581712 122255 581768
rect 120766 581710 122255 581712
rect 200806 581770 200866 582352
rect 203333 581770 203399 581773
rect 200806 581768 203399 581770
rect 200806 581712 203338 581768
rect 203394 581712 203399 581768
rect 200806 581710 203399 581712
rect 280846 581770 280906 582352
rect 282085 581770 282151 581773
rect 280846 581768 282151 581770
rect 280846 581712 282090 581768
rect 282146 581712 282151 581768
rect 280846 581710 282151 581712
rect 122189 581707 122255 581710
rect 203333 581707 203399 581710
rect 282085 581707 282151 581710
rect 430757 581090 430823 581093
rect 428812 581088 430823 581090
rect 428812 581032 430762 581088
rect 430818 581032 430823 581088
rect 428812 581030 430823 581032
rect 430757 581027 430823 581030
rect 513005 580818 513071 580821
rect 509956 580816 513071 580818
rect 509956 580760 513010 580816
rect 513066 580760 513071 580816
rect 509956 580758 513071 580760
rect 513005 580755 513071 580758
rect 317965 580410 318031 580413
rect 317965 580408 320068 580410
rect 317965 580352 317970 580408
rect 318026 580352 320068 580408
rect 317965 580350 320068 580352
rect 317965 580347 318031 580350
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 57329 579730 57395 579733
rect 137461 579730 137527 579733
rect 216673 579730 216739 579733
rect 57329 579728 59554 579730
rect 57329 579672 57334 579728
rect 57390 579686 59554 579728
rect 137461 579728 139410 579730
rect 57390 579672 60076 579686
rect 57329 579670 60076 579672
rect 57329 579667 57395 579670
rect 59494 579626 60076 579670
rect 137461 579672 137466 579728
rect 137522 579672 139410 579728
rect 137461 579670 139410 579672
rect 137461 579667 137527 579670
rect 139350 579662 139410 579670
rect 216673 579728 219450 579730
rect 216673 579672 216678 579728
rect 216734 579672 219450 579728
rect 216673 579670 219450 579672
rect 216673 579667 216739 579670
rect 219390 579662 219450 579670
rect 139350 579602 140032 579662
rect 219390 579602 220064 579662
rect 120766 578370 120826 578952
rect 122281 578370 122347 578373
rect 120766 578368 122347 578370
rect 120766 578312 122286 578368
rect 122342 578312 122347 578368
rect 120766 578310 122347 578312
rect 200806 578370 200866 578952
rect 202321 578370 202387 578373
rect 200806 578368 202387 578370
rect 200806 578312 202326 578368
rect 202382 578312 202387 578368
rect 200806 578310 202387 578312
rect 280846 578370 280906 578952
rect 283557 578370 283623 578373
rect 280846 578368 283623 578370
rect 280846 578312 283562 578368
rect 283618 578312 283623 578368
rect 280846 578310 283623 578312
rect 122281 578307 122347 578310
rect 202321 578307 202387 578310
rect 283557 578307 283623 578310
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect 57053 576874 57119 576877
rect 59494 576874 60076 576910
rect 57053 576872 60076 576874
rect 57053 576816 57058 576872
rect 57114 576850 60076 576872
rect 138657 576874 138723 576877
rect 139534 576874 140116 576910
rect 138657 576872 140116 576874
rect 57114 576816 59554 576850
rect 57053 576814 59554 576816
rect 138657 576816 138662 576872
rect 138718 576850 140116 576872
rect 219157 576874 219223 576877
rect 219758 576874 220156 576910
rect 219157 576872 220156 576874
rect 138718 576816 139594 576850
rect 138657 576814 139594 576816
rect 219157 576816 219162 576872
rect 219218 576850 220156 576872
rect 219218 576816 219818 576850
rect 219157 576814 219818 576816
rect 57053 576811 57119 576814
rect 138657 576811 138723 576814
rect 219157 576811 219223 576814
rect 430849 576330 430915 576333
rect 428812 576328 430915 576330
rect 428812 576272 430854 576328
rect 430910 576272 430915 576328
rect 428812 576270 430915 576272
rect 430849 576267 430915 576270
rect 201125 576262 201191 576265
rect 200836 576260 201191 576262
rect 120766 575650 120826 576232
rect 200836 576204 201130 576260
rect 201186 576204 201191 576260
rect 200836 576202 201191 576204
rect 201125 576199 201191 576202
rect 123661 575650 123727 575653
rect 120766 575648 123727 575650
rect 120766 575592 123666 575648
rect 123722 575592 123727 575648
rect 120766 575590 123727 575592
rect 280846 575650 280906 576232
rect 282177 575650 282243 575653
rect 280846 575648 282243 575650
rect 280846 575592 282182 575648
rect 282238 575592 282243 575648
rect 280846 575590 282243 575592
rect 123661 575587 123727 575590
rect 282177 575587 282243 575590
rect 316769 575650 316835 575653
rect 316769 575648 320068 575650
rect 316769 575592 316774 575648
rect 316830 575592 320068 575648
rect 316769 575590 320068 575592
rect 316769 575587 316835 575590
rect 58433 573474 58499 573477
rect 59494 573474 60076 573510
rect 58433 573472 60076 573474
rect 58433 573416 58438 573472
rect 58494 573450 60076 573472
rect 137185 573474 137251 573477
rect 139534 573474 140116 573510
rect 137185 573472 140116 573474
rect 58494 573416 59554 573450
rect 58433 573414 59554 573416
rect 137185 573416 137190 573472
rect 137246 573450 140116 573472
rect 217501 573474 217567 573477
rect 219758 573474 220156 573510
rect 217501 573472 220156 573474
rect 137246 573416 139594 573450
rect 137185 573414 139594 573416
rect 217501 573416 217506 573472
rect 217562 573450 220156 573472
rect 217562 573416 219818 573450
rect 217501 573414 219818 573416
rect 58433 573411 58499 573414
rect 137185 573411 137251 573414
rect 217501 573411 217567 573414
rect 121177 572862 121243 572865
rect 281165 572862 281231 572865
rect 120796 572860 121243 572862
rect 120796 572804 121182 572860
rect 121238 572804 121243 572860
rect 280876 572860 281231 572862
rect 120796 572802 121243 572804
rect 121177 572799 121243 572802
rect 200806 572794 200866 572832
rect 280876 572804 281170 572860
rect 281226 572804 281231 572860
rect 280876 572802 281231 572804
rect 281165 572799 281231 572802
rect 203425 572794 203491 572797
rect 200806 572792 203491 572794
rect 200806 572736 203430 572792
rect 203486 572736 203491 572792
rect 200806 572734 203491 572736
rect 203425 572731 203491 572734
rect 430941 571570 431007 571573
rect 428812 571568 431007 571570
rect 428812 571512 430946 571568
rect 431002 571512 431007 571568
rect 428812 571510 431007 571512
rect 430941 571507 431007 571510
rect 316769 570890 316835 570893
rect 316769 570888 320068 570890
rect 316769 570832 316774 570888
rect 316830 570832 320068 570888
rect 316769 570830 320068 570832
rect 316769 570827 316835 570830
rect 59537 570790 59603 570793
rect 59537 570788 60076 570790
rect 59537 570732 59542 570788
rect 59598 570732 60076 570788
rect 59537 570730 60076 570732
rect 139209 570754 139275 570757
rect 139534 570754 140116 570790
rect 139209 570752 140116 570754
rect 59537 570727 59603 570730
rect 139209 570696 139214 570752
rect 139270 570730 140116 570752
rect 216673 570754 216739 570757
rect 219758 570754 220156 570790
rect 216673 570752 220156 570754
rect 139270 570696 139594 570730
rect 139209 570694 139594 570696
rect 216673 570696 216678 570752
rect 216734 570730 220156 570752
rect 216734 570696 219818 570730
rect 216673 570694 219818 570696
rect 139209 570691 139275 570694
rect 216673 570691 216739 570694
rect 201217 570142 201283 570145
rect 200836 570140 201283 570142
rect 120766 570074 120826 570112
rect 200836 570084 201222 570140
rect 201278 570084 201283 570140
rect 200836 570082 201283 570084
rect 201217 570079 201283 570082
rect 123569 570074 123635 570077
rect 120766 570072 123635 570074
rect 120766 570016 123574 570072
rect 123630 570016 123635 570072
rect 120766 570014 123635 570016
rect 280846 570074 280906 570112
rect 281073 570074 281139 570077
rect 280846 570072 281139 570074
rect 280846 570016 281078 570072
rect 281134 570016 281139 570072
rect 280846 570014 281139 570016
rect 123569 570011 123635 570014
rect 281073 570011 281139 570014
rect -960 566796 480 567036
rect 428414 566269 428474 566780
rect 428365 566264 428474 566269
rect 428365 566208 428370 566264
rect 428426 566208 428474 566264
rect 428365 566206 428474 566208
rect 428365 566203 428431 566206
rect 317965 566130 318031 566133
rect 317965 566128 320068 566130
rect 317965 566072 317970 566128
rect 318026 566072 320068 566128
rect 317965 566070 320068 566072
rect 317965 566067 318031 566070
rect 583520 564212 584960 564452
rect 431033 562050 431099 562053
rect 428812 562048 431099 562050
rect 428812 561992 431038 562048
rect 431094 561992 431099 562048
rect 428812 561990 431099 561992
rect 431033 561987 431099 561990
rect 317965 561370 318031 561373
rect 317965 561368 320068 561370
rect 317965 561312 317970 561368
rect 318026 561312 320068 561368
rect 317965 561310 320068 561312
rect 317965 561307 318031 561310
rect 429653 557290 429719 557293
rect 428812 557288 429719 557290
rect 428812 557232 429658 557288
rect 429714 557232 429719 557288
rect 428812 557230 429719 557232
rect 429653 557227 429719 557230
rect 317413 556610 317479 556613
rect 317413 556608 320068 556610
rect 317413 556552 317418 556608
rect 317474 556552 320068 556608
rect 317413 556550 320068 556552
rect 317413 556547 317479 556550
rect -960 553740 480 553980
rect 431125 552530 431191 552533
rect 428812 552528 431191 552530
rect 428812 552472 431130 552528
rect 431186 552472 431191 552528
rect 428812 552470 431191 552472
rect 431125 552467 431191 552470
rect 318057 551850 318123 551853
rect 318057 551848 320068 551850
rect 318057 551792 318062 551848
rect 318118 551792 320068 551848
rect 318057 551790 320068 551792
rect 318057 551787 318123 551790
rect 583520 551020 584960 551260
rect 241513 550082 241579 550085
rect 300301 550082 300367 550085
rect 241513 550080 300367 550082
rect 241513 550024 241518 550080
rect 241574 550024 300306 550080
rect 300362 550024 300367 550080
rect 241513 550022 300367 550024
rect 241513 550019 241579 550022
rect 300301 550019 300367 550022
rect 248689 549946 248755 549949
rect 318057 549946 318123 549949
rect 248689 549944 318123 549946
rect 248689 549888 248694 549944
rect 248750 549888 318062 549944
rect 318118 549888 318123 549944
rect 248689 549886 318123 549888
rect 248689 549883 248755 549886
rect 318057 549883 318123 549886
rect 258717 549810 258783 549813
rect 303061 549810 303127 549813
rect 258717 549808 303127 549810
rect 258717 549752 258722 549808
rect 258778 549752 303066 549808
rect 303122 549752 303127 549808
rect 258717 549750 303127 549752
rect 258717 549747 258783 549750
rect 303061 549747 303127 549750
rect 255129 549674 255195 549677
rect 300577 549674 300643 549677
rect 255129 549672 300643 549674
rect 255129 549616 255134 549672
rect 255190 549616 300582 549672
rect 300638 549616 300643 549672
rect 255129 549614 300643 549616
rect 255129 549611 255195 549614
rect 300577 549611 300643 549614
rect 290917 549538 290983 549541
rect 301497 549538 301563 549541
rect 290917 549536 301563 549538
rect 290917 549480 290922 549536
rect 290978 549480 301502 549536
rect 301558 549480 301563 549536
rect 290917 549478 301563 549480
rect 290917 549475 290983 549478
rect 301497 549475 301563 549478
rect 286685 549402 286751 549405
rect 304349 549402 304415 549405
rect 286685 549400 304415 549402
rect 286685 549344 286690 549400
rect 286746 549344 304354 549400
rect 304410 549344 304415 549400
rect 286685 549342 304415 549344
rect 286685 549339 286751 549342
rect 304349 549339 304415 549342
rect 294505 548178 294571 548181
rect 294505 548176 296730 548178
rect 294505 548120 294510 548176
rect 294566 548120 296730 548176
rect 294505 548118 296730 548120
rect 294505 548115 294571 548118
rect 296670 548042 296730 548118
rect 315573 548042 315639 548045
rect 296670 548040 315639 548042
rect 296670 547984 315578 548040
rect 315634 547984 315639 548040
rect 296670 547982 315639 547984
rect 315573 547979 315639 547982
rect 3417 547906 3483 547909
rect 301589 547906 301655 547909
rect 3417 547904 301655 547906
rect 3417 547848 3422 547904
rect 3478 547848 301594 547904
rect 301650 547848 301655 547904
rect 3417 547846 301655 547848
rect 3417 547843 3483 547846
rect 301589 547843 301655 547846
rect 431217 547770 431283 547773
rect 428812 547768 431283 547770
rect 428812 547712 431222 547768
rect 431278 547712 431283 547768
rect 428812 547710 431283 547712
rect 431217 547707 431283 547710
rect 317965 547090 318031 547093
rect 317965 547088 320068 547090
rect 317965 547032 317970 547088
rect 318026 547032 320068 547088
rect 317965 547030 320068 547032
rect 317965 547027 318031 547030
rect 431309 543010 431375 543013
rect 428812 543008 431375 543010
rect 428812 542952 431314 543008
rect 431370 542952 431375 543008
rect 428812 542950 431375 542952
rect 431309 542947 431375 542950
rect 317965 542330 318031 542333
rect 317965 542328 320068 542330
rect 317965 542272 317970 542328
rect 318026 542272 320068 542328
rect 317965 542270 320068 542272
rect 317965 542267 318031 542270
rect -960 540684 480 540924
rect 302785 540426 302851 540429
rect 299828 540424 302851 540426
rect 299828 540368 302790 540424
rect 302846 540368 302851 540424
rect 299828 540366 302851 540368
rect 302785 540363 302851 540366
rect 429377 538250 429443 538253
rect 428812 538248 429443 538250
rect 428812 538192 429382 538248
rect 429438 538192 429443 538248
rect 428812 538190 429443 538192
rect 429377 538187 429443 538190
rect 583520 537692 584960 537932
rect 318701 537570 318767 537573
rect 318701 537568 320068 537570
rect 318701 537512 318706 537568
rect 318762 537512 320068 537568
rect 318701 537510 320068 537512
rect 318701 537507 318767 537510
rect 431401 533490 431467 533493
rect 428812 533488 431467 533490
rect 428812 533432 431406 533488
rect 431462 533432 431467 533488
rect 428812 533430 431467 533432
rect 431401 533427 431467 533430
rect 318609 532810 318675 532813
rect 318609 532808 320068 532810
rect 318609 532752 318614 532808
rect 318670 532752 320068 532808
rect 318609 532750 320068 532752
rect 318609 532747 318675 532750
rect 427813 528594 427879 528597
rect 428230 528594 428290 528700
rect 427813 528592 428290 528594
rect 427813 528536 427818 528592
rect 427874 528536 428290 528592
rect 427813 528534 428290 528536
rect 427813 528531 427879 528534
rect -960 527764 480 528004
rect 300301 527098 300367 527101
rect 430798 527098 430804 527100
rect 300301 527096 430804 527098
rect 300301 527040 300306 527096
rect 300362 527040 430804 527096
rect 300301 527038 430804 527040
rect 300301 527035 300367 527038
rect 430798 527036 430804 527038
rect 430868 527036 430874 527100
rect 303061 526962 303127 526965
rect 430614 526962 430620 526964
rect 303061 526960 430620 526962
rect 303061 526904 303066 526960
rect 303122 526904 430620 526960
rect 303061 526902 430620 526904
rect 303061 526899 303127 526902
rect 430614 526900 430620 526902
rect 430684 526900 430690 526964
rect 302325 525466 302391 525469
rect 299828 525464 302391 525466
rect 299828 525408 302330 525464
rect 302386 525408 302391 525464
rect 299828 525406 302391 525408
rect 302325 525403 302391 525406
rect 583520 524364 584960 524604
rect 368238 518060 368244 518124
rect 368308 518122 368314 518124
rect 506606 518122 506612 518124
rect 368308 518062 506612 518122
rect 368308 518060 368314 518062
rect 506606 518060 506612 518062
rect 506676 518060 506682 518124
rect 57881 517986 57947 517989
rect 57881 517984 60076 517986
rect 57881 517928 57886 517984
rect 57942 517928 60076 517984
rect 57881 517926 60076 517928
rect 57881 517923 57947 517926
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 302233 510506 302299 510509
rect 299828 510504 302299 510506
rect 299828 510448 302238 510504
rect 302294 510448 302299 510504
rect 299828 510446 302299 510448
rect 302233 510443 302299 510446
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 302233 495546 302299 495549
rect 299828 495544 302299 495546
rect 299828 495488 302238 495544
rect 302294 495488 302299 495544
rect 299828 495486 302299 495488
rect 302233 495483 302299 495486
rect 360878 489092 360884 489156
rect 360948 489154 360954 489156
rect 391933 489154 391999 489157
rect 360948 489152 391999 489154
rect 360948 489096 391938 489152
rect 391994 489096 391999 489152
rect 360948 489094 391999 489096
rect 360948 489092 360954 489094
rect 391933 489091 391999 489094
rect -960 488596 480 488836
rect 364926 487732 364932 487796
rect 364996 487794 365002 487796
rect 506473 487794 506539 487797
rect 364996 487792 506539 487794
rect 364996 487736 506478 487792
rect 506534 487736 506539 487792
rect 364996 487734 506539 487736
rect 364996 487732 365002 487734
rect 506473 487731 506539 487734
rect 363454 486372 363460 486436
rect 363524 486434 363530 486436
rect 488574 486434 488580 486436
rect 363524 486374 488580 486434
rect 363524 486372 363530 486374
rect 488574 486372 488580 486374
rect 488644 486372 488650 486436
rect 68461 485754 68527 485757
rect 77293 485754 77359 485757
rect 68461 485752 77359 485754
rect 68461 485696 68466 485752
rect 68522 485696 77298 485752
rect 77354 485696 77359 485752
rect 68461 485694 77359 485696
rect 68461 485691 68527 485694
rect 77293 485691 77359 485694
rect 187049 485754 187115 485757
rect 199326 485754 199332 485756
rect 187049 485752 199332 485754
rect 187049 485696 187054 485752
rect 187110 485696 199332 485752
rect 187049 485694 199332 485696
rect 187049 485691 187115 485694
rect 199326 485692 199332 485694
rect 199396 485692 199402 485756
rect 233601 485754 233667 485757
rect 366214 485754 366220 485756
rect 233601 485752 366220 485754
rect 233601 485696 233606 485752
rect 233662 485696 366220 485752
rect 233601 485694 366220 485696
rect 233601 485691 233667 485694
rect 366214 485692 366220 485694
rect 366284 485692 366290 485756
rect 55070 485556 55076 485620
rect 55140 485618 55146 485620
rect 73797 485618 73863 485621
rect 55140 485616 73863 485618
rect 55140 485560 73802 485616
rect 73858 485560 73863 485616
rect 55140 485558 73863 485560
rect 55140 485556 55146 485558
rect 73797 485555 73863 485558
rect 171133 485618 171199 485621
rect 198222 485618 198228 485620
rect 171133 485616 198228 485618
rect 171133 485560 171138 485616
rect 171194 485560 198228 485616
rect 171133 485558 198228 485560
rect 171133 485555 171199 485558
rect 198222 485556 198228 485558
rect 198292 485556 198298 485620
rect 205633 485618 205699 485621
rect 206870 485618 206876 485620
rect 205633 485616 206876 485618
rect 205633 485560 205638 485616
rect 205694 485560 206876 485616
rect 205633 485558 206876 485560
rect 205633 485555 205699 485558
rect 206870 485556 206876 485558
rect 206940 485556 206946 485620
rect 208393 485618 208459 485621
rect 209630 485618 209636 485620
rect 208393 485616 209636 485618
rect 208393 485560 208398 485616
rect 208454 485560 209636 485616
rect 208393 485558 209636 485560
rect 208393 485555 208459 485558
rect 209630 485556 209636 485558
rect 209700 485556 209706 485620
rect 235809 485618 235875 485621
rect 371918 485618 371924 485620
rect 235809 485616 371924 485618
rect 235809 485560 235814 485616
rect 235870 485560 371924 485616
rect 235809 485558 371924 485560
rect 235809 485555 235875 485558
rect 371918 485556 371924 485558
rect 371988 485556 371994 485620
rect 54886 485420 54892 485484
rect 54956 485482 54962 485484
rect 76005 485482 76071 485485
rect 54956 485480 76071 485482
rect 54956 485424 76010 485480
rect 76066 485424 76071 485480
rect 54956 485422 76071 485424
rect 54956 485420 54962 485422
rect 76005 485419 76071 485422
rect 148225 485482 148291 485485
rect 198038 485482 198044 485484
rect 148225 485480 198044 485482
rect 148225 485424 148230 485480
rect 148286 485424 198044 485480
rect 148225 485422 198044 485424
rect 148225 485419 148291 485422
rect 198038 485420 198044 485422
rect 198108 485420 198114 485484
rect 232313 485482 232379 485485
rect 371734 485482 371740 485484
rect 232313 485480 371740 485482
rect 232313 485424 232318 485480
rect 232374 485424 371740 485480
rect 232313 485422 371740 485424
rect 232313 485419 232379 485422
rect 371734 485420 371740 485422
rect 371804 485420 371810 485484
rect 44950 485284 44956 485348
rect 45020 485346 45026 485348
rect 66345 485346 66411 485349
rect 45020 485344 66411 485346
rect 45020 485288 66350 485344
rect 66406 485288 66411 485344
rect 45020 485286 66411 485288
rect 45020 485284 45026 485286
rect 66345 485283 66411 485286
rect 73889 485346 73955 485349
rect 95325 485346 95391 485349
rect 73889 485344 95391 485346
rect 73889 485288 73894 485344
rect 73950 485288 95330 485344
rect 95386 485288 95391 485344
rect 73889 485286 95391 485288
rect 73889 485283 73955 485286
rect 95325 485283 95391 485286
rect 145649 485346 145715 485349
rect 197854 485346 197860 485348
rect 145649 485344 197860 485346
rect 145649 485288 145654 485344
rect 145710 485288 197860 485344
rect 145649 485286 197860 485288
rect 145649 485283 145715 485286
rect 197854 485284 197860 485286
rect 197924 485284 197930 485348
rect 199142 485284 199148 485348
rect 199212 485346 199218 485348
rect 218697 485346 218763 485349
rect 199212 485344 218763 485346
rect 199212 485288 218702 485344
rect 218758 485288 218763 485344
rect 199212 485286 218763 485288
rect 199212 485284 199218 485286
rect 218697 485283 218763 485286
rect 231761 485346 231827 485349
rect 370446 485346 370452 485348
rect 231761 485344 370452 485346
rect 231761 485288 231766 485344
rect 231822 485288 370452 485344
rect 231761 485286 370452 485288
rect 231761 485283 231827 485286
rect 370446 485284 370452 485286
rect 370516 485284 370522 485348
rect 57830 485148 57836 485212
rect 57900 485210 57906 485212
rect 91369 485210 91435 485213
rect 57900 485208 91435 485210
rect 57900 485152 91374 485208
rect 91430 485152 91435 485208
rect 57900 485150 91435 485152
rect 57900 485148 57906 485150
rect 91369 485147 91435 485150
rect 147581 485210 147647 485213
rect 200614 485210 200620 485212
rect 147581 485208 200620 485210
rect 147581 485152 147586 485208
rect 147642 485152 200620 485208
rect 147581 485150 200620 485152
rect 147581 485147 147647 485150
rect 200614 485148 200620 485150
rect 200684 485148 200690 485212
rect 205633 485210 205699 485213
rect 206318 485210 206324 485212
rect 205633 485208 206324 485210
rect 205633 485152 205638 485208
rect 205694 485152 206324 485208
rect 205633 485150 206324 485152
rect 205633 485147 205699 485150
rect 206318 485148 206324 485150
rect 206388 485148 206394 485212
rect 219198 485148 219204 485212
rect 219268 485210 219274 485212
rect 226149 485210 226215 485213
rect 219268 485208 226215 485210
rect 219268 485152 226154 485208
rect 226210 485152 226215 485208
rect 219268 485150 226215 485152
rect 219268 485148 219274 485150
rect 226149 485147 226215 485150
rect 234337 485210 234403 485213
rect 373758 485210 373764 485212
rect 234337 485208 373764 485210
rect 234337 485152 234342 485208
rect 234398 485152 373764 485208
rect 234337 485150 373764 485152
rect 234337 485147 234403 485150
rect 373758 485148 373764 485150
rect 373828 485148 373834 485212
rect 375966 485148 375972 485212
rect 376036 485210 376042 485212
rect 511993 485210 512059 485213
rect 376036 485208 512059 485210
rect 376036 485152 511998 485208
rect 512054 485152 512059 485208
rect 376036 485150 512059 485152
rect 376036 485148 376042 485150
rect 511993 485147 512059 485150
rect 53465 485074 53531 485077
rect 94037 485074 94103 485077
rect 53465 485072 94103 485074
rect 53465 485016 53470 485072
rect 53526 485016 94042 485072
rect 94098 485016 94103 485072
rect 53465 485014 94103 485016
rect 53465 485011 53531 485014
rect 94037 485011 94103 485014
rect 145465 485074 145531 485077
rect 202270 485074 202276 485076
rect 145465 485072 202276 485074
rect 145465 485016 145470 485072
rect 145526 485016 202276 485072
rect 145465 485014 202276 485016
rect 145465 485011 145531 485014
rect 202270 485012 202276 485014
rect 202340 485012 202346 485076
rect 203609 485074 203675 485077
rect 217542 485074 217548 485076
rect 203609 485072 217548 485074
rect 203609 485016 203614 485072
rect 203670 485016 217548 485072
rect 203609 485014 217548 485016
rect 203609 485011 203675 485014
rect 217542 485012 217548 485014
rect 217612 485012 217618 485076
rect 223481 485074 223547 485077
rect 376150 485074 376156 485076
rect 223481 485072 376156 485074
rect 223481 485016 223486 485072
rect 223542 485016 376156 485072
rect 223481 485014 376156 485016
rect 223481 485011 223547 485014
rect 376150 485012 376156 485014
rect 376220 485012 376226 485076
rect 59118 484876 59124 484940
rect 59188 484938 59194 484940
rect 68921 484938 68987 484941
rect 59188 484936 68987 484938
rect 59188 484880 68926 484936
rect 68982 484880 68987 484936
rect 59188 484878 68987 484880
rect 59188 484876 59194 484878
rect 68921 484875 68987 484878
rect 185761 484938 185827 484941
rect 196566 484938 196572 484940
rect 185761 484936 196572 484938
rect 185761 484880 185766 484936
rect 185822 484880 196572 484936
rect 185761 484878 196572 484880
rect 185761 484875 185827 484878
rect 196566 484876 196572 484878
rect 196636 484876 196642 484940
rect 197445 484938 197511 484941
rect 198406 484938 198412 484940
rect 197445 484936 198412 484938
rect 197445 484880 197450 484936
rect 197506 484880 198412 484936
rect 197445 484878 198412 484880
rect 197445 484875 197511 484878
rect 198406 484876 198412 484878
rect 198476 484876 198482 484940
rect 201493 484938 201559 484941
rect 202454 484938 202460 484940
rect 201493 484936 202460 484938
rect 201493 484880 201498 484936
rect 201554 484880 202460 484936
rect 201493 484878 202460 484880
rect 201493 484875 201559 484878
rect 202454 484876 202460 484878
rect 202524 484876 202530 484940
rect 211153 484938 211219 484941
rect 211654 484938 211660 484940
rect 211153 484936 211660 484938
rect 211153 484880 211158 484936
rect 211214 484880 211660 484936
rect 211153 484878 211660 484880
rect 211153 484875 211219 484878
rect 211654 484876 211660 484878
rect 211724 484876 211730 484940
rect 235901 484938 235967 484941
rect 360694 484938 360700 484940
rect 235901 484936 360700 484938
rect 235901 484880 235906 484936
rect 235962 484880 360700 484936
rect 235901 484878 360700 484880
rect 235901 484875 235967 484878
rect 360694 484876 360700 484878
rect 360764 484876 360770 484940
rect 59302 484740 59308 484804
rect 59372 484802 59378 484804
rect 72509 484802 72575 484805
rect 59372 484800 72575 484802
rect 59372 484744 72514 484800
rect 72570 484744 72575 484800
rect 59372 484742 72575 484744
rect 59372 484740 59378 484742
rect 72509 484739 72575 484742
rect 200481 484802 200547 484805
rect 200982 484802 200988 484804
rect 200481 484800 200988 484802
rect 200481 484744 200486 484800
rect 200542 484744 200988 484800
rect 200481 484742 200988 484744
rect 200481 484739 200547 484742
rect 200982 484740 200988 484742
rect 201052 484740 201058 484804
rect 211245 484802 211311 484805
rect 211838 484802 211844 484804
rect 211245 484800 211844 484802
rect 211245 484744 211250 484800
rect 211306 484744 211844 484800
rect 211245 484742 211844 484744
rect 211245 484739 211311 484742
rect 211838 484740 211844 484742
rect 211908 484740 211914 484804
rect 76649 484530 76715 484533
rect 80789 484530 80855 484533
rect 76649 484528 80855 484530
rect 76649 484472 76654 484528
rect 76710 484472 80794 484528
rect 80850 484472 80855 484528
rect 76649 484470 80855 484472
rect 76649 484467 76715 484470
rect 80789 484467 80855 484470
rect 200297 484530 200363 484533
rect 201350 484530 201356 484532
rect 200297 484528 201356 484530
rect 200297 484472 200302 484528
rect 200358 484472 201356 484528
rect 200297 484470 201356 484472
rect 200297 484467 200363 484470
rect 201350 484468 201356 484470
rect 201420 484468 201426 484532
rect 205725 484530 205791 484533
rect 206686 484530 206692 484532
rect 205725 484528 206692 484530
rect 205725 484472 205730 484528
rect 205786 484472 206692 484528
rect 205725 484470 206692 484472
rect 205725 484467 205791 484470
rect 206686 484468 206692 484470
rect 206756 484468 206762 484532
rect 214833 484530 214899 484533
rect 216990 484530 216996 484532
rect 214833 484528 216996 484530
rect 214833 484472 214838 484528
rect 214894 484472 216996 484528
rect 214833 484470 216996 484472
rect 214833 484467 214899 484470
rect 216990 484468 216996 484470
rect 217060 484468 217066 484532
rect 219934 484468 219940 484532
rect 220004 484530 220010 484532
rect 224861 484530 224927 484533
rect 220004 484528 224927 484530
rect 220004 484472 224866 484528
rect 224922 484472 224927 484528
rect 583520 484516 584960 484756
rect 220004 484470 224927 484472
rect 220004 484468 220010 484470
rect 224861 484467 224927 484470
rect 164509 484258 164575 484261
rect 164509 484256 171150 484258
rect 164509 484200 164514 484256
rect 164570 484200 171150 484256
rect 164509 484198 171150 484200
rect 164509 484195 164575 484198
rect 171090 483986 171150 484198
rect 216254 483986 216260 483988
rect 171090 483926 216260 483986
rect 216254 483924 216260 483926
rect 216324 483924 216330 483988
rect 156505 483850 156571 483853
rect 213862 483850 213868 483852
rect 156505 483848 213868 483850
rect 156505 483792 156510 483848
rect 156566 483792 213868 483848
rect 156505 483790 213868 483792
rect 156505 483787 156571 483790
rect 213862 483788 213868 483790
rect 213932 483788 213938 483852
rect 144821 483714 144887 483717
rect 214414 483714 214420 483716
rect 144821 483712 214420 483714
rect 144821 483656 144826 483712
rect 144882 483656 214420 483712
rect 144821 483654 214420 483656
rect 144821 483651 144887 483654
rect 214414 483652 214420 483654
rect 214484 483652 214490 483716
rect 57094 482700 57100 482764
rect 57164 482762 57170 482764
rect 121361 482762 121427 482765
rect 57164 482760 121427 482762
rect 57164 482704 121366 482760
rect 121422 482704 121427 482760
rect 57164 482702 121427 482704
rect 57164 482700 57170 482702
rect 121361 482699 121427 482702
rect 48129 482626 48195 482629
rect 120073 482626 120139 482629
rect 48129 482624 120139 482626
rect 48129 482568 48134 482624
rect 48190 482568 120078 482624
rect 120134 482568 120139 482624
rect 48129 482566 120139 482568
rect 48129 482563 48195 482566
rect 120073 482563 120139 482566
rect 277117 482626 277183 482629
rect 359774 482626 359780 482628
rect 277117 482624 359780 482626
rect 277117 482568 277122 482624
rect 277178 482568 359780 482624
rect 277117 482566 359780 482568
rect 277117 482563 277183 482566
rect 359774 482564 359780 482566
rect 359844 482564 359850 482628
rect 48037 482490 48103 482493
rect 120441 482490 120507 482493
rect 48037 482488 120507 482490
rect 48037 482432 48042 482488
rect 48098 482432 120446 482488
rect 120502 482432 120507 482488
rect 48037 482430 120507 482432
rect 48037 482427 48103 482430
rect 120441 482427 120507 482430
rect 154481 482490 154547 482493
rect 212574 482490 212580 482492
rect 154481 482488 212580 482490
rect 154481 482432 154486 482488
rect 154542 482432 212580 482488
rect 154481 482430 212580 482432
rect 154481 482427 154547 482430
rect 212574 482428 212580 482430
rect 212644 482428 212650 482492
rect 236361 482490 236427 482493
rect 375414 482490 375420 482492
rect 236361 482488 375420 482490
rect 236361 482432 236366 482488
rect 236422 482432 375420 482488
rect 236361 482430 375420 482432
rect 236361 482427 236427 482430
rect 375414 482428 375420 482430
rect 375484 482428 375490 482492
rect 46606 482292 46612 482356
rect 46676 482354 46682 482356
rect 124397 482354 124463 482357
rect 46676 482352 124463 482354
rect 46676 482296 124402 482352
rect 124458 482296 124463 482352
rect 46676 482294 124463 482296
rect 46676 482292 46682 482294
rect 124397 482291 124463 482294
rect 148041 482354 148107 482357
rect 215886 482354 215892 482356
rect 148041 482352 215892 482354
rect 148041 482296 148046 482352
rect 148102 482296 215892 482352
rect 148041 482294 215892 482296
rect 148041 482291 148107 482294
rect 215886 482292 215892 482294
rect 215956 482292 215962 482356
rect 222561 482354 222627 482357
rect 374678 482354 374684 482356
rect 222561 482352 374684 482354
rect 222561 482296 222566 482352
rect 222622 482296 374684 482352
rect 222561 482294 374684 482296
rect 222561 482291 222627 482294
rect 374678 482292 374684 482294
rect 374748 482292 374754 482356
rect 3509 482218 3575 482221
rect 312537 482218 312603 482221
rect 3509 482216 312603 482218
rect 3509 482160 3514 482216
rect 3570 482160 312542 482216
rect 312598 482160 312603 482216
rect 3509 482158 312603 482160
rect 3509 482155 3575 482158
rect 312537 482155 312603 482158
rect 280705 481130 280771 481133
rect 377254 481130 377260 481132
rect 280705 481128 377260 481130
rect 280705 481072 280710 481128
rect 280766 481072 377260 481128
rect 280705 481070 377260 481072
rect 280705 481067 280771 481070
rect 377254 481068 377260 481070
rect 377324 481068 377330 481132
rect 179321 480994 179387 480997
rect 217174 480994 217180 480996
rect 179321 480992 217180 480994
rect 179321 480936 179326 480992
rect 179382 480936 217180 480992
rect 179321 480934 217180 480936
rect 179321 480931 179387 480934
rect 217174 480932 217180 480934
rect 217244 480932 217250 480996
rect 247309 480994 247375 480997
rect 374862 480994 374868 480996
rect 247309 480992 374868 480994
rect 247309 480936 247314 480992
rect 247370 480936 374868 480992
rect 247309 480934 374868 480936
rect 247309 480931 247375 480934
rect 374862 480932 374868 480934
rect 374932 480932 374938 480996
rect 147213 480858 147279 480861
rect 203190 480858 203196 480860
rect 147213 480856 203196 480858
rect 147213 480800 147218 480856
rect 147274 480800 203196 480856
rect 147213 480798 203196 480800
rect 147213 480795 147279 480798
rect 203190 480796 203196 480798
rect 203260 480796 203266 480860
rect 233969 480858 234035 480861
rect 378726 480858 378732 480860
rect 233969 480856 378732 480858
rect 233969 480800 233974 480856
rect 234030 480800 378732 480856
rect 233969 480798 378732 480800
rect 233969 480795 234035 480798
rect 378726 480796 378732 480798
rect 378796 480796 378802 480860
rect 59077 479906 59143 479909
rect 95509 479906 95575 479909
rect 59077 479904 95575 479906
rect 59077 479848 59082 479904
rect 59138 479848 95514 479904
rect 95570 479848 95575 479904
rect 59077 479846 95575 479848
rect 59077 479843 59143 479846
rect 95509 479843 95575 479846
rect 57462 479708 57468 479772
rect 57532 479770 57538 479772
rect 118785 479770 118851 479773
rect 57532 479768 118851 479770
rect 57532 479712 118790 479768
rect 118846 479712 118851 479768
rect 57532 479710 118851 479712
rect 57532 479708 57538 479710
rect 118785 479707 118851 479710
rect 172053 479770 172119 479773
rect 213126 479770 213132 479772
rect 172053 479768 213132 479770
rect 172053 479712 172058 479768
rect 172114 479712 213132 479768
rect 172053 479710 213132 479712
rect 172053 479707 172119 479710
rect 213126 479708 213132 479710
rect 213196 479708 213202 479772
rect 256325 479770 256391 479773
rect 359406 479770 359412 479772
rect 256325 479768 359412 479770
rect 256325 479712 256330 479768
rect 256386 479712 359412 479768
rect 256325 479710 359412 479712
rect 256325 479707 256391 479710
rect 359406 479708 359412 479710
rect 359476 479708 359482 479772
rect 59813 479634 59879 479637
rect 124489 479634 124555 479637
rect 59813 479632 124555 479634
rect 59813 479576 59818 479632
rect 59874 479576 124494 479632
rect 124550 479576 124555 479632
rect 59813 479574 124555 479576
rect 59813 479571 59879 479574
rect 124489 479571 124555 479574
rect 154665 479634 154731 479637
rect 215334 479634 215340 479636
rect 154665 479632 215340 479634
rect 154665 479576 154670 479632
rect 154726 479576 215340 479632
rect 154665 479574 215340 479576
rect 154665 479571 154731 479574
rect 215334 479572 215340 479574
rect 215404 479572 215410 479636
rect 229829 479634 229895 479637
rect 374494 479634 374500 479636
rect 229829 479632 374500 479634
rect 229829 479576 229834 479632
rect 229890 479576 374500 479632
rect 229829 479574 374500 479576
rect 229829 479571 229895 479574
rect 374494 479572 374500 479574
rect 374564 479572 374570 479636
rect 50521 479498 50587 479501
rect 121913 479498 121979 479501
rect 50521 479496 121979 479498
rect 50521 479440 50526 479496
rect 50582 479440 121918 479496
rect 121974 479440 121979 479496
rect 50521 479438 121979 479440
rect 50521 479435 50587 479438
rect 121913 479435 121979 479438
rect 148317 479498 148383 479501
rect 208894 479498 208900 479500
rect 148317 479496 208900 479498
rect 148317 479440 148322 479496
rect 148378 479440 208900 479496
rect 148317 479438 208900 479440
rect 148317 479435 148383 479438
rect 208894 479436 208900 479438
rect 208964 479436 208970 479500
rect 210366 479436 210372 479500
rect 210436 479498 210442 479500
rect 512085 479498 512151 479501
rect 210436 479496 512151 479498
rect 210436 479440 512090 479496
rect 512146 479440 512151 479496
rect 210436 479438 512151 479440
rect 210436 479436 210442 479438
rect 512085 479435 512151 479438
rect 297173 478546 297239 478549
rect 377438 478546 377444 478548
rect 297173 478544 377444 478546
rect 297173 478488 297178 478544
rect 297234 478488 377444 478544
rect 297173 478486 377444 478488
rect 297173 478483 297239 478486
rect 377438 478484 377444 478486
rect 377508 478484 377514 478548
rect 145741 478410 145807 478413
rect 205030 478410 205036 478412
rect 145741 478408 205036 478410
rect 145741 478352 145746 478408
rect 145802 478352 205036 478408
rect 145741 478350 205036 478352
rect 145741 478347 145807 478350
rect 205030 478348 205036 478350
rect 205100 478348 205106 478412
rect 234613 478410 234679 478413
rect 357566 478410 357572 478412
rect 234613 478408 357572 478410
rect 234613 478352 234618 478408
rect 234674 478352 357572 478408
rect 234613 478350 357572 478352
rect 234613 478347 234679 478350
rect 357566 478348 357572 478350
rect 357636 478348 357642 478412
rect 151353 478274 151419 478277
rect 214598 478274 214604 478276
rect 151353 478272 214604 478274
rect 151353 478216 151358 478272
rect 151414 478216 214604 478272
rect 151353 478214 214604 478216
rect 151353 478211 151419 478214
rect 214598 478212 214604 478214
rect 214668 478212 214674 478276
rect 223573 478274 223639 478277
rect 378910 478274 378916 478276
rect 223573 478272 378916 478274
rect 223573 478216 223578 478272
rect 223634 478216 378916 478272
rect 223573 478214 378916 478216
rect 223573 478211 223639 478214
rect 378910 478212 378916 478214
rect 378980 478212 378986 478276
rect 204846 478076 204852 478140
rect 204916 478138 204922 478140
rect 457529 478138 457595 478141
rect 204916 478136 457595 478138
rect 204916 478080 457534 478136
rect 457590 478080 457595 478136
rect 204916 478078 457595 478080
rect 204916 478076 204922 478078
rect 457529 478075 457595 478078
rect 46790 476852 46796 476916
rect 46860 476914 46866 476916
rect 123661 476914 123727 476917
rect 46860 476912 123727 476914
rect 46860 476856 123666 476912
rect 123722 476856 123727 476912
rect 46860 476854 123727 476856
rect 46860 476852 46866 476854
rect 123661 476851 123727 476854
rect 163773 476914 163839 476917
rect 213310 476914 213316 476916
rect 163773 476912 213316 476914
rect 163773 476856 163778 476912
rect 163834 476856 213316 476912
rect 163773 476854 213316 476856
rect 163773 476851 163839 476854
rect 213310 476852 213316 476854
rect 213380 476852 213386 476916
rect 227989 476914 228055 476917
rect 357934 476914 357940 476916
rect 227989 476912 357940 476914
rect 227989 476856 227994 476912
rect 228050 476856 357940 476912
rect 227989 476854 357940 476856
rect 227989 476851 228055 476854
rect 357934 476852 357940 476854
rect 358004 476852 358010 476916
rect 44766 476716 44772 476780
rect 44836 476778 44842 476780
rect 126329 476778 126395 476781
rect 44836 476776 126395 476778
rect 44836 476720 126334 476776
rect 126390 476720 126395 476776
rect 44836 476718 126395 476720
rect 44836 476716 44842 476718
rect 126329 476715 126395 476718
rect 157517 476778 157583 476781
rect 209814 476778 209820 476780
rect 157517 476776 209820 476778
rect 157517 476720 157522 476776
rect 157578 476720 209820 476776
rect 157517 476718 209820 476720
rect 157517 476715 157583 476718
rect 209814 476716 209820 476718
rect 209884 476716 209890 476780
rect 230749 476778 230815 476781
rect 379094 476778 379100 476780
rect 230749 476776 379100 476778
rect 230749 476720 230754 476776
rect 230810 476720 379100 476776
rect 230749 476718 379100 476720
rect 230749 476715 230815 476718
rect 379094 476716 379100 476718
rect 379164 476716 379170 476780
rect 254117 475962 254183 475965
rect 376886 475962 376892 475964
rect 254117 475960 376892 475962
rect 254117 475904 254122 475960
rect 254178 475904 376892 475960
rect 254117 475902 376892 475904
rect 254117 475899 254183 475902
rect 376886 475900 376892 475902
rect 376956 475900 376962 475964
rect 231945 475826 232011 475829
rect 367686 475826 367692 475828
rect 231945 475824 367692 475826
rect -960 475540 480 475780
rect 231945 475768 231950 475824
rect 232006 475768 367692 475824
rect 231945 475766 367692 475768
rect 231945 475763 232011 475766
rect 367686 475764 367692 475766
rect 367756 475764 367762 475828
rect 161657 475690 161723 475693
rect 207974 475690 207980 475692
rect 161657 475688 207980 475690
rect 161657 475632 161662 475688
rect 161718 475632 207980 475688
rect 161657 475630 207980 475632
rect 161657 475627 161723 475630
rect 207974 475628 207980 475630
rect 208044 475628 208050 475692
rect 240317 475690 240383 475693
rect 379462 475690 379468 475692
rect 240317 475688 379468 475690
rect 240317 475632 240322 475688
rect 240378 475632 379468 475688
rect 240317 475630 379468 475632
rect 240317 475627 240383 475630
rect 379462 475628 379468 475630
rect 379532 475628 379538 475692
rect 156781 475554 156847 475557
rect 218646 475554 218652 475556
rect 156781 475552 218652 475554
rect 156781 475496 156786 475552
rect 156842 475496 218652 475552
rect 156781 475494 218652 475496
rect 156781 475491 156847 475494
rect 218646 475492 218652 475494
rect 218716 475492 218722 475556
rect 226517 475554 226583 475557
rect 379278 475554 379284 475556
rect 226517 475552 379284 475554
rect 226517 475496 226522 475552
rect 226578 475496 379284 475552
rect 226517 475494 379284 475496
rect 226517 475491 226583 475494
rect 379278 475492 379284 475494
rect 379348 475492 379354 475556
rect 202086 475356 202092 475420
rect 202156 475418 202162 475420
rect 483013 475418 483079 475421
rect 202156 475416 483079 475418
rect 202156 475360 483018 475416
rect 483074 475360 483079 475416
rect 202156 475358 483079 475360
rect 202156 475356 202162 475358
rect 483013 475355 483079 475358
rect 153193 474330 153259 474333
rect 218830 474330 218836 474332
rect 153193 474328 218836 474330
rect 153193 474272 153198 474328
rect 153254 474272 218836 474328
rect 153193 474270 218836 474272
rect 153193 474267 153259 474270
rect 218830 474268 218836 474270
rect 218900 474268 218906 474332
rect 127341 474194 127407 474197
rect 196750 474194 196756 474196
rect 127341 474192 196756 474194
rect 127341 474136 127346 474192
rect 127402 474136 196756 474192
rect 127341 474134 196756 474136
rect 127341 474131 127407 474134
rect 196750 474132 196756 474134
rect 196820 474132 196826 474196
rect 143533 474058 143599 474061
rect 216070 474058 216076 474060
rect 143533 474056 216076 474058
rect 143533 474000 143538 474056
rect 143594 474000 216076 474056
rect 143533 473998 216076 474000
rect 143533 473995 143599 473998
rect 216070 473996 216076 473998
rect 216140 473996 216146 474060
rect 171225 472698 171291 472701
rect 203006 472698 203012 472700
rect 171225 472696 203012 472698
rect 171225 472640 171230 472696
rect 171286 472640 203012 472696
rect 171225 472638 203012 472640
rect 171225 472635 171291 472638
rect 203006 472636 203012 472638
rect 203076 472636 203082 472700
rect 152733 472562 152799 472565
rect 204294 472562 204300 472564
rect 152733 472560 204300 472562
rect 152733 472504 152738 472560
rect 152794 472504 204300 472560
rect 152733 472502 204300 472504
rect 152733 472499 152799 472502
rect 204294 472500 204300 472502
rect 204364 472500 204370 472564
rect 365110 472500 365116 472564
rect 365180 472562 365186 472564
rect 476062 472562 476068 472564
rect 365180 472502 476068 472562
rect 365180 472500 365186 472502
rect 476062 472500 476068 472502
rect 476132 472500 476138 472564
rect 182725 471882 182791 471885
rect 199510 471882 199516 471884
rect 182725 471880 199516 471882
rect 182725 471824 182730 471880
rect 182786 471824 199516 471880
rect 182725 471822 199516 471824
rect 182725 471819 182791 471822
rect 199510 471820 199516 471822
rect 199580 471820 199586 471884
rect 59169 471746 59235 471749
rect 91921 471746 91987 471749
rect 59169 471744 91987 471746
rect 59169 471688 59174 471744
rect 59230 471688 91926 471744
rect 91982 471688 91987 471744
rect 59169 471686 91987 471688
rect 59169 471683 59235 471686
rect 91921 471683 91987 471686
rect 183645 471746 183711 471749
rect 217358 471746 217364 471748
rect 183645 471744 217364 471746
rect 183645 471688 183650 471744
rect 183706 471688 217364 471744
rect 183645 471686 217364 471688
rect 183645 471683 183711 471686
rect 217358 471684 217364 471686
rect 217428 471684 217434 471748
rect 55029 471610 55095 471613
rect 88517 471610 88583 471613
rect 55029 471608 88583 471610
rect 55029 471552 55034 471608
rect 55090 471552 88522 471608
rect 88578 471552 88583 471608
rect 55029 471550 88583 471552
rect 55029 471547 55095 471550
rect 88517 471547 88583 471550
rect 172605 471610 172671 471613
rect 211981 471610 212047 471613
rect 172605 471608 212047 471610
rect 172605 471552 172610 471608
rect 172666 471552 211986 471608
rect 212042 471552 212047 471608
rect 172605 471550 212047 471552
rect 172605 471547 172671 471550
rect 211981 471547 212047 471550
rect 54201 471474 54267 471477
rect 88425 471474 88491 471477
rect 54201 471472 88491 471474
rect 54201 471416 54206 471472
rect 54262 471416 88430 471472
rect 88486 471416 88491 471472
rect 54201 471414 88491 471416
rect 54201 471411 54267 471414
rect 88425 471411 88491 471414
rect 162853 471474 162919 471477
rect 203701 471474 203767 471477
rect 162853 471472 203767 471474
rect 162853 471416 162858 471472
rect 162914 471416 203706 471472
rect 203762 471416 203767 471472
rect 162853 471414 203767 471416
rect 162853 471411 162919 471414
rect 203701 471411 203767 471414
rect 56133 471338 56199 471341
rect 89805 471338 89871 471341
rect 56133 471336 89871 471338
rect 56133 471280 56138 471336
rect 56194 471280 89810 471336
rect 89866 471280 89871 471336
rect 56133 471278 89871 471280
rect 56133 471275 56199 471278
rect 89805 471275 89871 471278
rect 161565 471338 161631 471341
rect 203517 471338 203583 471341
rect 161565 471336 203583 471338
rect 161565 471280 161570 471336
rect 161626 471280 203522 471336
rect 203578 471280 203583 471336
rect 583520 471324 584960 471564
rect 161565 471278 203583 471280
rect 161565 471275 161631 471278
rect 203517 471275 203583 471278
rect 53281 471202 53347 471205
rect 87505 471202 87571 471205
rect 53281 471200 87571 471202
rect 53281 471144 53286 471200
rect 53342 471144 87510 471200
rect 87566 471144 87571 471200
rect 53281 471142 87571 471144
rect 53281 471139 53347 471142
rect 87505 471139 87571 471142
rect 161749 471202 161815 471205
rect 214741 471202 214807 471205
rect 161749 471200 214807 471202
rect 161749 471144 161754 471200
rect 161810 471144 214746 471200
rect 214802 471144 214807 471200
rect 161749 471142 214807 471144
rect 161749 471139 161815 471142
rect 214741 471139 214807 471142
rect 298185 471202 298251 471205
rect 377622 471202 377628 471204
rect 298185 471200 377628 471202
rect 298185 471144 298190 471200
rect 298246 471144 377628 471200
rect 298185 471142 377628 471144
rect 298185 471139 298251 471142
rect 377622 471140 377628 471142
rect 377692 471140 377698 471204
rect 169845 469978 169911 469981
rect 206134 469978 206140 469980
rect 169845 469976 206140 469978
rect 169845 469920 169850 469976
rect 169906 469920 206140 469976
rect 169845 469918 206140 469920
rect 169845 469915 169911 469918
rect 206134 469916 206140 469918
rect 206204 469916 206210 469980
rect 58934 469780 58940 469844
rect 59004 469842 59010 469844
rect 67817 469842 67883 469845
rect 59004 469840 67883 469842
rect 59004 469784 67822 469840
rect 67878 469784 67883 469840
rect 59004 469782 67883 469784
rect 59004 469780 59010 469782
rect 67817 469779 67883 469782
rect 160093 469842 160159 469845
rect 200798 469842 200804 469844
rect 160093 469840 200804 469842
rect 160093 469784 160098 469840
rect 160154 469784 200804 469840
rect 160093 469782 200804 469784
rect 160093 469779 160159 469782
rect 200798 469780 200804 469782
rect 200868 469780 200874 469844
rect 47894 469100 47900 469164
rect 47964 469162 47970 469164
rect 69197 469162 69263 469165
rect 47964 469160 69263 469162
rect 47964 469104 69202 469160
rect 69258 469104 69263 469160
rect 47964 469102 69263 469104
rect 47964 469100 47970 469102
rect 69197 469099 69263 469102
rect 48630 468964 48636 469028
rect 48700 469026 48706 469028
rect 70577 469026 70643 469029
rect 48700 469024 70643 469026
rect 48700 468968 70582 469024
rect 70638 468968 70643 469024
rect 48700 468966 70643 468968
rect 48700 468964 48706 468966
rect 70577 468963 70643 468966
rect 169753 469026 169819 469029
rect 202321 469026 202387 469029
rect 169753 469024 202387 469026
rect 169753 468968 169758 469024
rect 169814 468968 202326 469024
rect 202382 468968 202387 469024
rect 169753 468966 202387 468968
rect 169753 468963 169819 468966
rect 202321 468963 202387 468966
rect 55622 468828 55628 468892
rect 55692 468890 55698 468892
rect 78857 468890 78923 468893
rect 55692 468888 78923 468890
rect 55692 468832 78862 468888
rect 78918 468832 78923 468888
rect 55692 468830 78923 468832
rect 55692 468828 55698 468830
rect 78857 468827 78923 468830
rect 167269 468890 167335 468893
rect 206461 468890 206527 468893
rect 167269 468888 206527 468890
rect 167269 468832 167274 468888
rect 167330 468832 206466 468888
rect 206522 468832 206527 468888
rect 167269 468830 206527 468832
rect 167269 468827 167335 468830
rect 206461 468827 206527 468830
rect 53598 468692 53604 468756
rect 53668 468754 53674 468756
rect 78949 468754 79015 468757
rect 53668 468752 79015 468754
rect 53668 468696 78954 468752
rect 79010 468696 79015 468752
rect 53668 468694 79015 468696
rect 53668 468692 53674 468694
rect 78949 468691 79015 468694
rect 168373 468754 168439 468757
rect 209129 468754 209195 468757
rect 168373 468752 209195 468754
rect 168373 468696 168378 468752
rect 168434 468696 209134 468752
rect 209190 468696 209195 468752
rect 168373 468694 209195 468696
rect 168373 468691 168439 468694
rect 209129 468691 209195 468694
rect 50470 468556 50476 468620
rect 50540 468618 50546 468620
rect 77385 468618 77451 468621
rect 50540 468616 77451 468618
rect 50540 468560 77390 468616
rect 77446 468560 77451 468616
rect 50540 468558 77451 468560
rect 50540 468556 50546 468558
rect 77385 468555 77451 468558
rect 167085 468618 167151 468621
rect 210601 468618 210667 468621
rect 167085 468616 210667 468618
rect 167085 468560 167090 468616
rect 167146 468560 210606 468616
rect 210662 468560 210667 468616
rect 167085 468558 210667 468560
rect 167085 468555 167151 468558
rect 210601 468555 210667 468558
rect 50838 468420 50844 468484
rect 50908 468482 50914 468484
rect 78765 468482 78831 468485
rect 50908 468480 78831 468482
rect 50908 468424 78770 468480
rect 78826 468424 78831 468480
rect 50908 468422 78831 468424
rect 50908 468420 50914 468422
rect 78765 468419 78831 468422
rect 168557 468482 168623 468485
rect 213494 468482 213500 468484
rect 168557 468480 213500 468482
rect 168557 468424 168562 468480
rect 168618 468424 213500 468480
rect 168557 468422 213500 468424
rect 168557 468419 168623 468422
rect 213494 468420 213500 468422
rect 213564 468420 213570 468484
rect 265065 468482 265131 468485
rect 359590 468482 359596 468484
rect 265065 468480 359596 468482
rect 265065 468424 265070 468480
rect 265126 468424 359596 468480
rect 265065 468422 359596 468424
rect 265065 468419 265131 468422
rect 359590 468420 359596 468422
rect 359660 468420 359666 468484
rect 58750 468284 58756 468348
rect 58820 468346 58826 468348
rect 67725 468346 67791 468349
rect 58820 468344 67791 468346
rect 58820 468288 67730 468344
rect 67786 468288 67791 468344
rect 58820 468286 67791 468288
rect 58820 468284 58826 468286
rect 67725 468283 67791 468286
rect 48078 467876 48084 467940
rect 48148 467938 48154 467940
rect 48221 467938 48287 467941
rect 50705 467940 50771 467941
rect 50654 467938 50660 467940
rect 48148 467936 48287 467938
rect 48148 467880 48226 467936
rect 48282 467880 48287 467936
rect 48148 467878 48287 467880
rect 50614 467878 50660 467938
rect 50724 467936 50771 467940
rect 50766 467880 50771 467936
rect 48148 467876 48154 467878
rect 48221 467875 48287 467878
rect 50654 467876 50660 467878
rect 50724 467876 50771 467880
rect 50705 467875 50771 467876
rect 154573 467258 154639 467261
rect 208342 467258 208348 467260
rect 154573 467256 208348 467258
rect 154573 467200 154578 467256
rect 154634 467200 208348 467256
rect 154573 467198 208348 467200
rect 154573 467195 154639 467198
rect 208342 467196 208348 467198
rect 208412 467196 208418 467260
rect 60222 467060 60228 467124
rect 60292 467122 60298 467124
rect 73337 467122 73403 467125
rect 60292 467120 73403 467122
rect 60292 467064 73342 467120
rect 73398 467064 73403 467120
rect 60292 467062 73403 467064
rect 60292 467060 60298 467062
rect 73337 467059 73403 467062
rect 151813 467122 151879 467125
rect 209998 467122 210004 467124
rect 151813 467120 210004 467122
rect 151813 467064 151818 467120
rect 151874 467064 210004 467120
rect 151813 467062 210004 467064
rect 151813 467059 151879 467062
rect 209998 467060 210004 467062
rect 210068 467060 210074 467124
rect 179638 466924 179644 466988
rect 179708 466986 179714 466988
rect 180149 466986 180215 466989
rect 179708 466984 180215 466986
rect 179708 466928 180154 466984
rect 180210 466928 180215 466984
rect 179708 466926 180215 466928
rect 179708 466924 179714 466926
rect 180149 466923 180215 466926
rect 178033 466578 178099 466581
rect 190913 466580 190979 466581
rect 338481 466580 338547 466581
rect 339769 466580 339835 466581
rect 350993 466580 351059 466581
rect 178350 466578 178356 466580
rect 178033 466576 178356 466578
rect 178033 466520 178038 466576
rect 178094 466520 178356 466576
rect 178033 466518 178356 466520
rect 178033 466515 178099 466518
rect 178350 466516 178356 466518
rect 178420 466516 178426 466580
rect 190862 466578 190868 466580
rect 190822 466518 190868 466578
rect 190932 466576 190979 466580
rect 338430 466578 338436 466580
rect 190974 466520 190979 466576
rect 190862 466516 190868 466518
rect 190932 466516 190979 466520
rect 338390 466518 338436 466578
rect 338500 466576 338547 466580
rect 339718 466578 339724 466580
rect 338542 466520 338547 466576
rect 338430 466516 338436 466518
rect 338500 466516 338547 466520
rect 339678 466518 339724 466578
rect 339788 466576 339835 466580
rect 350942 466578 350948 466580
rect 339830 466520 339835 466576
rect 339718 466516 339724 466518
rect 339788 466516 339835 466520
rect 350902 466518 350948 466578
rect 351012 466576 351059 466580
rect 351054 466520 351059 466576
rect 350942 466516 350948 466518
rect 351012 466516 351059 466520
rect 190913 466515 190979 466516
rect 338481 466515 338547 466516
rect 339769 466515 339835 466516
rect 350993 466515 351059 466516
rect 498193 466578 498259 466581
rect 499757 466580 499823 466581
rect 510889 466580 510955 466581
rect 498510 466578 498516 466580
rect 498193 466576 498516 466578
rect 498193 466520 498198 466576
rect 498254 466520 498516 466576
rect 498193 466518 498516 466520
rect 498193 466515 498259 466518
rect 498510 466516 498516 466518
rect 498580 466516 498586 466580
rect 499757 466576 499804 466580
rect 499868 466578 499874 466580
rect 510838 466578 510844 466580
rect 499757 466520 499762 466576
rect 499757 466516 499804 466520
rect 499868 466518 499914 466578
rect 510798 466518 510844 466578
rect 510908 466576 510955 466580
rect 510950 466520 510955 466576
rect 499868 466516 499874 466518
rect 510838 466516 510844 466518
rect 510908 466516 510955 466520
rect 499757 466515 499823 466516
rect 510889 466515 510955 466516
rect 54702 466380 54708 466444
rect 54772 466442 54778 466444
rect 71773 466442 71839 466445
rect 54772 466440 71839 466442
rect 54772 466384 71778 466440
rect 71834 466384 71839 466440
rect 54772 466382 71839 466384
rect 54772 466380 54778 466382
rect 71773 466379 71839 466382
rect 57646 466244 57652 466308
rect 57716 466306 57722 466308
rect 76557 466306 76623 466309
rect 57716 466304 76623 466306
rect 57716 466248 76562 466304
rect 76618 466248 76623 466304
rect 57716 466246 76623 466248
rect 57716 466244 57722 466246
rect 76557 466243 76623 466246
rect 48446 466108 48452 466172
rect 48516 466170 48522 466172
rect 48516 466110 55230 466170
rect 48516 466108 48522 466110
rect 53230 465972 53236 466036
rect 53300 466034 53306 466036
rect 53649 466034 53715 466037
rect 53300 466032 53715 466034
rect 53300 465976 53654 466032
rect 53710 465976 53715 466032
rect 53300 465974 53715 465976
rect 55170 466034 55230 466110
rect 55438 466108 55444 466172
rect 55508 466170 55514 466172
rect 74625 466170 74691 466173
rect 55508 466168 74691 466170
rect 55508 466112 74630 466168
rect 74686 466112 74691 466168
rect 55508 466110 74691 466112
rect 55508 466108 55514 466110
rect 74625 466107 74691 466110
rect 180057 466170 180123 466173
rect 198774 466170 198780 466172
rect 180057 466168 198780 466170
rect 180057 466112 180062 466168
rect 180118 466112 198780 466168
rect 180057 466110 198780 466112
rect 180057 466107 180123 466110
rect 198774 466108 198780 466110
rect 198844 466108 198850 466172
rect 70393 466034 70459 466037
rect 55170 466032 70459 466034
rect 55170 465976 70398 466032
rect 70454 465976 70459 466032
rect 55170 465974 70459 465976
rect 53300 465972 53306 465974
rect 53649 465971 53715 465974
rect 70393 465971 70459 465974
rect 166993 466034 167059 466037
rect 203609 466034 203675 466037
rect 166993 466032 203675 466034
rect 166993 465976 166998 466032
rect 167054 465976 203614 466032
rect 203670 465976 203675 466032
rect 166993 465974 203675 465976
rect 166993 465971 167059 465974
rect 203609 465971 203675 465974
rect 52126 465836 52132 465900
rect 52196 465898 52202 465900
rect 74533 465898 74599 465901
rect 52196 465896 74599 465898
rect 52196 465840 74538 465896
rect 74594 465840 74599 465896
rect 52196 465838 74599 465840
rect 52196 465836 52202 465838
rect 74533 465835 74599 465838
rect 165797 465898 165863 465901
rect 205214 465898 205220 465900
rect 165797 465896 205220 465898
rect 165797 465840 165802 465896
rect 165858 465840 205220 465896
rect 165797 465838 205220 465840
rect 165797 465835 165863 465838
rect 205214 465836 205220 465838
rect 205284 465836 205290 465900
rect 52310 465700 52316 465764
rect 52380 465762 52386 465764
rect 76005 465762 76071 465765
rect 52380 465760 76071 465762
rect 52380 465704 76010 465760
rect 76066 465704 76071 465760
rect 52380 465702 76071 465704
rect 52380 465700 52386 465702
rect 76005 465699 76071 465702
rect 165613 465762 165679 465765
rect 218973 465762 219039 465765
rect 165613 465760 219039 465762
rect 165613 465704 165618 465760
rect 165674 465704 218978 465760
rect 219034 465704 219039 465760
rect 165613 465702 219039 465704
rect 165613 465699 165679 465702
rect 218973 465699 219039 465702
rect 292573 465762 292639 465765
rect 359958 465762 359964 465764
rect 292573 465760 359964 465762
rect 292573 465704 292578 465760
rect 292634 465704 359964 465760
rect 292573 465702 359964 465704
rect 292573 465699 292639 465702
rect 359958 465700 359964 465702
rect 360028 465700 360034 465764
rect 58566 465564 58572 465628
rect 58636 465626 58642 465628
rect 69105 465626 69171 465629
rect 58636 465624 69171 465626
rect 58636 465568 69110 465624
rect 69166 465568 69171 465624
rect 58636 465566 69171 465568
rect 58636 465564 58642 465566
rect 69105 465563 69171 465566
rect 51758 465156 51764 465220
rect 51828 465218 51834 465220
rect 52361 465218 52427 465221
rect 51828 465216 52427 465218
rect 51828 465160 52366 465216
rect 52422 465160 52427 465216
rect 51828 465158 52427 465160
rect 51828 465156 51834 465158
rect 52361 465155 52427 465158
rect 171133 464402 171199 464405
rect 208158 464402 208164 464404
rect 171133 464400 208164 464402
rect 171133 464344 171138 464400
rect 171194 464344 208164 464400
rect 171133 464342 208164 464344
rect 171133 464339 171199 464342
rect 208158 464340 208164 464342
rect 208228 464340 208234 464404
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 196558 460186 196618 460190
rect 198917 460186 198983 460189
rect 196558 460184 198983 460186
rect 196558 460128 198922 460184
rect 198978 460128 198983 460184
rect 196558 460126 198983 460128
rect 356562 460186 356622 460190
rect 358813 460186 358879 460189
rect 356562 460184 358879 460186
rect 356562 460128 358818 460184
rect 358874 460128 358879 460184
rect 356562 460126 358879 460128
rect 198917 460123 198983 460126
rect 358813 460123 358879 460126
rect 516558 459642 516618 460190
rect 518893 459642 518959 459645
rect 519537 459642 519603 459645
rect 516558 459640 519603 459642
rect 516558 459584 518898 459640
rect 518954 459584 519542 459640
rect 519598 459584 519603 459640
rect 516558 459582 519603 459584
rect 518893 459579 518959 459582
rect 519537 459579 519603 459582
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 57237 417346 57303 417349
rect 60002 417346 60062 417894
rect 216673 417890 216739 417893
rect 219390 417890 220064 417924
rect 216673 417888 220064 417890
rect 216673 417832 216678 417888
rect 216734 417864 220064 417888
rect 377581 417890 377647 417893
rect 379470 417890 380052 417924
rect 377581 417888 380052 417890
rect 216734 417832 219450 417864
rect 216673 417830 219450 417832
rect 377581 417832 377586 417888
rect 377642 417864 380052 417888
rect 377642 417832 379530 417864
rect 377581 417830 379530 417832
rect 216673 417827 216739 417830
rect 377581 417827 377647 417830
rect 357566 417420 357572 417484
rect 357636 417482 357642 417484
rect 358629 417482 358695 417485
rect 357636 417480 358695 417482
rect 357636 417424 358634 417480
rect 358690 417424 358695 417480
rect 357636 417422 358695 417424
rect 357636 417420 357642 417422
rect 358629 417419 358695 417422
rect 57237 417344 60062 417346
rect 57237 417288 57242 417344
rect 57298 417288 60062 417344
rect 57237 417286 60062 417288
rect 57237 417283 57303 417286
rect 57881 417210 57947 417213
rect 57881 417208 60062 417210
rect 57881 417152 57886 417208
rect 57942 417152 60062 417208
rect 57881 417150 60062 417152
rect 57881 417147 57947 417150
rect 60002 416942 60062 417150
rect 217961 416938 218027 416941
rect 219390 416938 220064 416972
rect 217961 416936 220064 416938
rect 217961 416880 217966 416936
rect 218022 416912 220064 416936
rect 377213 416938 377279 416941
rect 377857 416938 377923 416941
rect 379470 416938 380052 416972
rect 377213 416936 380052 416938
rect 218022 416880 219450 416912
rect 217961 416878 219450 416880
rect 377213 416880 377218 416936
rect 377274 416880 377862 416936
rect 377918 416912 380052 416936
rect 377918 416880 379530 416912
rect 377213 416878 379530 416880
rect 217961 416875 218027 416878
rect 377213 416875 377279 416878
rect 377857 416875 377923 416878
rect 57881 414218 57947 414221
rect 60002 414218 60062 414766
rect 217041 414762 217107 414765
rect 219390 414762 220064 414796
rect 217041 414760 220064 414762
rect 217041 414704 217046 414760
rect 217102 414736 220064 414760
rect 377673 414762 377739 414765
rect 379470 414762 380052 414796
rect 377673 414760 380052 414762
rect 217102 414704 219450 414736
rect 217041 414702 219450 414704
rect 377673 414704 377678 414760
rect 377734 414736 380052 414760
rect 377734 414704 379530 414736
rect 377673 414702 379530 414704
rect 217041 414699 217107 414702
rect 377673 414699 377739 414702
rect 57881 414216 60062 414218
rect 57881 414160 57886 414216
rect 57942 414160 60062 414216
rect 57881 414158 60062 414160
rect 57881 414155 57947 414158
rect 204294 413884 204300 413948
rect 204364 413946 204370 413948
rect 205541 413946 205607 413949
rect 204364 413944 205607 413946
rect 204364 413888 205546 413944
rect 205602 413888 205607 413944
rect 204364 413886 205607 413888
rect 204364 413884 204370 413886
rect 205541 413883 205607 413886
rect 377489 413946 377555 413949
rect 377949 413946 378015 413949
rect 377489 413944 379530 413946
rect 377489 413888 377494 413944
rect 377550 413888 377954 413944
rect 378010 413888 379530 413944
rect 377489 413886 379530 413888
rect 377489 413883 377555 413886
rect 377949 413883 378015 413886
rect 379470 413844 379530 413886
rect 57881 413266 57947 413269
rect 60002 413266 60062 413814
rect 216857 413810 216923 413813
rect 219390 413810 220064 413844
rect 216857 413808 220064 413810
rect 216857 413752 216862 413808
rect 216918 413784 220064 413808
rect 379470 413784 380052 413844
rect 216918 413752 219450 413784
rect 216857 413750 219450 413752
rect 216857 413747 216923 413750
rect 57881 413264 60062 413266
rect 57881 413208 57886 413264
rect 57942 413208 60062 413264
rect 57881 413206 60062 413208
rect 57881 413203 57947 413206
rect 57881 411498 57947 411501
rect 60002 411498 60062 412046
rect 217685 412042 217751 412045
rect 219390 412042 220064 412076
rect 217685 412040 220064 412042
rect 217685 411984 217690 412040
rect 217746 412016 220064 412040
rect 377121 412042 377187 412045
rect 377489 412042 377555 412045
rect 379470 412042 380052 412076
rect 377121 412040 380052 412042
rect 217746 411984 219450 412016
rect 217685 411982 219450 411984
rect 377121 411984 377126 412040
rect 377182 411984 377494 412040
rect 377550 412016 380052 412040
rect 377550 411984 379530 412016
rect 377121 411982 379530 411984
rect 217685 411979 217751 411982
rect 377121 411979 377187 411982
rect 377489 411979 377555 411982
rect 57881 411496 60062 411498
rect 57881 411440 57886 411496
rect 57942 411440 60062 411496
rect 57881 411438 60062 411440
rect 57881 411435 57947 411438
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 56961 410410 57027 410413
rect 60002 410410 60062 410958
rect 216673 410954 216739 410957
rect 219390 410954 220064 410988
rect 216673 410952 220064 410954
rect 216673 410896 216678 410952
rect 216734 410928 220064 410952
rect 377213 410954 377279 410957
rect 377765 410954 377831 410957
rect 379470 410954 380052 410988
rect 377213 410952 380052 410954
rect 216734 410896 219450 410928
rect 216673 410894 219450 410896
rect 377213 410896 377218 410952
rect 377274 410896 377770 410952
rect 377826 410928 380052 410952
rect 377826 410896 379530 410928
rect 377213 410894 379530 410896
rect 216673 410891 216739 410894
rect 377213 410891 377279 410894
rect 377765 410891 377831 410894
rect 56961 410408 60062 410410
rect 56961 410352 56966 410408
rect 57022 410352 60062 410408
rect 56961 410350 60062 410352
rect 56961 410347 57027 410350
rect 57881 408642 57947 408645
rect 60002 408642 60062 409190
rect 217317 409186 217383 409189
rect 217869 409186 217935 409189
rect 219390 409186 220064 409220
rect 217317 409184 220064 409186
rect 217317 409128 217322 409184
rect 217378 409128 217874 409184
rect 217930 409160 220064 409184
rect 377397 409186 377463 409189
rect 378041 409186 378107 409189
rect 379470 409186 380052 409220
rect 377397 409184 380052 409186
rect 217930 409128 219450 409160
rect 217317 409126 219450 409128
rect 377397 409128 377402 409184
rect 377458 409128 378046 409184
rect 378102 409160 380052 409184
rect 378102 409128 379530 409160
rect 377397 409126 379530 409128
rect 217317 409123 217383 409126
rect 217869 409123 217935 409126
rect 377397 409123 377463 409126
rect 378041 409123 378107 409126
rect 57881 408640 60062 408642
rect 57881 408584 57886 408640
rect 57942 408584 60062 408640
rect 57881 408582 60062 408584
rect 57881 408579 57947 408582
rect 578877 404970 578943 404973
rect 583520 404970 584960 405060
rect 578877 404968 584960 404970
rect 578877 404912 578882 404968
rect 578938 404912 584960 404968
rect 578877 404910 584960 404912
rect 578877 404907 578943 404910
rect 583520 404820 584960 404910
rect 196558 400346 196618 400350
rect 199469 400346 199535 400349
rect 199837 400346 199903 400349
rect 196558 400344 199903 400346
rect 196558 400288 199474 400344
rect 199530 400288 199842 400344
rect 199898 400288 199903 400344
rect 196558 400286 199903 400288
rect 356562 400346 356622 400350
rect 359825 400346 359891 400349
rect 356562 400344 359891 400346
rect 356562 400288 359830 400344
rect 359886 400288 359891 400344
rect 356562 400286 359891 400288
rect 516558 400346 516618 400350
rect 518985 400346 519051 400349
rect 516558 400344 519051 400346
rect 516558 400288 518990 400344
rect 519046 400288 519051 400344
rect 516558 400286 519051 400288
rect 199469 400283 199535 400286
rect 199837 400283 199903 400286
rect 359825 400283 359891 400286
rect 518985 400283 519051 400286
rect 196558 397626 196618 398718
rect 356562 398170 356622 398718
rect 359089 398170 359155 398173
rect 356562 398168 359155 398170
rect 356562 398112 359094 398168
rect 359150 398112 359155 398168
rect 356562 398110 359155 398112
rect 516558 398170 516618 398718
rect 519077 398170 519143 398173
rect 516558 398168 519143 398170
rect 516558 398112 519082 398168
rect 519138 398112 519143 398168
rect 516558 398110 519143 398112
rect 359089 398107 359155 398110
rect 519077 398107 519143 398110
rect -960 397340 480 397580
rect 196558 397566 199026 397626
rect 198966 397493 199026 397566
rect 198966 397488 199075 397493
rect 198966 397432 199014 397488
rect 199070 397432 199075 397488
rect 198966 397430 199075 397432
rect 199009 397427 199075 397430
rect 196558 396810 196618 397358
rect 199653 396810 199719 396813
rect 196558 396808 199719 396810
rect 196558 396752 199658 396808
rect 199714 396752 199719 396808
rect 196558 396750 199719 396752
rect 356562 396810 356622 397358
rect 358997 396810 359063 396813
rect 356562 396808 359063 396810
rect 356562 396752 359002 396808
rect 359058 396752 359063 396808
rect 356562 396750 359063 396752
rect 516558 396810 516618 397358
rect 519261 396810 519327 396813
rect 516558 396808 519327 396810
rect 516558 396752 519266 396808
rect 519322 396752 519327 396808
rect 516558 396750 519327 396752
rect 199653 396747 199719 396750
rect 358997 396747 359063 396750
rect 519261 396747 519327 396750
rect 199285 395994 199351 395997
rect 199929 395994 199995 395997
rect 197126 395992 199995 395994
rect 197126 395936 199290 395992
rect 199346 395936 199934 395992
rect 199990 395936 199995 395992
rect 197126 395934 199995 395936
rect 197126 395892 197186 395934
rect 199285 395931 199351 395934
rect 199929 395931 199995 395934
rect 196604 395832 197186 395892
rect 356562 395314 356622 395862
rect 359181 395314 359247 395317
rect 356562 395312 359247 395314
rect 356562 395256 359186 395312
rect 359242 395256 359247 395312
rect 356562 395254 359247 395256
rect 516558 395314 516618 395862
rect 519169 395314 519235 395317
rect 516558 395312 519235 395314
rect 516558 395256 519174 395312
rect 519230 395256 519235 395312
rect 516558 395254 519235 395256
rect 359181 395251 359247 395254
rect 519169 395251 519235 395254
rect 196558 394634 196618 394638
rect 199377 394634 199443 394637
rect 199745 394634 199811 394637
rect 196558 394632 199811 394634
rect 196558 394576 199382 394632
rect 199438 394576 199750 394632
rect 199806 394576 199811 394632
rect 196558 394574 199811 394576
rect 199377 394571 199443 394574
rect 199745 394571 199811 394574
rect 356562 394090 356622 394638
rect 358905 394090 358971 394093
rect 356562 394088 358971 394090
rect 356562 394032 358910 394088
rect 358966 394032 358971 394088
rect 356562 394030 358971 394032
rect 516558 394090 516618 394638
rect 519353 394090 519419 394093
rect 516558 394088 519419 394090
rect 516558 394032 519358 394088
rect 519414 394032 519419 394088
rect 516558 394030 519419 394032
rect 358905 394027 358971 394030
rect 519353 394027 519419 394030
rect 583520 391628 584960 391868
rect 57881 391506 57947 391509
rect 57881 391504 60062 391506
rect 57881 391448 57886 391504
rect 57942 391448 60062 391504
rect 57881 391446 60062 391448
rect 57881 391443 57947 391446
rect 60002 390966 60062 391446
rect 216673 390962 216739 390965
rect 219390 390962 220064 390996
rect 216673 390960 220064 390962
rect 216673 390904 216678 390960
rect 216734 390936 220064 390960
rect 376937 390962 377003 390965
rect 379470 390962 380052 390996
rect 376937 390960 380052 390962
rect 216734 390904 219450 390936
rect 216673 390902 219450 390904
rect 376937 390904 376942 390960
rect 376998 390936 380052 390960
rect 376998 390904 379530 390936
rect 376937 390902 379530 390904
rect 216673 390899 216739 390902
rect 376937 390899 377003 390902
rect 208342 390628 208348 390692
rect 208412 390690 208418 390692
rect 209681 390690 209747 390693
rect 208412 390688 209747 390690
rect 208412 390632 209686 390688
rect 209742 390632 209747 390688
rect 208412 390630 209747 390632
rect 208412 390628 208418 390630
rect 209681 390627 209747 390630
rect 57605 389738 57671 389741
rect 57605 389736 60062 389738
rect 57605 389680 57610 389736
rect 57666 389680 60062 389736
rect 57605 389678 60062 389680
rect 57605 389675 57671 389678
rect 60002 389334 60062 389678
rect 216673 389330 216739 389333
rect 219390 389330 220064 389364
rect 216673 389328 220064 389330
rect 216673 389272 216678 389328
rect 216734 389304 220064 389328
rect 376937 389330 377003 389333
rect 379470 389330 380052 389364
rect 376937 389328 380052 389330
rect 216734 389272 219450 389304
rect 216673 389270 219450 389272
rect 376937 389272 376942 389328
rect 376998 389304 380052 389328
rect 376998 389272 379530 389304
rect 376937 389270 379530 389272
rect 216673 389267 216739 389270
rect 376937 389267 377003 389270
rect 57605 389058 57671 389061
rect 60002 389058 60062 389062
rect 57605 389056 60062 389058
rect 57605 389000 57610 389056
rect 57666 389000 60062 389056
rect 57605 388998 60062 389000
rect 216673 389058 216739 389061
rect 219390 389058 220064 389092
rect 216673 389056 220064 389058
rect 216673 389000 216678 389056
rect 216734 389032 220064 389056
rect 376937 389058 377003 389061
rect 379470 389058 380052 389092
rect 376937 389056 380052 389058
rect 216734 389000 219450 389032
rect 216673 388998 219450 389000
rect 376937 389000 376942 389056
rect 376998 389032 380052 389056
rect 376998 389000 379530 389032
rect 376937 388998 379530 389000
rect 57605 388995 57671 388998
rect 216673 388995 216739 388998
rect 376937 388995 377003 388998
rect 56685 388650 56751 388653
rect 57646 388650 57652 388652
rect 56685 388648 57652 388650
rect 56685 388592 56690 388648
rect 56746 388592 57652 388648
rect 56685 388590 57652 388592
rect 56685 388587 56751 388590
rect 57646 388588 57652 388590
rect 57716 388588 57722 388652
rect 57646 388452 57652 388516
rect 57716 388514 57722 388516
rect 58525 388514 58591 388517
rect 57716 388512 58591 388514
rect 57716 388456 58530 388512
rect 58586 388456 58591 388512
rect 57716 388454 58591 388456
rect 57716 388452 57722 388454
rect 58525 388451 58591 388454
rect -960 384284 480 384524
rect 198406 380972 198412 381036
rect 198476 381034 198482 381036
rect 198641 381034 198707 381037
rect 198476 381032 198707 381034
rect 198476 380976 198646 381032
rect 198702 380976 198707 381032
rect 198476 380974 198707 380976
rect 198476 380972 198482 380974
rect 198641 380971 198707 380974
rect 210734 380972 210740 381036
rect 210804 381034 210810 381036
rect 212901 381034 212967 381037
rect 376937 381036 377003 381037
rect 376886 381034 376892 381036
rect 210804 381032 212967 381034
rect 210804 380976 212906 381032
rect 212962 380976 212967 381032
rect 210804 380974 212967 380976
rect 376846 380974 376892 381034
rect 376956 381032 377003 381036
rect 376998 380976 377003 381032
rect 210804 380972 210810 380974
rect 212901 380971 212967 380974
rect 376886 380972 376892 380974
rect 376956 380972 377003 380976
rect 376937 380971 377003 380972
rect 52361 380898 52427 380901
rect 217869 380898 217935 380901
rect 52361 380896 217935 380898
rect 52361 380840 52366 380896
rect 52422 380840 217874 380896
rect 217930 380840 217935 380896
rect 52361 380838 217935 380840
rect 52361 380835 52427 380838
rect 217869 380835 217935 380838
rect 235993 380900 236059 380901
rect 237097 380900 237163 380901
rect 243077 380900 243143 380901
rect 245377 380900 245443 380901
rect 247585 380900 247651 380901
rect 254485 380900 254551 380901
rect 255865 380900 255931 380901
rect 256969 380900 257035 380901
rect 276013 380900 276079 380901
rect 235993 380896 236054 380900
rect 235993 380840 235998 380896
rect 235993 380836 236054 380840
rect 236118 380898 236124 380900
rect 236118 380838 236150 380898
rect 237097 380896 237142 380900
rect 237206 380898 237212 380900
rect 237097 380840 237102 380896
rect 236118 380836 236124 380838
rect 237097 380836 237142 380840
rect 237206 380838 237254 380898
rect 243077 380896 243126 380900
rect 243190 380898 243196 380900
rect 243077 380840 243082 380896
rect 237206 380836 237212 380838
rect 243077 380836 243126 380840
rect 243190 380838 243234 380898
rect 245377 380896 245438 380900
rect 245377 380840 245382 380896
rect 243190 380836 243196 380838
rect 245377 380836 245438 380840
rect 245502 380898 245508 380900
rect 245502 380838 245534 380898
rect 247585 380896 247614 380900
rect 247678 380898 247684 380900
rect 247585 380840 247590 380896
rect 245502 380836 245508 380838
rect 247585 380836 247614 380840
rect 247678 380838 247742 380898
rect 254485 380896 254550 380900
rect 254485 380840 254490 380896
rect 254546 380840 254550 380896
rect 247678 380836 247684 380838
rect 254485 380836 254550 380840
rect 254614 380898 254620 380900
rect 254614 380838 254642 380898
rect 255865 380896 255910 380900
rect 255974 380898 255980 380900
rect 255865 380840 255870 380896
rect 254614 380836 254620 380838
rect 255865 380836 255910 380840
rect 255974 380838 256022 380898
rect 256969 380896 256998 380900
rect 257062 380898 257068 380900
rect 269776 380898 269782 380900
rect 256969 380840 256974 380896
rect 255974 380836 255980 380838
rect 256969 380836 256998 380840
rect 257062 380838 257126 380898
rect 267690 380838 269782 380898
rect 257062 380836 257068 380838
rect 235993 380835 236059 380836
rect 237097 380835 237163 380836
rect 243077 380835 243143 380836
rect 245377 380835 245443 380836
rect 247585 380835 247651 380836
rect 254485 380835 254551 380836
rect 255865 380835 255931 380836
rect 256969 380835 257035 380836
rect 76048 380700 76054 380764
rect 76118 380762 76124 380764
rect 202873 380762 202939 380765
rect 76118 380760 202939 380762
rect 76118 380704 202878 380760
rect 202934 380704 202939 380760
rect 76118 380702 202939 380704
rect 76118 380700 76124 380702
rect 202873 380699 202939 380702
rect 215477 380762 215543 380765
rect 216581 380762 216647 380765
rect 263928 380762 263934 380764
rect 215477 380760 263934 380762
rect 215477 380704 215482 380760
rect 215538 380704 216586 380760
rect 216642 380704 263934 380760
rect 215477 380702 263934 380704
rect 215477 380699 215543 380702
rect 216581 380699 216647 380702
rect 263928 380700 263934 380702
rect 263998 380700 264004 380764
rect 83120 380564 83126 380628
rect 83190 380626 83196 380628
rect 207013 380626 207079 380629
rect 83190 380624 207079 380626
rect 83190 380568 207018 380624
rect 207074 380568 207079 380624
rect 83190 380566 207079 380568
rect 83190 380564 83196 380566
rect 207013 380563 207079 380566
rect 207933 380626 207999 380629
rect 212625 380626 212691 380629
rect 259453 380628 259519 380629
rect 265249 380628 265315 380629
rect 258080 380626 258086 380628
rect 207933 380624 258086 380626
rect 207933 380568 207938 380624
rect 207994 380568 212630 380624
rect 212686 380568 258086 380624
rect 207933 380566 258086 380568
rect 207933 380563 207999 380566
rect 212625 380563 212691 380566
rect 258080 380564 258086 380566
rect 258150 380564 258156 380628
rect 259440 380626 259446 380628
rect 259362 380566 259446 380626
rect 259510 380624 259519 380628
rect 259514 380568 259519 380624
rect 259440 380564 259446 380566
rect 259510 380564 259519 380568
rect 260664 380564 260670 380628
rect 260734 380564 260740 380628
rect 265249 380624 265294 380628
rect 265358 380626 265364 380628
rect 265249 380568 265254 380624
rect 265249 380564 265294 380568
rect 265358 380566 265406 380626
rect 265358 380564 265364 380566
rect 259453 380563 259519 380564
rect 84510 380428 84516 380492
rect 84580 380490 84586 380492
rect 208393 380490 208459 380493
rect 84580 380488 208459 380490
rect 84580 380432 208398 380488
rect 208454 380432 208459 380488
rect 84580 380430 208459 380432
rect 84580 380428 84586 380430
rect 208393 380427 208459 380430
rect 216622 380428 216628 380492
rect 216692 380490 216698 380492
rect 216990 380490 216996 380492
rect 216692 380430 216996 380490
rect 216692 380428 216698 380430
rect 216990 380428 216996 380430
rect 217060 380490 217066 380492
rect 260672 380490 260732 380564
rect 265249 380563 265315 380564
rect 217060 380430 260732 380490
rect 217060 380428 217066 380430
rect 105813 380356 105879 380357
rect 110965 380356 111031 380357
rect 113541 380356 113607 380357
rect 115933 380356 115999 380357
rect 118325 380356 118391 380357
rect 120901 380356 120967 380357
rect 123569 380356 123635 380357
rect 128353 380356 128419 380357
rect 133505 380356 133571 380357
rect 135897 380356 135963 380357
rect 138473 380356 138539 380357
rect 148593 380356 148659 380357
rect 155953 380356 156019 380357
rect 158529 380356 158595 380357
rect 160921 380356 160987 380357
rect 163497 380356 163563 380357
rect 166073 380356 166139 380357
rect 105813 380352 105860 380356
rect 105924 380354 105930 380356
rect 105813 380296 105818 380352
rect 105813 380292 105860 380296
rect 105924 380294 105970 380354
rect 110965 380352 111012 380356
rect 111076 380354 111082 380356
rect 110965 380296 110970 380352
rect 105924 380292 105930 380294
rect 110965 380292 111012 380296
rect 111076 380294 111122 380354
rect 113541 380352 113588 380356
rect 113652 380354 113658 380356
rect 113541 380296 113546 380352
rect 111076 380292 111082 380294
rect 113541 380292 113588 380296
rect 113652 380294 113698 380354
rect 115933 380352 115980 380356
rect 116044 380354 116050 380356
rect 115933 380296 115938 380352
rect 113652 380292 113658 380294
rect 115933 380292 115980 380296
rect 116044 380294 116090 380354
rect 118325 380352 118372 380356
rect 118436 380354 118442 380356
rect 118325 380296 118330 380352
rect 116044 380292 116050 380294
rect 118325 380292 118372 380296
rect 118436 380294 118482 380354
rect 120901 380352 120948 380356
rect 121012 380354 121018 380356
rect 123518 380354 123524 380356
rect 120901 380296 120906 380352
rect 118436 380292 118442 380294
rect 120901 380292 120948 380296
rect 121012 380294 121058 380354
rect 123478 380294 123524 380354
rect 123588 380352 123635 380356
rect 128302 380354 128308 380356
rect 123630 380296 123635 380352
rect 121012 380292 121018 380294
rect 123518 380292 123524 380294
rect 123588 380292 123635 380296
rect 128262 380294 128308 380354
rect 128372 380352 128419 380356
rect 133454 380354 133460 380356
rect 128414 380296 128419 380352
rect 128302 380292 128308 380294
rect 128372 380292 128419 380296
rect 133414 380294 133460 380354
rect 133524 380352 133571 380356
rect 135846 380354 135852 380356
rect 133566 380296 133571 380352
rect 133454 380292 133460 380294
rect 133524 380292 133571 380296
rect 135806 380294 135852 380354
rect 135916 380352 135963 380356
rect 138422 380354 138428 380356
rect 135958 380296 135963 380352
rect 135846 380292 135852 380294
rect 135916 380292 135963 380296
rect 138382 380294 138428 380354
rect 138492 380352 138539 380356
rect 148542 380354 148548 380356
rect 138534 380296 138539 380352
rect 138422 380292 138428 380294
rect 138492 380292 138539 380296
rect 148502 380294 148548 380354
rect 148612 380352 148659 380356
rect 155902 380354 155908 380356
rect 148654 380296 148659 380352
rect 148542 380292 148548 380294
rect 148612 380292 148659 380296
rect 155862 380294 155908 380354
rect 155972 380352 156019 380356
rect 158478 380354 158484 380356
rect 156014 380296 156019 380352
rect 155902 380292 155908 380294
rect 155972 380292 156019 380296
rect 158438 380294 158484 380354
rect 158548 380352 158595 380356
rect 160870 380354 160876 380356
rect 158590 380296 158595 380352
rect 158478 380292 158484 380294
rect 158548 380292 158595 380296
rect 160830 380294 160876 380354
rect 160940 380352 160987 380356
rect 163446 380354 163452 380356
rect 160982 380296 160987 380352
rect 160870 380292 160876 380294
rect 160940 380292 160987 380296
rect 163406 380294 163452 380354
rect 163516 380352 163563 380356
rect 166022 380354 166028 380356
rect 163558 380296 163563 380352
rect 163446 380292 163452 380294
rect 163516 380292 163563 380296
rect 165982 380294 166028 380354
rect 166092 380352 166139 380356
rect 166134 380296 166139 380352
rect 166022 380292 166028 380294
rect 166092 380292 166139 380296
rect 105813 380291 105879 380292
rect 110965 380291 111031 380292
rect 113541 380291 113607 380292
rect 115933 380291 115999 380292
rect 118325 380291 118391 380292
rect 120901 380291 120967 380292
rect 123569 380291 123635 380292
rect 128353 380291 128419 380292
rect 133505 380291 133571 380292
rect 135897 380291 135963 380292
rect 138473 380291 138539 380292
rect 148593 380291 148659 380292
rect 155953 380291 156019 380292
rect 158529 380291 158595 380292
rect 160921 380291 160987 380292
rect 163497 380291 163563 380292
rect 166073 380291 166139 380292
rect 203885 380354 203951 380357
rect 218513 380354 218579 380357
rect 244273 380356 244339 380357
rect 244222 380354 244228 380356
rect 203885 380352 218579 380354
rect 203885 380296 203890 380352
rect 203946 380296 218518 380352
rect 218574 380296 218579 380352
rect 203885 380294 218579 380296
rect 244182 380294 244228 380354
rect 244292 380352 244339 380356
rect 244334 380296 244339 380352
rect 203885 380291 203951 380294
rect 218513 380291 218579 380294
rect 244222 380292 244228 380294
rect 244292 380292 244339 380296
rect 244273 380291 244339 380292
rect 119102 380156 119108 380220
rect 119172 380218 119178 380220
rect 207013 380218 207079 380221
rect 119172 380216 207079 380218
rect 119172 380160 207018 380216
rect 207074 380160 207079 380216
rect 119172 380158 207079 380160
rect 119172 380156 119178 380158
rect 207013 380155 207079 380158
rect 51758 379476 51764 379540
rect 51828 379538 51834 379540
rect 52269 379538 52335 379541
rect 51828 379536 52335 379538
rect 51828 379480 52274 379536
rect 52330 379480 52335 379536
rect 51828 379478 52335 379480
rect 51828 379476 51834 379478
rect 52269 379475 52335 379478
rect 200982 379476 200988 379540
rect 201052 379538 201058 379540
rect 201309 379538 201375 379541
rect 201052 379536 201375 379538
rect 201052 379480 201314 379536
rect 201370 379480 201375 379536
rect 201052 379478 201375 379480
rect 201052 379476 201058 379478
rect 201309 379475 201375 379478
rect 202454 379476 202460 379540
rect 202524 379538 202530 379540
rect 202781 379538 202847 379541
rect 202524 379536 202847 379538
rect 202524 379480 202786 379536
rect 202842 379480 202847 379536
rect 202524 379478 202847 379480
rect 202524 379476 202530 379478
rect 202781 379475 202847 379478
rect 206185 379538 206251 379541
rect 206318 379538 206324 379540
rect 206185 379536 206324 379538
rect 206185 379480 206190 379536
rect 206246 379480 206324 379536
rect 206185 379478 206324 379480
rect 206185 379475 206251 379478
rect 206318 379476 206324 379478
rect 206388 379476 206394 379540
rect 217133 379538 217199 379541
rect 217869 379538 217935 379541
rect 217133 379536 217935 379538
rect 217133 379480 217138 379536
rect 217194 379480 217874 379536
rect 217930 379480 217935 379536
rect 217133 379478 217935 379480
rect 217133 379475 217199 379478
rect 217869 379475 217935 379478
rect 218053 379538 218119 379541
rect 218053 379536 218162 379538
rect 218053 379480 218058 379536
rect 218114 379480 218162 379536
rect 218053 379475 218162 379480
rect 46105 379402 46171 379405
rect 78254 379402 78260 379404
rect 46105 379400 78260 379402
rect 46105 379344 46110 379400
rect 46166 379344 78260 379400
rect 46105 379342 78260 379344
rect 46105 379339 46171 379342
rect 78254 379340 78260 379342
rect 78324 379340 78330 379404
rect 80329 379402 80395 379405
rect 85481 379404 85547 379405
rect 86585 379404 86651 379405
rect 87689 379404 87755 379405
rect 80462 379402 80468 379404
rect 80329 379400 80468 379402
rect 80329 379344 80334 379400
rect 80390 379344 80468 379400
rect 80329 379342 80468 379344
rect 80329 379339 80395 379342
rect 80462 379340 80468 379342
rect 80532 379340 80538 379404
rect 85430 379402 85436 379404
rect 85390 379342 85436 379402
rect 85500 379400 85547 379404
rect 86534 379402 86540 379404
rect 85542 379344 85547 379400
rect 85430 379340 85436 379342
rect 85500 379340 85547 379344
rect 86494 379342 86540 379402
rect 86604 379400 86651 379404
rect 87638 379402 87644 379404
rect 86646 379344 86651 379400
rect 86534 379340 86540 379342
rect 86604 379340 86651 379344
rect 87598 379342 87644 379402
rect 87708 379400 87755 379404
rect 87750 379344 87755 379400
rect 87638 379340 87644 379342
rect 87708 379340 87755 379344
rect 85481 379339 85547 379340
rect 86585 379339 86651 379340
rect 87689 379339 87755 379340
rect 88333 379404 88399 379405
rect 88793 379404 88859 379405
rect 88333 379400 88380 379404
rect 88444 379402 88450 379404
rect 88742 379402 88748 379404
rect 88333 379344 88338 379400
rect 88333 379340 88380 379344
rect 88444 379342 88490 379402
rect 88702 379342 88748 379402
rect 88812 379400 88859 379404
rect 88854 379344 88859 379400
rect 88444 379340 88450 379342
rect 88742 379340 88748 379342
rect 88812 379340 88859 379344
rect 88333 379339 88399 379340
rect 88793 379339 88859 379340
rect 90633 379402 90699 379405
rect 91369 379404 91435 379405
rect 90766 379402 90772 379404
rect 90633 379400 90772 379402
rect 90633 379344 90638 379400
rect 90694 379344 90772 379400
rect 90633 379342 90772 379344
rect 90633 379339 90699 379342
rect 90766 379340 90772 379342
rect 90836 379340 90842 379404
rect 91318 379402 91324 379404
rect 91278 379342 91324 379402
rect 91388 379400 91435 379404
rect 91430 379344 91435 379400
rect 91318 379340 91324 379342
rect 91388 379340 91435 379344
rect 91369 379339 91435 379340
rect 92381 379404 92447 379405
rect 92381 379400 92428 379404
rect 92492 379402 92498 379404
rect 92381 379344 92386 379400
rect 92381 379340 92428 379344
rect 92492 379342 92538 379402
rect 92492 379340 92498 379342
rect 93342 379340 93348 379404
rect 93412 379402 93418 379404
rect 93577 379402 93643 379405
rect 93412 379400 93643 379402
rect 93412 379344 93582 379400
rect 93638 379344 93643 379400
rect 93412 379342 93643 379344
rect 93412 379340 93418 379342
rect 92381 379339 92447 379340
rect 93577 379339 93643 379342
rect 96061 379404 96127 379405
rect 96061 379400 96108 379404
rect 96172 379402 96178 379404
rect 98177 379402 98243 379405
rect 101029 379404 101095 379405
rect 98494 379402 98500 379404
rect 96061 379344 96066 379400
rect 96061 379340 96108 379344
rect 96172 379342 96218 379402
rect 98177 379400 98500 379402
rect 98177 379344 98182 379400
rect 98238 379344 98500 379400
rect 98177 379342 98500 379344
rect 96172 379340 96178 379342
rect 96061 379339 96127 379340
rect 98177 379339 98243 379342
rect 98494 379340 98500 379342
rect 98564 379340 98570 379404
rect 101029 379400 101076 379404
rect 101140 379402 101146 379404
rect 101029 379344 101034 379400
rect 101029 379340 101076 379344
rect 101140 379342 101186 379402
rect 101140 379340 101146 379342
rect 103278 379340 103284 379404
rect 103348 379402 103354 379404
rect 103513 379402 103579 379405
rect 105353 379404 105419 379405
rect 105302 379402 105308 379404
rect 103348 379400 103579 379402
rect 103348 379344 103518 379400
rect 103574 379344 103579 379400
rect 103348 379342 103579 379344
rect 105262 379342 105308 379402
rect 105372 379400 105419 379404
rect 105414 379344 105419 379400
rect 103348 379340 103354 379342
rect 101029 379339 101095 379340
rect 103513 379339 103579 379342
rect 105302 379340 105308 379342
rect 105372 379340 105419 379344
rect 105353 379339 105419 379340
rect 108205 379404 108271 379405
rect 108849 379404 108915 379405
rect 111241 379404 111307 379405
rect 112345 379404 112411 379405
rect 113449 379404 113515 379405
rect 108205 379400 108252 379404
rect 108316 379402 108322 379404
rect 108798 379402 108804 379404
rect 108205 379344 108210 379400
rect 108205 379340 108252 379344
rect 108316 379342 108362 379402
rect 108758 379342 108804 379402
rect 108868 379400 108915 379404
rect 111190 379402 111196 379404
rect 108910 379344 108915 379400
rect 108316 379340 108322 379342
rect 108798 379340 108804 379342
rect 108868 379340 108915 379344
rect 111150 379342 111196 379402
rect 111260 379400 111307 379404
rect 112294 379402 112300 379404
rect 111302 379344 111307 379400
rect 111190 379340 111196 379342
rect 111260 379340 111307 379344
rect 112254 379342 112300 379402
rect 112364 379400 112411 379404
rect 113398 379402 113404 379404
rect 112406 379344 112411 379400
rect 112294 379340 112300 379342
rect 112364 379340 112411 379344
rect 113358 379342 113404 379402
rect 113468 379400 113515 379404
rect 113510 379344 113515 379400
rect 113398 379340 113404 379342
rect 113468 379340 113515 379344
rect 108205 379339 108271 379340
rect 108849 379339 108915 379340
rect 111241 379339 111307 379340
rect 112345 379339 112411 379340
rect 113449 379339 113515 379340
rect 114461 379404 114527 379405
rect 115841 379404 115907 379405
rect 141049 379404 141115 379405
rect 143625 379404 143691 379405
rect 146017 379404 146083 379405
rect 150985 379404 151051 379405
rect 153561 379404 153627 379405
rect 114461 379400 114508 379404
rect 114572 379402 114578 379404
rect 115790 379402 115796 379404
rect 114461 379344 114466 379400
rect 114461 379340 114508 379344
rect 114572 379342 114618 379402
rect 115750 379342 115796 379402
rect 115860 379400 115907 379404
rect 140998 379402 141004 379404
rect 115902 379344 115907 379400
rect 114572 379340 114578 379342
rect 115790 379340 115796 379342
rect 115860 379340 115907 379344
rect 140958 379342 141004 379402
rect 141068 379400 141115 379404
rect 143574 379402 143580 379404
rect 141110 379344 141115 379400
rect 140998 379340 141004 379342
rect 141068 379340 141115 379344
rect 143534 379342 143580 379402
rect 143644 379400 143691 379404
rect 145966 379402 145972 379404
rect 143686 379344 143691 379400
rect 143574 379340 143580 379342
rect 143644 379340 143691 379344
rect 145926 379342 145972 379402
rect 146036 379400 146083 379404
rect 150934 379402 150940 379404
rect 146078 379344 146083 379400
rect 145966 379340 145972 379342
rect 146036 379340 146083 379344
rect 150894 379342 150940 379402
rect 151004 379400 151051 379404
rect 153510 379402 153516 379404
rect 151046 379344 151051 379400
rect 150934 379340 150940 379342
rect 151004 379340 151051 379344
rect 153470 379342 153516 379402
rect 153580 379400 153627 379404
rect 153622 379344 153627 379400
rect 153510 379340 153516 379342
rect 153580 379340 153627 379344
rect 114461 379339 114527 379340
rect 115841 379339 115907 379340
rect 141049 379339 141115 379340
rect 143625 379339 143691 379340
rect 146017 379339 146083 379340
rect 150985 379339 151051 379340
rect 153561 379339 153627 379340
rect 199009 379402 199075 379405
rect 199142 379402 199148 379404
rect 199009 379400 199148 379402
rect 199009 379344 199014 379400
rect 199070 379344 199148 379400
rect 199009 379342 199148 379344
rect 199009 379339 199075 379342
rect 199142 379340 199148 379342
rect 199212 379340 199218 379404
rect 47485 379266 47551 379269
rect 79542 379266 79548 379268
rect 47485 379264 79548 379266
rect 47485 379208 47490 379264
rect 47546 379208 79548 379264
rect 47485 379206 79548 379208
rect 47485 379203 47551 379206
rect 79542 379204 79548 379206
rect 79612 379266 79618 379268
rect 79612 379206 84210 379266
rect 79612 379204 79618 379206
rect 84150 379130 84210 379206
rect 90030 379204 90036 379268
rect 90100 379266 90106 379268
rect 90725 379266 90791 379269
rect 90100 379264 90791 379266
rect 90100 379208 90730 379264
rect 90786 379208 90791 379264
rect 90100 379206 90791 379208
rect 90100 379204 90106 379206
rect 90725 379203 90791 379206
rect 93485 379266 93551 379269
rect 95969 379268 96035 379269
rect 93710 379266 93716 379268
rect 93485 379264 93716 379266
rect 93485 379208 93490 379264
rect 93546 379208 93716 379264
rect 93485 379206 93716 379208
rect 93485 379203 93551 379206
rect 93710 379204 93716 379206
rect 93780 379204 93786 379268
rect 95918 379266 95924 379268
rect 95878 379206 95924 379266
rect 95988 379264 96035 379268
rect 96030 379208 96035 379264
rect 95918 379204 95924 379206
rect 95988 379204 96035 379208
rect 98126 379204 98132 379268
rect 98196 379266 98202 379268
rect 98361 379266 98427 379269
rect 99465 379268 99531 379269
rect 102961 379268 103027 379269
rect 99414 379266 99420 379268
rect 98196 379264 98427 379266
rect 98196 379208 98366 379264
rect 98422 379208 98427 379264
rect 98196 379206 98427 379208
rect 99374 379206 99420 379266
rect 99484 379264 99531 379268
rect 102910 379266 102916 379268
rect 99526 379208 99531 379264
rect 98196 379204 98202 379206
rect 95969 379203 96035 379204
rect 98361 379203 98427 379206
rect 99414 379204 99420 379206
rect 99484 379204 99531 379208
rect 102870 379206 102916 379266
rect 102980 379264 103027 379268
rect 103022 379208 103027 379264
rect 102910 379204 102916 379206
rect 102980 379204 103027 379208
rect 109718 379204 109724 379268
rect 109788 379266 109794 379268
rect 109788 379206 208778 379266
rect 109788 379204 109794 379206
rect 99465 379203 99531 379204
rect 102961 379203 103027 379204
rect 208485 379130 208551 379133
rect 84150 379128 208551 379130
rect 84150 379072 208490 379128
rect 208546 379072 208551 379128
rect 84150 379070 208551 379072
rect 208718 379130 208778 379206
rect 209814 379204 209820 379268
rect 209884 379266 209890 379268
rect 210969 379266 211035 379269
rect 209884 379264 211035 379266
rect 209884 379208 210974 379264
rect 211030 379208 211035 379264
rect 209884 379206 211035 379208
rect 209884 379204 209890 379206
rect 210969 379203 211035 379206
rect 209497 379130 209563 379133
rect 218102 379130 218162 379475
rect 267690 379402 267750 380838
rect 269776 380836 269782 380838
rect 269846 380836 269852 380900
rect 276013 380896 276038 380900
rect 276102 380898 276108 380900
rect 370405 380898 370471 380901
rect 485944 380898 485950 380900
rect 276013 380840 276018 380896
rect 276013 380836 276038 380840
rect 276102 380838 276170 380898
rect 370405 380896 485950 380898
rect 370405 380840 370410 380896
rect 370466 380840 485950 380896
rect 370405 380838 485950 380840
rect 276102 380836 276108 380838
rect 276013 380835 276079 380836
rect 370405 380835 370471 380838
rect 485944 380836 485950 380838
rect 486014 380836 486020 380900
rect 421097 380764 421163 380765
rect 421072 380762 421078 380764
rect 421006 380702 421078 380762
rect 421142 380760 421163 380764
rect 421158 380704 421163 380760
rect 421072 380700 421078 380702
rect 421142 380700 421163 380704
rect 421097 380699 421163 380700
rect 421741 380764 421807 380765
rect 425973 380764 426039 380765
rect 433609 380764 433675 380765
rect 421741 380760 421758 380764
rect 421822 380762 421828 380764
rect 425968 380762 425974 380764
rect 421741 380704 421746 380760
rect 421741 380700 421758 380704
rect 421822 380702 421898 380762
rect 425882 380702 425974 380762
rect 421822 380700 421828 380702
rect 425968 380700 425974 380702
rect 426038 380700 426044 380764
rect 433584 380762 433590 380764
rect 433518 380702 433590 380762
rect 433654 380760 433675 380764
rect 433670 380704 433675 380760
rect 433584 380700 433590 380702
rect 433654 380700 433675 380704
rect 421741 380699 421807 380700
rect 425973 380699 426039 380700
rect 433609 380699 433675 380700
rect 434345 380764 434411 380765
rect 436001 380764 436067 380765
rect 438485 380764 438551 380765
rect 440877 380764 440943 380765
rect 443453 380764 443519 380765
rect 434345 380760 434406 380764
rect 434345 380704 434350 380760
rect 434345 380700 434406 380704
rect 434470 380762 434476 380764
rect 434470 380702 434502 380762
rect 436001 380760 436038 380764
rect 436102 380762 436108 380764
rect 438480 380762 438486 380764
rect 436001 380704 436006 380760
rect 434470 380700 434476 380702
rect 436001 380700 436038 380704
rect 436102 380702 436158 380762
rect 438394 380702 438486 380762
rect 436102 380700 436108 380702
rect 438480 380700 438486 380702
rect 438550 380700 438556 380764
rect 440877 380760 440934 380764
rect 440998 380762 441004 380764
rect 440877 380704 440882 380760
rect 440877 380700 440934 380704
rect 440998 380702 441034 380762
rect 443453 380760 443518 380764
rect 443453 380704 443458 380760
rect 443514 380704 443518 380760
rect 440998 380700 441004 380702
rect 443453 380700 443518 380704
rect 443582 380762 443588 380764
rect 443582 380702 443610 380762
rect 443582 380700 443588 380702
rect 434345 380699 434411 380700
rect 436001 380699 436067 380700
rect 438485 380699 438551 380700
rect 440877 380699 440943 380700
rect 443453 380699 443519 380700
rect 270953 380628 271019 380629
rect 408677 380628 408743 380629
rect 413461 380628 413527 380629
rect 422845 380628 422911 380629
rect 425237 380628 425303 380629
rect 436921 380628 436987 380629
rect 465901 380628 465967 380629
rect 270953 380624 271006 380628
rect 271070 380626 271076 380628
rect 270953 380568 270958 380624
rect 270953 380564 271006 380568
rect 271070 380566 271110 380626
rect 408677 380624 408702 380628
rect 408766 380626 408772 380628
rect 413456 380626 413462 380628
rect 408677 380568 408682 380624
rect 271070 380564 271076 380566
rect 408677 380564 408702 380568
rect 408766 380566 408834 380626
rect 413370 380566 413462 380626
rect 408766 380564 408772 380566
rect 413456 380564 413462 380566
rect 413526 380564 413532 380628
rect 422840 380626 422846 380628
rect 422754 380566 422846 380626
rect 422840 380564 422846 380566
rect 422910 380564 422916 380628
rect 425237 380624 425294 380628
rect 425358 380626 425364 380628
rect 425237 380568 425242 380624
rect 425237 380564 425294 380568
rect 425358 380566 425394 380626
rect 436921 380624 436990 380628
rect 436921 380568 436926 380624
rect 436982 380568 436990 380624
rect 425358 380564 425364 380566
rect 436921 380564 436990 380568
rect 437054 380626 437060 380628
rect 437054 380566 437078 380626
rect 465901 380624 465958 380628
rect 466022 380626 466028 380628
rect 465901 380568 465906 380624
rect 437054 380564 437060 380566
rect 465901 380564 465958 380568
rect 466022 380566 466058 380626
rect 466022 380564 466028 380566
rect 270953 380563 271019 380564
rect 408677 380563 408743 380564
rect 413461 380563 413527 380564
rect 422845 380563 422911 380564
rect 425237 380563 425303 380564
rect 436921 380563 436987 380564
rect 465901 380563 465967 380564
rect 376569 379538 376635 379541
rect 376886 379538 376892 379540
rect 376569 379536 376892 379538
rect 376569 379480 376574 379536
rect 376630 379480 376892 379536
rect 376569 379478 376892 379480
rect 376569 379475 376635 379478
rect 376886 379476 376892 379478
rect 376956 379476 376962 379540
rect 238710 379342 267750 379402
rect 268653 379404 268719 379405
rect 271045 379404 271111 379405
rect 268653 379400 268700 379404
rect 268764 379402 268770 379404
rect 268653 379344 268658 379400
rect 238710 379266 238770 379342
rect 268653 379340 268700 379344
rect 268764 379342 268810 379402
rect 271045 379400 271092 379404
rect 271156 379402 271162 379404
rect 271965 379402 272031 379405
rect 273253 379404 273319 379405
rect 274357 379404 274423 379405
rect 275645 379404 275711 379405
rect 285949 379404 286015 379405
rect 272190 379402 272196 379404
rect 271045 379344 271050 379400
rect 268764 379340 268770 379342
rect 271045 379340 271092 379344
rect 271156 379342 271202 379402
rect 271965 379400 272196 379402
rect 271965 379344 271970 379400
rect 272026 379344 272196 379400
rect 271965 379342 272196 379344
rect 271156 379340 271162 379342
rect 268653 379339 268719 379340
rect 271045 379339 271111 379340
rect 271965 379339 272031 379342
rect 272190 379340 272196 379342
rect 272260 379340 272266 379404
rect 273253 379400 273300 379404
rect 273364 379402 273370 379404
rect 273253 379344 273258 379400
rect 273253 379340 273300 379344
rect 273364 379342 273410 379402
rect 274357 379400 274404 379404
rect 274468 379402 274474 379404
rect 274357 379344 274362 379400
rect 273364 379340 273370 379342
rect 274357 379340 274404 379344
rect 274468 379342 274514 379402
rect 275645 379400 275692 379404
rect 275756 379402 275762 379404
rect 275645 379344 275650 379400
rect 274468 379340 274474 379342
rect 275645 379340 275692 379344
rect 275756 379342 275802 379402
rect 285949 379400 285996 379404
rect 286060 379402 286066 379404
rect 287605 379402 287671 379405
rect 290917 379404 290983 379405
rect 293309 379404 293375 379405
rect 295885 379404 295951 379405
rect 288198 379402 288204 379404
rect 285949 379344 285954 379400
rect 275756 379340 275762 379342
rect 285949 379340 285996 379344
rect 286060 379342 286106 379402
rect 287605 379400 288204 379402
rect 287605 379344 287610 379400
rect 287666 379344 288204 379400
rect 287605 379342 288204 379344
rect 286060 379340 286066 379342
rect 273253 379339 273319 379340
rect 274357 379339 274423 379340
rect 275645 379339 275711 379340
rect 285949 379339 286015 379340
rect 287605 379339 287671 379342
rect 288198 379340 288204 379342
rect 288268 379340 288274 379404
rect 290917 379400 290964 379404
rect 291028 379402 291034 379404
rect 290917 379344 290922 379400
rect 290917 379340 290964 379344
rect 291028 379342 291074 379402
rect 293309 379400 293356 379404
rect 293420 379402 293426 379404
rect 293309 379344 293314 379400
rect 291028 379340 291034 379342
rect 293309 379340 293356 379344
rect 293420 379342 293466 379402
rect 295885 379400 295932 379404
rect 295996 379402 296002 379404
rect 298093 379402 298159 379405
rect 300853 379404 300919 379405
rect 298502 379402 298508 379404
rect 295885 379344 295890 379400
rect 293420 379340 293426 379342
rect 295885 379340 295932 379344
rect 295996 379342 296042 379402
rect 298093 379400 298508 379402
rect 298093 379344 298098 379400
rect 298154 379344 298508 379400
rect 298093 379342 298508 379344
rect 295996 379340 296002 379342
rect 290917 379339 290983 379340
rect 293309 379339 293375 379340
rect 295885 379339 295951 379340
rect 298093 379339 298159 379342
rect 298502 379340 298508 379342
rect 298572 379340 298578 379404
rect 300853 379400 300900 379404
rect 300964 379402 300970 379404
rect 303061 379402 303127 379405
rect 303470 379402 303476 379404
rect 300853 379344 300858 379400
rect 300853 379340 300900 379344
rect 300964 379342 301010 379402
rect 303061 379400 303476 379402
rect 303061 379344 303066 379400
rect 303122 379344 303476 379400
rect 303061 379342 303476 379344
rect 300964 379340 300970 379342
rect 300853 379339 300919 379340
rect 303061 379339 303127 379342
rect 303470 379340 303476 379342
rect 303540 379340 303546 379404
rect 305729 379402 305795 379405
rect 308397 379404 308463 379405
rect 310973 379404 311039 379405
rect 313365 379404 313431 379405
rect 315757 379404 315823 379405
rect 318333 379404 318399 379405
rect 323301 379404 323367 379405
rect 305862 379402 305868 379404
rect 305729 379400 305868 379402
rect 305729 379344 305734 379400
rect 305790 379344 305868 379400
rect 305729 379342 305868 379344
rect 305729 379339 305795 379342
rect 305862 379340 305868 379342
rect 305932 379340 305938 379404
rect 308397 379400 308444 379404
rect 308508 379402 308514 379404
rect 308397 379344 308402 379400
rect 308397 379340 308444 379344
rect 308508 379342 308554 379402
rect 310973 379400 311020 379404
rect 311084 379402 311090 379404
rect 310973 379344 310978 379400
rect 308508 379340 308514 379342
rect 310973 379340 311020 379344
rect 311084 379342 311130 379402
rect 313365 379400 313412 379404
rect 313476 379402 313482 379404
rect 313365 379344 313370 379400
rect 311084 379340 311090 379342
rect 313365 379340 313412 379344
rect 313476 379342 313522 379402
rect 315757 379400 315804 379404
rect 315868 379402 315874 379404
rect 315757 379344 315762 379400
rect 313476 379340 313482 379342
rect 315757 379340 315804 379344
rect 315868 379342 315914 379402
rect 318333 379400 318380 379404
rect 318444 379402 318450 379404
rect 318333 379344 318338 379400
rect 315868 379340 315874 379342
rect 318333 379340 318380 379344
rect 318444 379342 318490 379402
rect 323301 379400 323348 379404
rect 323412 379402 323418 379404
rect 323301 379344 323306 379400
rect 318444 379340 318450 379342
rect 323301 379340 323348 379344
rect 323412 379342 323458 379402
rect 323412 379340 323418 379342
rect 377438 379340 377444 379404
rect 377508 379402 377514 379404
rect 380985 379402 381051 379405
rect 377508 379400 381051 379402
rect 377508 379344 380990 379400
rect 381046 379344 381051 379400
rect 377508 379342 381051 379344
rect 377508 379340 377514 379342
rect 308397 379339 308463 379340
rect 310973 379339 311039 379340
rect 313365 379339 313431 379340
rect 315757 379339 315823 379340
rect 318333 379339 318399 379340
rect 323301 379339 323367 379340
rect 380985 379339 381051 379342
rect 396165 379402 396231 379405
rect 397126 379402 397132 379404
rect 396165 379400 397132 379402
rect 396165 379344 396170 379400
rect 396226 379344 397132 379400
rect 396165 379342 397132 379344
rect 396165 379339 396231 379342
rect 397126 379340 397132 379342
rect 397196 379340 397202 379404
rect 400438 379402 400444 379404
rect 398054 379342 400444 379402
rect 219390 379206 238770 379266
rect 245653 379266 245719 379269
rect 248597 379268 248663 379269
rect 250069 379268 250135 379269
rect 251173 379268 251239 379269
rect 252277 379268 252343 379269
rect 253381 379268 253447 379269
rect 261661 379268 261727 379269
rect 273437 379268 273503 379269
rect 277025 379268 277091 379269
rect 246430 379266 246436 379268
rect 245653 379264 246436 379266
rect 245653 379208 245658 379264
rect 245714 379208 246436 379264
rect 245653 379206 246436 379208
rect 219390 379130 219450 379206
rect 245653 379203 245719 379206
rect 246430 379204 246436 379206
rect 246500 379204 246506 379268
rect 248597 379264 248644 379268
rect 248708 379266 248714 379268
rect 248597 379208 248602 379264
rect 248597 379204 248644 379208
rect 248708 379206 248754 379266
rect 250069 379264 250116 379268
rect 250180 379266 250186 379268
rect 250069 379208 250074 379264
rect 248708 379204 248714 379206
rect 250069 379204 250116 379208
rect 250180 379206 250226 379266
rect 251173 379264 251220 379268
rect 251284 379266 251290 379268
rect 251173 379208 251178 379264
rect 250180 379204 250186 379206
rect 251173 379204 251220 379208
rect 251284 379206 251330 379266
rect 252277 379264 252324 379268
rect 252388 379266 252394 379268
rect 252277 379208 252282 379264
rect 251284 379204 251290 379206
rect 252277 379204 252324 379208
rect 252388 379206 252434 379266
rect 253381 379264 253428 379268
rect 253492 379266 253498 379268
rect 253381 379208 253386 379264
rect 252388 379204 252394 379206
rect 253381 379204 253428 379208
rect 253492 379206 253538 379266
rect 261661 379264 261708 379268
rect 261772 379266 261778 379268
rect 261661 379208 261666 379264
rect 253492 379204 253498 379206
rect 261661 379204 261708 379208
rect 261772 379206 261818 379266
rect 273437 379264 273484 379268
rect 273548 379266 273554 379268
rect 276974 379266 276980 379268
rect 273437 379208 273442 379264
rect 261772 379204 261778 379206
rect 273437 379204 273484 379208
rect 273548 379206 273594 379266
rect 276934 379206 276980 379266
rect 277044 379264 277091 379268
rect 277086 379208 277091 379264
rect 273548 379204 273554 379206
rect 276974 379204 276980 379206
rect 277044 379204 277091 379208
rect 248597 379203 248663 379204
rect 250069 379203 250135 379204
rect 251173 379203 251239 379204
rect 252277 379203 252343 379204
rect 253381 379203 253447 379204
rect 261661 379203 261727 379204
rect 273437 379203 273503 379204
rect 277025 379203 277091 379204
rect 277853 379266 277919 379269
rect 279141 379268 279207 379269
rect 280797 379268 280863 379269
rect 278446 379266 278452 379268
rect 277853 379264 278452 379266
rect 277853 379208 277858 379264
rect 277914 379208 278452 379264
rect 277853 379206 278452 379208
rect 277853 379203 277919 379206
rect 278446 379204 278452 379206
rect 278516 379204 278522 379268
rect 279141 379264 279188 379268
rect 279252 379266 279258 379268
rect 279141 379208 279146 379264
rect 279141 379204 279188 379208
rect 279252 379206 279298 379266
rect 280797 379264 280844 379268
rect 280908 379266 280914 379268
rect 283005 379266 283071 379269
rect 325877 379268 325943 379269
rect 283414 379266 283420 379268
rect 280797 379208 280802 379264
rect 279252 379204 279258 379206
rect 280797 379204 280844 379208
rect 280908 379206 280954 379266
rect 283005 379264 283420 379266
rect 283005 379208 283010 379264
rect 283066 379208 283420 379264
rect 283005 379206 283420 379208
rect 280908 379204 280914 379206
rect 279141 379203 279207 379204
rect 280797 379203 280863 379204
rect 283005 379203 283071 379206
rect 283414 379204 283420 379206
rect 283484 379204 283490 379268
rect 325877 379264 325924 379268
rect 325988 379266 325994 379268
rect 373901 379266 373967 379269
rect 398054 379266 398114 379342
rect 400438 379340 400444 379342
rect 400508 379340 400514 379404
rect 405733 379402 405799 379405
rect 407573 379404 407639 379405
rect 408309 379404 408375 379405
rect 406510 379402 406516 379404
rect 405733 379400 406516 379402
rect 405733 379344 405738 379400
rect 405794 379344 406516 379400
rect 405733 379342 406516 379344
rect 405733 379339 405799 379342
rect 406510 379340 406516 379342
rect 406580 379340 406586 379404
rect 407573 379400 407620 379404
rect 407684 379402 407690 379404
rect 407573 379344 407578 379400
rect 407573 379340 407620 379344
rect 407684 379342 407730 379402
rect 408309 379400 408356 379404
rect 408420 379402 408426 379404
rect 410609 379402 410675 379405
rect 411253 379404 411319 379405
rect 412357 379404 412423 379405
rect 410742 379402 410748 379404
rect 408309 379344 408314 379400
rect 407684 379340 407690 379342
rect 408309 379340 408356 379344
rect 408420 379342 408466 379402
rect 410609 379400 410748 379402
rect 410609 379344 410614 379400
rect 410670 379344 410748 379400
rect 410609 379342 410748 379344
rect 408420 379340 408426 379342
rect 407573 379339 407639 379340
rect 408309 379339 408375 379340
rect 410609 379339 410675 379342
rect 410742 379340 410748 379342
rect 410812 379340 410818 379404
rect 411253 379400 411300 379404
rect 411364 379402 411370 379404
rect 411253 379344 411258 379400
rect 411253 379340 411300 379344
rect 411364 379342 411410 379402
rect 412357 379400 412404 379404
rect 412468 379402 412474 379404
rect 413093 379402 413159 379405
rect 423397 379404 423463 379405
rect 427445 379404 427511 379405
rect 439037 379404 439103 379405
rect 445845 379404 445911 379405
rect 413502 379402 413508 379404
rect 412357 379344 412362 379400
rect 411364 379340 411370 379342
rect 412357 379340 412404 379344
rect 412468 379342 412514 379402
rect 413093 379400 413508 379402
rect 413093 379344 413098 379400
rect 413154 379344 413508 379400
rect 413093 379342 413508 379344
rect 412468 379340 412474 379342
rect 411253 379339 411319 379340
rect 412357 379339 412423 379340
rect 413093 379339 413159 379342
rect 413502 379340 413508 379342
rect 413572 379340 413578 379404
rect 423397 379400 423444 379404
rect 423508 379402 423514 379404
rect 423397 379344 423402 379400
rect 423397 379340 423444 379344
rect 423508 379342 423554 379402
rect 427445 379400 427492 379404
rect 427556 379402 427562 379404
rect 427445 379344 427450 379400
rect 423508 379340 423514 379342
rect 427445 379340 427492 379344
rect 427556 379342 427602 379402
rect 439037 379400 439084 379404
rect 439148 379402 439154 379404
rect 439037 379344 439042 379400
rect 427556 379340 427562 379342
rect 439037 379340 439084 379344
rect 439148 379342 439194 379402
rect 445845 379400 445892 379404
rect 445956 379402 445962 379404
rect 448145 379402 448211 379405
rect 450997 379404 451063 379405
rect 448278 379402 448284 379404
rect 445845 379344 445850 379400
rect 439148 379340 439154 379342
rect 445845 379340 445892 379344
rect 445956 379342 446002 379402
rect 448145 379400 448284 379402
rect 448145 379344 448150 379400
rect 448206 379344 448284 379400
rect 448145 379342 448284 379344
rect 445956 379340 445962 379342
rect 423397 379339 423463 379340
rect 427445 379339 427511 379340
rect 439037 379339 439103 379340
rect 445845 379339 445911 379340
rect 448145 379339 448211 379342
rect 448278 379340 448284 379342
rect 448348 379340 448354 379404
rect 450997 379400 451044 379404
rect 451108 379402 451114 379404
rect 452745 379402 452811 379405
rect 453430 379402 453436 379404
rect 450997 379344 451002 379400
rect 450997 379340 451044 379344
rect 451108 379342 451154 379402
rect 452745 379400 453436 379402
rect 452745 379344 452750 379400
rect 452806 379344 453436 379400
rect 452745 379342 453436 379344
rect 451108 379340 451114 379342
rect 450997 379339 451063 379340
rect 452745 379339 452811 379342
rect 453430 379340 453436 379342
rect 453500 379340 453506 379404
rect 455505 379402 455571 379405
rect 458357 379404 458423 379405
rect 455822 379402 455828 379404
rect 455505 379400 455828 379402
rect 455505 379344 455510 379400
rect 455566 379344 455828 379400
rect 455505 379342 455828 379344
rect 455505 379339 455571 379342
rect 455822 379340 455828 379342
rect 455892 379340 455898 379404
rect 458357 379400 458404 379404
rect 458468 379402 458474 379404
rect 458357 379344 458362 379400
rect 458357 379340 458404 379344
rect 458468 379342 458514 379402
rect 458468 379340 458474 379342
rect 458357 379339 458423 379340
rect 402973 379268 403039 379269
rect 405365 379268 405431 379269
rect 409965 379268 410031 379269
rect 414565 379268 414631 379269
rect 325877 379208 325882 379264
rect 325877 379204 325924 379208
rect 325988 379206 326034 379266
rect 373901 379264 398114 379266
rect 373901 379208 373906 379264
rect 373962 379208 398114 379264
rect 373901 379206 398114 379208
rect 325988 379204 325994 379206
rect 325877 379203 325943 379204
rect 373901 379203 373967 379206
rect 401726 379204 401732 379268
rect 401796 379204 401802 379268
rect 402973 379264 403020 379268
rect 403084 379266 403090 379268
rect 402973 379208 402978 379264
rect 402973 379204 403020 379208
rect 403084 379206 403130 379266
rect 405365 379264 405412 379268
rect 405476 379266 405482 379268
rect 405365 379208 405370 379264
rect 403084 379204 403090 379206
rect 405365 379204 405412 379208
rect 405476 379206 405522 379266
rect 409965 379264 410012 379268
rect 410076 379266 410082 379268
rect 409965 379208 409970 379264
rect 405476 379204 405482 379206
rect 409965 379204 410012 379208
rect 410076 379206 410122 379266
rect 414565 379264 414612 379268
rect 414676 379266 414682 379268
rect 415393 379266 415459 379269
rect 416037 379268 416103 379269
rect 415894 379266 415900 379268
rect 414565 379208 414570 379264
rect 410076 379204 410082 379206
rect 414565 379204 414612 379208
rect 414676 379206 414722 379266
rect 415393 379264 415900 379266
rect 415393 379208 415398 379264
rect 415454 379208 415900 379264
rect 415393 379206 415900 379208
rect 414676 379204 414682 379206
rect 208718 379128 219450 379130
rect 208718 379072 209502 379128
rect 209558 379072 219450 379128
rect 208718 379070 219450 379072
rect 222009 379130 222075 379133
rect 240542 379130 240548 379132
rect 222009 379128 240548 379130
rect 222009 379072 222014 379128
rect 222070 379072 240548 379128
rect 222009 379070 240548 379072
rect 208485 379067 208551 379070
rect 209497 379067 209563 379070
rect 222009 379067 222075 379070
rect 240542 379068 240548 379070
rect 240612 379130 240618 379132
rect 241462 379130 241468 379132
rect 240612 379070 241468 379130
rect 240612 379068 240618 379070
rect 241462 379068 241468 379070
rect 241532 379068 241538 379132
rect 253197 379130 253263 379133
rect 369669 379130 369735 379133
rect 401734 379130 401794 379204
rect 402973 379203 403039 379204
rect 405365 379203 405431 379204
rect 409965 379203 410031 379204
rect 414565 379203 414631 379204
rect 415393 379203 415459 379206
rect 415894 379204 415900 379206
rect 415964 379204 415970 379268
rect 416037 379264 416084 379268
rect 416148 379266 416154 379268
rect 418337 379266 418403 379269
rect 419390 379266 419396 379268
rect 416037 379208 416042 379264
rect 416037 379204 416084 379208
rect 416148 379206 416194 379266
rect 418337 379264 419396 379266
rect 418337 379208 418342 379264
rect 418398 379208 419396 379264
rect 418337 379206 419396 379208
rect 416148 379204 416154 379206
rect 416037 379203 416103 379204
rect 418337 379203 418403 379206
rect 419390 379204 419396 379206
rect 419460 379204 419466 379268
rect 437749 379266 437815 379269
rect 463509 379268 463575 379269
rect 473445 379268 473511 379269
rect 437974 379266 437980 379268
rect 437749 379264 437980 379266
rect 437749 379208 437754 379264
rect 437810 379208 437980 379264
rect 437749 379206 437980 379208
rect 437749 379203 437815 379206
rect 437974 379204 437980 379206
rect 438044 379204 438050 379268
rect 463509 379264 463556 379268
rect 463620 379266 463626 379268
rect 463509 379208 463514 379264
rect 463509 379204 463556 379208
rect 463620 379206 463666 379266
rect 473445 379264 473492 379268
rect 473556 379266 473562 379268
rect 474733 379266 474799 379269
rect 480805 379268 480871 379269
rect 503069 379268 503135 379269
rect 503529 379268 503595 379269
rect 475878 379266 475884 379268
rect 473445 379208 473450 379264
rect 463620 379204 463626 379206
rect 473445 379204 473492 379208
rect 473556 379206 473602 379266
rect 474733 379264 475884 379266
rect 474733 379208 474738 379264
rect 474794 379208 475884 379264
rect 474733 379206 475884 379208
rect 473556 379204 473562 379206
rect 463509 379203 463575 379204
rect 473445 379203 473511 379204
rect 474733 379203 474799 379206
rect 475878 379204 475884 379206
rect 475948 379204 475954 379268
rect 480805 379264 480852 379268
rect 480916 379266 480922 379268
rect 480805 379208 480810 379264
rect 480805 379204 480852 379208
rect 480916 379206 480962 379266
rect 503069 379264 503116 379268
rect 503180 379266 503186 379268
rect 503069 379208 503074 379264
rect 480916 379204 480922 379206
rect 503069 379204 503116 379208
rect 503180 379206 503226 379266
rect 503180 379204 503186 379206
rect 503478 379204 503484 379268
rect 503548 379266 503595 379268
rect 503548 379264 503640 379266
rect 503590 379208 503640 379264
rect 503548 379206 503640 379208
rect 503548 379204 503595 379206
rect 480805 379203 480871 379204
rect 503069 379203 503135 379204
rect 503529 379203 503595 379204
rect 433374 379130 433380 379132
rect 253197 379128 401794 379130
rect 253197 379072 253202 379128
rect 253258 379072 369674 379128
rect 369730 379072 401794 379128
rect 253197 379070 401794 379072
rect 412590 379070 433380 379130
rect 253197 379067 253263 379070
rect 369669 379067 369735 379070
rect 51625 378994 51691 378997
rect 77201 378996 77267 378997
rect 57094 378994 57100 378996
rect 51625 378992 57100 378994
rect 51625 378936 51630 378992
rect 51686 378936 57100 378992
rect 51625 378934 57100 378936
rect 51625 378931 51691 378934
rect 57094 378932 57100 378934
rect 57164 378932 57170 378996
rect 77150 378994 77156 378996
rect 77110 378934 77156 378994
rect 77220 378992 77267 378996
rect 77262 378936 77267 378992
rect 77150 378932 77156 378934
rect 77220 378932 77267 378936
rect 78254 378932 78260 378996
rect 78324 378994 78330 378996
rect 208025 378994 208091 378997
rect 238150 378994 238156 378996
rect 78324 378992 238156 378994
rect 78324 378936 208030 378992
rect 208086 378936 238156 378992
rect 78324 378934 238156 378936
rect 78324 378932 78330 378934
rect 77201 378931 77267 378932
rect 208025 378931 208091 378934
rect 238150 378932 238156 378934
rect 238220 378994 238226 378996
rect 369761 378994 369827 378997
rect 397494 378994 397500 378996
rect 238220 378992 397500 378994
rect 238220 378936 369766 378992
rect 369822 378936 397500 378992
rect 238220 378934 397500 378936
rect 238220 378932 238226 378934
rect 369761 378931 369827 378934
rect 397494 378932 397500 378934
rect 397564 378932 397570 378996
rect 53230 378796 53236 378860
rect 53300 378858 53306 378860
rect 53557 378858 53623 378861
rect 53300 378856 53623 378858
rect 53300 378800 53562 378856
rect 53618 378800 53623 378856
rect 53300 378798 53623 378800
rect 53300 378796 53306 378798
rect 53557 378795 53623 378798
rect 81433 378858 81499 378861
rect 81934 378858 81940 378860
rect 81433 378856 81940 378858
rect 81433 378800 81438 378856
rect 81494 378800 81940 378856
rect 81433 378798 81940 378800
rect 81433 378795 81499 378798
rect 81934 378796 81940 378798
rect 82004 378858 82010 378860
rect 221641 378858 221707 378861
rect 82004 378856 221707 378858
rect 82004 378800 221646 378856
rect 221702 378800 221707 378856
rect 82004 378798 221707 378800
rect 82004 378796 82010 378798
rect 221641 378795 221707 378798
rect 241462 378796 241468 378860
rect 241532 378858 241538 378860
rect 373625 378858 373691 378861
rect 373901 378858 373967 378861
rect 241532 378856 373967 378858
rect 241532 378800 373630 378856
rect 373686 378800 373906 378856
rect 373962 378800 373967 378856
rect 241532 378798 373967 378800
rect 241532 378796 241538 378798
rect 373625 378795 373691 378798
rect 373901 378795 373967 378798
rect 380985 378858 381051 378861
rect 381169 378858 381235 378861
rect 412590 378858 412650 379070
rect 433374 379068 433380 379070
rect 433444 379068 433450 379132
rect 380985 378856 412650 378858
rect 380985 378800 380990 378856
rect 381046 378800 381174 378856
rect 381230 378800 412650 378856
rect 380985 378798 412650 378800
rect 418245 378858 418311 378861
rect 418470 378858 418476 378860
rect 418245 378856 418476 378858
rect 418245 378800 418250 378856
rect 418306 378800 418476 378856
rect 418245 378798 418476 378800
rect 380985 378795 381051 378798
rect 381169 378795 381235 378798
rect 418245 378795 418311 378798
rect 418470 378796 418476 378798
rect 418540 378796 418546 378860
rect 467925 378858 467991 378861
rect 470869 378860 470935 378861
rect 468518 378858 468524 378860
rect 467925 378856 468524 378858
rect 467925 378800 467930 378856
rect 467986 378800 468524 378856
rect 467925 378798 468524 378800
rect 467925 378795 467991 378798
rect 468518 378796 468524 378798
rect 468588 378796 468594 378860
rect 470869 378856 470916 378860
rect 470980 378858 470986 378860
rect 477585 378858 477651 378861
rect 483381 378860 483447 378861
rect 478454 378858 478460 378860
rect 470869 378800 470874 378856
rect 470869 378796 470916 378800
rect 470980 378798 471026 378858
rect 477585 378856 478460 378858
rect 477585 378800 477590 378856
rect 477646 378800 478460 378856
rect 477585 378798 478460 378800
rect 470980 378796 470986 378798
rect 470869 378795 470935 378796
rect 477585 378795 477651 378798
rect 478454 378796 478460 378798
rect 478524 378796 478530 378860
rect 483381 378856 483428 378860
rect 483492 378858 483498 378860
rect 483381 378800 483386 378856
rect 483381 378796 483428 378800
rect 483492 378798 483538 378858
rect 483492 378796 483498 378798
rect 483381 378795 483447 378796
rect 80329 378722 80395 378725
rect 220997 378722 221063 378725
rect 222009 378722 222075 378725
rect 80329 378720 222075 378722
rect 80329 378664 80334 378720
rect 80390 378664 221002 378720
rect 221058 378664 222014 378720
rect 222070 378664 222075 378720
rect 80329 378662 222075 378664
rect 80329 378659 80395 378662
rect 220997 378659 221063 378662
rect 222009 378659 222075 378662
rect 233877 378722 233943 378725
rect 239254 378722 239260 378724
rect 233877 378720 239260 378722
rect 233877 378664 233882 378720
rect 233938 378664 239260 378720
rect 233877 378662 239260 378664
rect 233877 378659 233943 378662
rect 239254 378660 239260 378662
rect 239324 378722 239330 378724
rect 239324 378662 369870 378722
rect 239324 378660 239330 378662
rect 94681 378588 94747 378589
rect 94630 378586 94636 378588
rect 94590 378526 94636 378586
rect 94700 378584 94747 378588
rect 94742 378528 94747 378584
rect 94630 378524 94636 378526
rect 94700 378524 94747 378528
rect 97022 378524 97028 378588
rect 97092 378586 97098 378588
rect 97717 378586 97783 378589
rect 97092 378584 97783 378586
rect 97092 378528 97722 378584
rect 97778 378528 97783 378584
rect 97092 378526 97783 378528
rect 97092 378524 97098 378526
rect 94681 378523 94747 378524
rect 97717 378523 97783 378526
rect 117078 378524 117084 378588
rect 117148 378586 117154 378588
rect 204805 378586 204871 378589
rect 117148 378584 204871 378586
rect 117148 378528 204810 378584
rect 204866 378528 204871 378584
rect 117148 378526 204871 378528
rect 117148 378524 117154 378526
rect 204805 378523 204871 378526
rect 209998 378524 210004 378588
rect 210068 378586 210074 378588
rect 211061 378586 211127 378589
rect 210068 378584 211127 378586
rect 210068 378528 211066 378584
rect 211122 378528 211127 378584
rect 210068 378526 211127 378528
rect 210068 378524 210074 378526
rect 211061 378523 211127 378526
rect 212441 378586 212507 378589
rect 221273 378586 221339 378589
rect 320909 378588 320975 378589
rect 278078 378586 278084 378588
rect 212441 378584 278084 378586
rect 212441 378528 212446 378584
rect 212502 378528 221278 378584
rect 221334 378528 278084 378584
rect 212441 378526 278084 378528
rect 212441 378523 212507 378526
rect 221273 378523 221339 378526
rect 278078 378524 278084 378526
rect 278148 378524 278154 378588
rect 320909 378584 320956 378588
rect 321020 378586 321026 378588
rect 320909 378528 320914 378584
rect 320909 378524 320956 378528
rect 321020 378526 321066 378586
rect 321020 378524 321026 378526
rect 320909 378523 320975 378524
rect 100753 378452 100819 378453
rect 104065 378452 104131 378453
rect 125961 378452 126027 378453
rect 100702 378450 100708 378452
rect 100662 378390 100708 378450
rect 100772 378448 100819 378452
rect 104014 378450 104020 378452
rect 100814 378392 100819 378448
rect 100702 378388 100708 378390
rect 100772 378388 100819 378392
rect 103974 378390 104020 378450
rect 104084 378448 104131 378452
rect 125910 378450 125916 378452
rect 104126 378392 104131 378448
rect 104014 378388 104020 378390
rect 104084 378388 104131 378392
rect 125870 378390 125916 378450
rect 125980 378448 126027 378452
rect 126022 378392 126027 378448
rect 125910 378388 125916 378390
rect 125980 378388 126027 378392
rect 100753 378387 100819 378388
rect 104065 378387 104131 378388
rect 125961 378387 126027 378388
rect 131021 378452 131087 378453
rect 131021 378448 131068 378452
rect 131132 378450 131138 378452
rect 131021 378392 131026 378448
rect 131021 378388 131068 378392
rect 131132 378390 131178 378450
rect 131132 378388 131138 378390
rect 183134 378388 183140 378452
rect 183204 378450 183210 378452
rect 183461 378450 183527 378453
rect 183204 378448 183527 378450
rect 183204 378392 183466 378448
rect 183522 378392 183527 378448
rect 183204 378390 183527 378392
rect 183204 378388 183210 378390
rect 131021 378387 131087 378388
rect 183461 378387 183527 378390
rect 208485 378450 208551 378453
rect 209405 378450 209471 378453
rect 233877 378450 233943 378453
rect 208485 378448 233943 378450
rect 208485 378392 208490 378448
rect 208546 378392 209410 378448
rect 209466 378392 233882 378448
rect 233938 378392 233943 378448
rect 208485 378390 233943 378392
rect 208485 378387 208551 378390
rect 209405 378387 209471 378390
rect 233877 378387 233943 378390
rect 248229 378452 248295 378453
rect 250621 378452 250687 378453
rect 253565 378452 253631 378453
rect 255957 378452 256023 378453
rect 258349 378452 258415 378453
rect 260925 378452 260991 378453
rect 263593 378452 263659 378453
rect 248229 378448 248276 378452
rect 248340 378450 248346 378452
rect 248229 378392 248234 378448
rect 248229 378388 248276 378392
rect 248340 378390 248386 378450
rect 250621 378448 250668 378452
rect 250732 378450 250738 378452
rect 250621 378392 250626 378448
rect 248340 378388 248346 378390
rect 250621 378388 250668 378392
rect 250732 378390 250778 378450
rect 253565 378448 253612 378452
rect 253676 378450 253682 378452
rect 253565 378392 253570 378448
rect 250732 378388 250738 378390
rect 253565 378388 253612 378392
rect 253676 378390 253722 378450
rect 255957 378448 256004 378452
rect 256068 378450 256074 378452
rect 255957 378392 255962 378448
rect 253676 378388 253682 378390
rect 255957 378388 256004 378392
rect 256068 378390 256114 378450
rect 258349 378448 258396 378452
rect 258460 378450 258466 378452
rect 258349 378392 258354 378448
rect 256068 378388 256074 378390
rect 258349 378388 258396 378392
rect 258460 378390 258506 378450
rect 260925 378448 260972 378452
rect 261036 378450 261042 378452
rect 263542 378450 263548 378452
rect 260925 378392 260930 378448
rect 258460 378388 258466 378390
rect 260925 378388 260972 378392
rect 261036 378390 261082 378450
rect 263502 378390 263548 378450
rect 263612 378448 263659 378452
rect 263654 378392 263659 378448
rect 261036 378388 261042 378390
rect 263542 378388 263548 378390
rect 263612 378388 263659 378392
rect 248229 378387 248295 378388
rect 250621 378387 250687 378388
rect 253565 378387 253631 378388
rect 255957 378387 256023 378388
rect 258349 378387 258415 378388
rect 260925 378387 260991 378388
rect 263593 378387 263659 378388
rect 265341 378450 265407 378453
rect 265934 378450 265940 378452
rect 265341 378448 265940 378450
rect 265341 378392 265346 378448
rect 265402 378392 265940 378448
rect 265341 378390 265940 378392
rect 265341 378387 265407 378390
rect 265934 378388 265940 378390
rect 266004 378388 266010 378452
rect 268101 378450 268167 378453
rect 343173 378452 343239 378453
rect 268326 378450 268332 378452
rect 268101 378448 268332 378450
rect 268101 378392 268106 378448
rect 268162 378392 268332 378448
rect 268101 378390 268332 378392
rect 268101 378387 268167 378390
rect 268326 378388 268332 378390
rect 268396 378388 268402 378452
rect 343173 378448 343220 378452
rect 343284 378450 343290 378452
rect 369810 378450 369870 378662
rect 377622 378660 377628 378724
rect 377692 378722 377698 378724
rect 435766 378722 435772 378724
rect 377692 378662 435772 378722
rect 377692 378660 377698 378662
rect 381126 378589 381186 378662
rect 435766 378660 435772 378662
rect 435836 378660 435842 378724
rect 381077 378584 381186 378589
rect 396073 378588 396139 378589
rect 396022 378586 396028 378588
rect 381077 378528 381082 378584
rect 381138 378528 381186 378584
rect 381077 378526 381186 378528
rect 395982 378526 396028 378586
rect 396092 378584 396139 378588
rect 396134 378528 396139 378584
rect 381077 378523 381143 378526
rect 396022 378524 396028 378526
rect 396092 378524 396139 378528
rect 396073 378523 396139 378524
rect 403617 378586 403683 378589
rect 428181 378588 428247 378589
rect 404118 378586 404124 378588
rect 403617 378584 404124 378586
rect 403617 378528 403622 378584
rect 403678 378528 404124 378584
rect 403617 378526 404124 378528
rect 403617 378523 403683 378526
rect 404118 378524 404124 378526
rect 404188 378524 404194 378588
rect 428181 378584 428228 378588
rect 428292 378586 428298 378588
rect 430665 378586 430731 378589
rect 430982 378586 430988 378588
rect 428181 378528 428186 378584
rect 428181 378524 428228 378528
rect 428292 378526 428338 378586
rect 430665 378584 430988 378586
rect 430665 378528 430670 378584
rect 430726 378528 430988 378584
rect 430665 378526 430988 378528
rect 428292 378524 428298 378526
rect 428181 378523 428247 378524
rect 430665 378523 430731 378526
rect 430982 378524 430988 378526
rect 431052 378524 431058 378588
rect 372521 378450 372587 378453
rect 399518 378450 399524 378452
rect 343173 378392 343178 378448
rect 343173 378388 343220 378392
rect 343284 378390 343330 378450
rect 369810 378448 399524 378450
rect 369810 378392 372526 378448
rect 372582 378392 399524 378448
rect 369810 378390 399524 378392
rect 343284 378388 343290 378390
rect 343173 378387 343239 378388
rect 372521 378387 372587 378390
rect 399518 378388 399524 378390
rect 399588 378388 399594 378452
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 101806 378252 101812 378316
rect 101876 378314 101882 378316
rect 101949 378314 102015 378317
rect 101876 378312 102015 378314
rect 101876 378256 101954 378312
rect 102010 378256 102015 378312
rect 101876 378254 102015 378256
rect 101876 378252 101882 378254
rect 101949 378251 102015 378254
rect 118182 378252 118188 378316
rect 118252 378314 118258 378316
rect 212441 378314 212507 378317
rect 118252 378312 212507 378314
rect 118252 378256 212446 378312
rect 212502 378256 212507 378312
rect 118252 378254 212507 378256
rect 118252 378252 118258 378254
rect 212441 378251 212507 378254
rect 221181 378314 221247 378317
rect 221641 378314 221707 378317
rect 241830 378314 241836 378316
rect 221181 378312 241836 378314
rect 221181 378256 221186 378312
rect 221242 378256 221646 378312
rect 221702 378256 241836 378312
rect 221181 378254 241836 378256
rect 221181 378251 221247 378254
rect 221641 378251 221707 378254
rect 241830 378252 241836 378254
rect 241900 378314 241906 378316
rect 253197 378314 253263 378317
rect 241900 378312 253263 378314
rect 241900 378256 253202 378312
rect 253258 378256 253263 378312
rect 241900 378254 253263 378256
rect 241900 378252 241906 378254
rect 253197 378251 253263 378254
rect 262765 378316 262831 378317
rect 266353 378316 266419 378317
rect 262765 378312 262812 378316
rect 262876 378314 262882 378316
rect 266302 378314 266308 378316
rect 262765 378256 262770 378312
rect 262765 378252 262812 378256
rect 262876 378254 262922 378314
rect 266262 378254 266308 378314
rect 266372 378312 266419 378316
rect 266414 378256 266419 378312
rect 262876 378252 262882 378254
rect 266302 378252 266308 378254
rect 266372 378252 266419 378256
rect 262765 378251 262831 378252
rect 266353 378251 266419 378252
rect 267549 378316 267615 378317
rect 267549 378312 267596 378316
rect 267660 378314 267666 378316
rect 267549 378256 267554 378312
rect 267549 378252 267596 378256
rect 267660 378254 267706 378314
rect 267660 378252 267666 378254
rect 343398 378252 343404 378316
rect 343468 378314 343474 378316
rect 343541 378314 343607 378317
rect 343468 378312 343607 378314
rect 343468 378256 343546 378312
rect 343602 378256 343607 378312
rect 343468 378254 343607 378256
rect 343468 378252 343474 378254
rect 267549 378251 267615 378252
rect 343541 378251 343607 378254
rect 428273 378314 428339 378317
rect 428590 378314 428596 378316
rect 428273 378312 428596 378314
rect 428273 378256 428278 378312
rect 428334 378256 428596 378312
rect 428273 378254 428596 378256
rect 428273 378251 428339 378254
rect 428590 378252 428596 378254
rect 428660 378252 428666 378316
rect 583520 378300 584960 378390
rect 106457 378180 106523 378181
rect 107561 378180 107627 378181
rect 106406 378178 106412 378180
rect 106366 378118 106412 378178
rect 106476 378176 106523 378180
rect 107510 378178 107516 378180
rect 106518 378120 106523 378176
rect 106406 378116 106412 378118
rect 106476 378116 106523 378120
rect 107470 378118 107516 378178
rect 107580 378176 107627 378180
rect 107622 378120 107627 378176
rect 107510 378116 107516 378118
rect 107580 378116 107627 378120
rect 106457 378115 106523 378116
rect 107561 378115 107627 378116
rect 182265 378178 182331 378181
rect 182817 378178 182883 378181
rect 183502 378178 183508 378180
rect 182265 378176 183508 378178
rect 182265 378120 182270 378176
rect 182326 378120 182822 378176
rect 182878 378120 183508 378176
rect 182265 378118 183508 378120
rect 182265 378115 182331 378118
rect 182817 378115 182883 378118
rect 183502 378116 183508 378118
rect 183572 378116 183578 378180
rect 204805 378178 204871 378181
rect 205449 378178 205515 378181
rect 276013 378178 276079 378181
rect 204805 378176 276079 378178
rect 204805 378120 204810 378176
rect 204866 378120 205454 378176
rect 205510 378120 276018 378176
rect 276074 378120 276079 378176
rect 204805 378118 276079 378120
rect 204805 378115 204871 378118
rect 205449 378115 205515 378118
rect 276013 378115 276079 378118
rect 376937 378178 377003 378181
rect 416957 378180 417023 378181
rect 418153 378180 418219 378181
rect 377990 378178 377996 378180
rect 376937 378176 377996 378178
rect 376937 378120 376942 378176
rect 376998 378120 377996 378176
rect 376937 378118 377996 378120
rect 376937 378115 377003 378118
rect 377990 378116 377996 378118
rect 378060 378116 378066 378180
rect 416957 378176 417004 378180
rect 417068 378178 417074 378180
rect 418102 378178 418108 378180
rect 416957 378120 416962 378176
rect 416957 378116 417004 378120
rect 417068 378118 417114 378178
rect 418062 378118 418108 378178
rect 418172 378176 418219 378180
rect 418214 378120 418219 378176
rect 417068 378116 417074 378118
rect 418102 378116 418108 378118
rect 418172 378116 418219 378120
rect 416957 378115 417023 378116
rect 418153 378115 418219 378116
rect 419809 378178 419875 378181
rect 423949 378180 424015 378181
rect 426433 378180 426499 378181
rect 420678 378178 420684 378180
rect 419809 378176 420684 378178
rect 419809 378120 419814 378176
rect 419870 378120 420684 378176
rect 419809 378118 420684 378120
rect 419809 378115 419875 378118
rect 420678 378116 420684 378118
rect 420748 378116 420754 378180
rect 423949 378176 423996 378180
rect 424060 378178 424066 378180
rect 426382 378178 426388 378180
rect 423949 378120 423954 378176
rect 423949 378116 423996 378120
rect 424060 378118 424106 378178
rect 426342 378118 426388 378178
rect 426452 378176 426499 378180
rect 426494 378120 426499 378176
rect 424060 378116 424066 378118
rect 426382 378116 426388 378118
rect 426452 378116 426499 378120
rect 423949 378115 424015 378116
rect 426433 378115 426499 378116
rect 429377 378178 429443 378181
rect 431125 378180 431191 378181
rect 432229 378180 432295 378181
rect 429694 378178 429700 378180
rect 429377 378176 429700 378178
rect 429377 378120 429382 378176
rect 429438 378120 429700 378176
rect 429377 378118 429700 378120
rect 429377 378115 429443 378118
rect 429694 378116 429700 378118
rect 429764 378116 429770 378180
rect 431125 378176 431172 378180
rect 431236 378178 431242 378180
rect 431125 378120 431130 378176
rect 431125 378116 431172 378120
rect 431236 378118 431282 378178
rect 432229 378176 432276 378180
rect 432340 378178 432346 378180
rect 432229 378120 432234 378176
rect 431236 378116 431242 378118
rect 432229 378116 432276 378120
rect 432340 378118 432386 378178
rect 432340 378116 432346 378118
rect 460974 378116 460980 378180
rect 461044 378116 461050 378180
rect 431125 378115 431191 378116
rect 432229 378115 432295 378116
rect 198733 378042 198799 378045
rect 273253 378042 273319 378045
rect 198733 378040 273319 378042
rect 198733 377984 198738 378040
rect 198794 377984 273258 378040
rect 273314 377984 273319 378040
rect 198733 377982 273319 377984
rect 198733 377979 198799 377982
rect 273253 377979 273319 377982
rect 359774 377980 359780 378044
rect 359844 378042 359850 378044
rect 460982 378042 461042 378116
rect 359844 377982 461042 378042
rect 359844 377980 359850 377982
rect 95969 377906 96035 377909
rect 211429 377906 211495 377909
rect 95969 377904 211495 377906
rect 95969 377848 95974 377904
rect 96030 377848 211434 377904
rect 211490 377848 211495 377904
rect 95969 377846 211495 377848
rect 95969 377843 96035 377846
rect 211429 377843 211495 377846
rect 211838 377844 211844 377908
rect 211908 377906 211914 377908
rect 212441 377906 212507 377909
rect 211908 377904 212507 377906
rect 211908 377848 212446 377904
rect 212502 377848 212507 377904
rect 211908 377846 212507 377848
rect 211908 377844 211914 377846
rect 212441 377843 212507 377846
rect 212574 377844 212580 377908
rect 212644 377906 212650 377908
rect 213821 377906 213887 377909
rect 212644 377904 213887 377906
rect 212644 377848 213826 377904
rect 213882 377848 213887 377904
rect 212644 377846 213887 377848
rect 212644 377844 212650 377846
rect 213821 377843 213887 377846
rect 215334 377844 215340 377908
rect 215404 377906 215410 377908
rect 215569 377906 215635 377909
rect 215404 377904 215635 377906
rect 215404 377848 215574 377904
rect 215630 377848 215635 377904
rect 215404 377846 215635 377848
rect 215404 377844 215410 377846
rect 215569 377843 215635 377846
rect 105353 377770 105419 377773
rect 215661 377770 215727 377773
rect 221365 377770 221431 377773
rect 221825 377770 221891 377773
rect 105353 377768 221891 377770
rect 105353 377712 105358 377768
rect 105414 377712 215666 377768
rect 215722 377712 221370 377768
rect 221426 377712 221830 377768
rect 221886 377712 221891 377768
rect 105353 377710 221891 377712
rect 105353 377707 105419 377710
rect 215661 377707 215727 377710
rect 221365 377707 221431 377710
rect 221825 377707 221891 377710
rect 98361 377634 98427 377637
rect 207933 377634 207999 377637
rect 98361 377632 207999 377634
rect 98361 377576 98366 377632
rect 98422 377576 207938 377632
rect 207994 377576 207999 377632
rect 98361 377574 207999 377576
rect 98361 377571 98427 377574
rect 207933 377571 207999 377574
rect 211429 377634 211495 377637
rect 212717 377634 212783 377637
rect 213269 377634 213335 377637
rect 211429 377632 213335 377634
rect 211429 377576 211434 377632
rect 211490 377576 212722 377632
rect 212778 377576 213274 377632
rect 213330 377576 213335 377632
rect 211429 377574 213335 377576
rect 211429 377571 211495 377574
rect 212717 377571 212783 377574
rect 213269 377571 213335 377574
rect 43437 377498 43503 377501
rect 199469 377498 199535 377501
rect 43437 377496 199535 377498
rect 43437 377440 43442 377496
rect 43498 377440 199474 377496
rect 199530 377440 199535 377496
rect 43437 377438 199535 377440
rect 43437 377435 43503 377438
rect 199469 377435 199535 377438
rect 211654 376620 211660 376684
rect 211724 376682 211730 376684
rect 212349 376682 212415 376685
rect 211724 376680 212415 376682
rect 211724 376624 212354 376680
rect 212410 376624 212415 376680
rect 211724 376622 212415 376624
rect 211724 376620 211730 376622
rect 212349 376619 212415 376622
rect 213862 376620 213868 376684
rect 213932 376682 213938 376684
rect 215201 376682 215267 376685
rect 213932 376680 215267 376682
rect 213932 376624 215206 376680
rect 215262 376624 215267 376680
rect 213932 376622 215267 376624
rect 213932 376620 213938 376622
rect 215201 376619 215267 376622
rect 216489 376682 216555 376685
rect 216622 376682 216628 376684
rect 216489 376680 216628 376682
rect 216489 376624 216494 376680
rect 216550 376624 216628 376680
rect 216489 376622 216628 376624
rect 216489 376619 216555 376622
rect 216622 376620 216628 376622
rect 216692 376620 216698 376684
rect 377254 376620 377260 376684
rect 377324 376682 377330 376684
rect 480805 376682 480871 376685
rect 377324 376680 480871 376682
rect 377324 376624 480810 376680
rect 480866 376624 480871 376680
rect 377324 376622 480871 376624
rect 377324 376620 377330 376622
rect 480805 376619 480871 376622
rect 217542 375260 217548 375324
rect 217612 375322 217618 375324
rect 325877 375322 325943 375325
rect 217612 375320 325943 375322
rect 217612 375264 325882 375320
rect 325938 375264 325943 375320
rect 217612 375262 325943 375264
rect 217612 375260 217618 375262
rect 325877 375259 325943 375262
rect 217501 375052 217567 375053
rect 217501 375048 217548 375052
rect 217612 375050 217618 375052
rect 217501 374992 217506 375048
rect 217501 374988 217548 374992
rect 217612 374990 217658 375050
rect 217612 374988 217618 374990
rect 217501 374987 217567 374988
rect 359958 374580 359964 374644
rect 360028 374642 360034 374644
rect 371785 374642 371851 374645
rect 419809 374642 419875 374645
rect 360028 374640 419875 374642
rect 360028 374584 371790 374640
rect 371846 374584 419814 374640
rect 419870 374584 419875 374640
rect 360028 374582 419875 374584
rect 360028 374580 360034 374582
rect 371785 374579 371851 374582
rect 419809 374579 419875 374582
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect 178585 358868 178651 358869
rect 179689 358868 179755 358869
rect 190913 358868 190979 358869
rect 338481 358868 338547 358869
rect 178534 358866 178540 358868
rect 178494 358806 178540 358866
rect 178604 358864 178651 358868
rect 179638 358866 179644 358868
rect 178646 358808 178651 358864
rect 178534 358804 178540 358806
rect 178604 358804 178651 358808
rect 179598 358806 179644 358866
rect 179708 358864 179755 358868
rect 190862 358866 190868 358868
rect 179750 358808 179755 358864
rect 179638 358804 179644 358806
rect 179708 358804 179755 358808
rect 190822 358806 190868 358866
rect 190932 358864 190979 358868
rect 338430 358866 338436 358868
rect 190974 358808 190979 358864
rect 190862 358804 190868 358806
rect 190932 358804 190979 358808
rect 338390 358806 338436 358866
rect 338500 358864 338547 358868
rect 338542 358808 338547 358864
rect 338430 358804 338436 358806
rect 338500 358804 338547 358808
rect 339718 358804 339724 358868
rect 339788 358866 339794 358868
rect 339861 358866 339927 358869
rect 339788 358864 339927 358866
rect 339788 358808 339866 358864
rect 339922 358808 339927 358864
rect 339788 358806 339927 358808
rect 339788 358804 339794 358806
rect 178585 358803 178651 358804
rect 179689 358803 179755 358804
rect 190913 358803 190979 358804
rect 338481 358803 338547 358804
rect 339861 358803 339927 358806
rect 350942 358804 350948 358868
rect 351012 358866 351018 358868
rect 351729 358866 351795 358869
rect 351012 358864 351795 358866
rect 351012 358808 351734 358864
rect 351790 358808 351795 358864
rect 351012 358806 351795 358808
rect 351012 358804 351018 358806
rect 351729 358803 351795 358806
rect 498510 358804 498516 358868
rect 498580 358866 498586 358868
rect 498929 358866 498995 358869
rect 498580 358864 498995 358866
rect 498580 358808 498934 358864
rect 498990 358808 498995 358864
rect 498580 358806 498995 358808
rect 498580 358804 498586 358806
rect 498929 358803 498995 358806
rect 499798 358804 499804 358868
rect 499868 358866 499874 358868
rect 500769 358866 500835 358869
rect 510889 358868 510955 358869
rect 510838 358866 510844 358868
rect 499868 358864 500835 358866
rect 499868 358808 500774 358864
rect 500830 358808 500835 358864
rect 499868 358806 500835 358808
rect 510798 358806 510844 358866
rect 510908 358864 510955 358868
rect 510950 358808 510955 358864
rect 499868 358804 499874 358806
rect 500769 358803 500835 358806
rect 510838 358804 510844 358806
rect 510908 358804 510955 358808
rect 510889 358803 510955 358804
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 196558 353154 196618 353190
rect 198825 353154 198891 353157
rect 196558 353152 198891 353154
rect 196558 353096 198830 353152
rect 198886 353096 198891 353152
rect 196558 353094 198891 353096
rect 356562 353154 356622 353190
rect 358905 353154 358971 353157
rect 356562 353152 358971 353154
rect 356562 353096 358910 353152
rect 358966 353096 358971 353152
rect 356562 353094 358971 353096
rect 198825 353091 198891 353094
rect 358905 353091 358971 353094
rect 516558 352882 516618 353190
rect 519261 352882 519327 352885
rect 519537 352882 519603 352885
rect 516558 352880 519603 352882
rect 516558 352824 519266 352880
rect 519322 352824 519542 352880
rect 519598 352824 519603 352880
rect 516558 352822 519603 352824
rect 519261 352819 519327 352822
rect 519537 352819 519603 352822
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 57513 311130 57579 311133
rect 57513 311128 60062 311130
rect 57513 311072 57518 311128
rect 57574 311072 60062 311128
rect 57513 311070 60062 311072
rect 57513 311067 57579 311070
rect 60002 310894 60062 311070
rect 217317 310994 217383 310997
rect 217501 310994 217567 310997
rect 217317 310992 219450 310994
rect 217317 310936 217322 310992
rect 217378 310936 217506 310992
rect 217562 310936 219450 310992
rect 217317 310934 219450 310936
rect 217317 310931 217383 310934
rect 217501 310931 217567 310934
rect 219390 310924 219450 310934
rect 219390 310864 220064 310924
rect 379838 310864 380052 310924
rect 376937 310858 377003 310861
rect 377581 310858 377647 310861
rect 379838 310858 379898 310864
rect 376937 310856 379898 310858
rect 376937 310800 376942 310856
rect 376998 310800 377586 310856
rect 377642 310800 379898 310856
rect 376937 310798 379898 310800
rect 376937 310795 377003 310798
rect 377581 310795 377647 310798
rect 377213 310042 377279 310045
rect 377857 310042 377923 310045
rect 377213 310040 379898 310042
rect 377213 309984 377218 310040
rect 377274 309984 377862 310040
rect 377918 309984 379898 310040
rect 377213 309982 379898 309984
rect 377213 309979 377279 309982
rect 377857 309979 377923 309982
rect 379838 309972 379898 309982
rect 56869 309906 56935 309909
rect 60002 309906 60062 309942
rect 219390 309912 220064 309972
rect 379838 309912 380052 309972
rect 56869 309904 60062 309906
rect 56869 309848 56874 309904
rect 56930 309848 60062 309904
rect 56869 309846 60062 309848
rect 216949 309906 217015 309909
rect 217961 309906 218027 309909
rect 219390 309906 219450 309912
rect 216949 309904 219450 309906
rect 216949 309848 216954 309904
rect 217010 309848 217966 309904
rect 218022 309848 219450 309904
rect 216949 309846 219450 309848
rect 56869 309843 56935 309846
rect 216949 309843 217015 309846
rect 217961 309843 218027 309846
rect 216673 309090 216739 309093
rect 217685 309090 217751 309093
rect 216673 309088 217751 309090
rect 216673 309032 216678 309088
rect 216734 309032 217690 309088
rect 217746 309032 217751 309088
rect 216673 309030 217751 309032
rect 216673 309027 216739 309030
rect 217685 309027 217751 309030
rect 57789 307866 57855 307869
rect 217685 307866 217751 307869
rect 377673 307866 377739 307869
rect 57789 307864 59922 307866
rect 57789 307808 57794 307864
rect 57850 307808 59922 307864
rect 57789 307806 59922 307808
rect 57789 307803 57855 307806
rect 59862 307796 59922 307806
rect 217685 307864 219450 307866
rect 217685 307808 217690 307864
rect 217746 307808 219450 307864
rect 217685 307806 219450 307808
rect 217685 307803 217751 307806
rect 219390 307796 219450 307806
rect 377673 307864 379898 307866
rect 377673 307808 377678 307864
rect 377734 307808 379898 307864
rect 377673 307806 379898 307808
rect 377673 307803 377739 307806
rect 379838 307796 379898 307806
rect 59862 307736 60032 307796
rect 219390 307736 220064 307796
rect 379838 307736 380052 307796
rect 216857 307730 216923 307733
rect 217409 307730 217475 307733
rect 216857 307728 217475 307730
rect 216857 307672 216862 307728
rect 216918 307672 217414 307728
rect 217470 307672 217475 307728
rect 216857 307670 217475 307672
rect 216857 307667 216923 307670
rect 217409 307667 217475 307670
rect 57697 306778 57763 306781
rect 60002 306778 60062 306814
rect 219390 306784 220064 306844
rect 379838 306784 380052 306844
rect 57697 306776 60062 306778
rect 57697 306720 57702 306776
rect 57758 306720 60062 306776
rect 57697 306718 60062 306720
rect 217409 306778 217475 306781
rect 219390 306778 219450 306784
rect 217409 306776 219450 306778
rect 217409 306720 217414 306776
rect 217470 306720 219450 306776
rect 217409 306718 219450 306720
rect 377949 306778 378015 306781
rect 379838 306778 379898 306784
rect 377949 306776 379898 306778
rect 377949 306720 377954 306776
rect 378010 306720 379898 306776
rect 377949 306718 379898 306720
rect 57697 306715 57763 306718
rect 217409 306715 217475 306718
rect 377949 306715 378015 306718
rect -960 306234 480 306324
rect -960 306174 674 306234
rect -960 306098 480 306174
rect 614 306098 674 306174
rect -960 306084 674 306098
rect 246 306038 674 306084
rect 246 305554 306 306038
rect 246 305494 6930 305554
rect 6870 305010 6930 305494
rect 54334 305010 54340 305012
rect 6870 304950 54340 305010
rect 54334 304948 54340 304950
rect 54404 304948 54410 305012
rect 57605 305010 57671 305013
rect 57789 305010 57855 305013
rect 60002 305010 60062 305046
rect 219390 305016 220064 305076
rect 379838 305016 380052 305076
rect 57605 305008 60062 305010
rect 57605 304952 57610 305008
rect 57666 304952 57794 305008
rect 57850 304952 60062 305008
rect 57605 304950 60062 304952
rect 217777 305010 217843 305013
rect 219390 305010 219450 305016
rect 217777 305008 219450 305010
rect 217777 304952 217782 305008
rect 217838 304952 219450 305008
rect 217777 304950 219450 304952
rect 377581 305010 377647 305013
rect 379838 305010 379898 305016
rect 377581 305008 379898 305010
rect 377581 304952 377586 305008
rect 377642 304952 379898 305008
rect 377581 304950 379898 304952
rect 57605 304947 57671 304950
rect 57789 304947 57855 304950
rect 217777 304947 217843 304950
rect 377581 304947 377647 304950
rect 57605 303650 57671 303653
rect 60002 303650 60062 303958
rect 219390 303928 220064 303988
rect 379838 303928 380052 303988
rect 217593 303922 217659 303925
rect 219390 303922 219450 303928
rect 217593 303920 219450 303922
rect 217593 303864 217598 303920
rect 217654 303864 219450 303920
rect 217593 303862 219450 303864
rect 377857 303922 377923 303925
rect 379838 303922 379898 303928
rect 377857 303920 379898 303922
rect 377857 303864 377862 303920
rect 377918 303864 379898 303920
rect 377857 303862 379898 303864
rect 217593 303859 217659 303862
rect 377857 303859 377923 303862
rect 57605 303648 60062 303650
rect 57605 303592 57610 303648
rect 57666 303592 60062 303648
rect 57605 303590 60062 303592
rect 57605 303587 57671 303590
rect 57421 301610 57487 301613
rect 60002 301610 60062 302190
rect 219390 302160 220064 302220
rect 379838 302160 380052 302220
rect 217133 302154 217199 302157
rect 219390 302154 219450 302160
rect 217133 302152 219450 302154
rect 217133 302096 217138 302152
rect 217194 302096 219450 302152
rect 217133 302094 219450 302096
rect 377397 302154 377463 302157
rect 378041 302154 378107 302157
rect 379838 302154 379898 302160
rect 377397 302152 379898 302154
rect 377397 302096 377402 302152
rect 377458 302096 378046 302152
rect 378102 302096 379898 302152
rect 377397 302094 379898 302096
rect 217133 302091 217199 302094
rect 377397 302091 377463 302094
rect 378041 302091 378107 302094
rect 57421 301608 60062 301610
rect 57421 301552 57426 301608
rect 57482 301552 60062 301608
rect 57421 301550 60062 301552
rect 57421 301547 57487 301550
rect 583520 298604 584960 298844
rect 518985 293858 519051 293861
rect 519353 293858 519419 293861
rect 516558 293856 519419 293858
rect 516558 293800 518990 293856
rect 519046 293800 519358 293856
rect 519414 293800 519419 293856
rect 516558 293798 519419 293800
rect 516558 293350 516618 293798
rect 518985 293795 519051 293798
rect 519353 293795 519419 293798
rect -960 293028 480 293268
rect 196558 292770 196618 293350
rect 199193 292770 199259 292773
rect 199653 292770 199719 292773
rect 196558 292768 199719 292770
rect 196558 292712 199198 292768
rect 199254 292712 199658 292768
rect 199714 292712 199719 292768
rect 196558 292710 199719 292712
rect 356562 292770 356622 293350
rect 359089 292770 359155 292773
rect 359273 292770 359339 292773
rect 356562 292768 359339 292770
rect 356562 292712 359094 292768
rect 359150 292712 359278 292768
rect 359334 292712 359339 292768
rect 356562 292710 359339 292712
rect 199193 292707 199259 292710
rect 199653 292707 199719 292710
rect 359089 292707 359155 292710
rect 359273 292707 359339 292710
rect 518893 292498 518959 292501
rect 519537 292498 519603 292501
rect 516558 292496 519603 292498
rect 516558 292440 518898 292496
rect 518954 292440 519542 292496
rect 519598 292440 519603 292496
rect 516558 292438 519603 292440
rect 359089 291818 359155 291821
rect 359549 291818 359615 291821
rect 356562 291816 359615 291818
rect 356562 291760 359094 291816
rect 359150 291760 359554 291816
rect 359610 291760 359615 291816
rect 356562 291758 359615 291760
rect 356562 291718 356622 291758
rect 359089 291755 359155 291758
rect 359549 291755 359615 291758
rect 516558 291718 516618 292438
rect 518893 292435 518959 292438
rect 519537 292435 519603 292438
rect 196558 291682 196618 291718
rect 198733 291682 198799 291685
rect 199469 291682 199535 291685
rect 196558 291680 199535 291682
rect 196558 291624 198738 291680
rect 198794 291624 199474 291680
rect 199530 291624 199535 291680
rect 196558 291622 199535 291624
rect 198733 291619 198799 291622
rect 199469 291619 199535 291622
rect 199101 291002 199167 291005
rect 199561 291002 199627 291005
rect 358997 291002 359063 291005
rect 359549 291002 359615 291005
rect 196558 291000 199627 291002
rect 196558 290944 199106 291000
rect 199162 290944 199566 291000
rect 199622 290944 199627 291000
rect 196558 290942 199627 290944
rect 196558 290358 196618 290942
rect 199101 290939 199167 290942
rect 199561 290939 199627 290942
rect 356562 291000 359615 291002
rect 356562 290944 359002 291000
rect 359058 290944 359554 291000
rect 359610 290944 359615 291000
rect 356562 290942 359615 290944
rect 356562 290358 356622 290942
rect 358997 290939 359063 290942
rect 359549 290939 359615 290942
rect 516558 290322 516618 290358
rect 519077 290322 519143 290325
rect 519629 290322 519695 290325
rect 516558 290320 519695 290322
rect 516558 290264 519082 290320
rect 519138 290264 519634 290320
rect 519690 290264 519695 290320
rect 516558 290262 519695 290264
rect 519077 290259 519143 290262
rect 519629 290259 519695 290262
rect 358813 289778 358879 289781
rect 359457 289778 359523 289781
rect 358813 289776 359523 289778
rect 358813 289720 358818 289776
rect 358874 289720 359462 289776
rect 359518 289720 359523 289776
rect 358813 289718 359523 289720
rect 358813 289715 358879 289718
rect 359457 289715 359523 289718
rect 196558 288826 196618 288862
rect 198917 288826 198983 288829
rect 196558 288824 198983 288826
rect 196558 288768 198922 288824
rect 198978 288768 198983 288824
rect 196558 288766 198983 288768
rect 356562 288826 356622 288862
rect 358813 288826 358879 288829
rect 356562 288824 358879 288826
rect 356562 288768 358818 288824
rect 358874 288768 358879 288824
rect 356562 288766 358879 288768
rect 516558 288826 516618 288862
rect 519169 288826 519235 288829
rect 520181 288826 520247 288829
rect 516558 288824 520247 288826
rect 516558 288768 519174 288824
rect 519230 288768 520186 288824
rect 520242 288768 520247 288824
rect 516558 288766 520247 288768
rect 198917 288763 198983 288766
rect 358813 288763 358879 288766
rect 519169 288763 519235 288766
rect 520181 288763 520247 288766
rect 199009 288418 199075 288421
rect 199745 288418 199811 288421
rect 199009 288416 199811 288418
rect 199009 288360 199014 288416
rect 199070 288360 199750 288416
rect 199806 288360 199811 288416
rect 199009 288358 199811 288360
rect 199009 288355 199075 288358
rect 199745 288355 199811 288358
rect 358997 288418 359063 288421
rect 359181 288418 359247 288421
rect 358997 288416 359247 288418
rect 358997 288360 359002 288416
rect 359058 288360 359186 288416
rect 359242 288360 359247 288416
rect 358997 288358 359247 288360
rect 358997 288355 359063 288358
rect 359181 288355 359247 288358
rect 196558 287602 196618 287638
rect 199009 287602 199075 287605
rect 196558 287600 199075 287602
rect 196558 287544 199014 287600
rect 199070 287544 199075 287600
rect 196558 287542 199075 287544
rect 356562 287602 356622 287638
rect 358997 287602 359063 287605
rect 356562 287600 359063 287602
rect 356562 287544 359002 287600
rect 359058 287544 359063 287600
rect 356562 287542 359063 287544
rect 516558 287602 516618 287638
rect 518985 287602 519051 287605
rect 516558 287600 519051 287602
rect 516558 287544 518990 287600
rect 519046 287544 519051 287600
rect 516558 287542 519051 287544
rect 199009 287539 199075 287542
rect 358997 287539 359063 287542
rect 518985 287539 519051 287542
rect 583520 285276 584960 285516
rect 58709 284202 58775 284205
rect 58709 284200 60062 284202
rect 58709 284144 58714 284200
rect 58770 284144 60062 284200
rect 58709 284142 60062 284144
rect 58709 284139 58775 284142
rect 60002 283966 60062 284142
rect 216673 284066 216739 284069
rect 376937 284066 377003 284069
rect 216673 284064 219450 284066
rect 216673 284008 216678 284064
rect 216734 284008 219450 284064
rect 216673 284006 219450 284008
rect 216673 284003 216739 284006
rect 219390 283996 219450 284006
rect 376937 284064 379530 284066
rect 376937 284008 376942 284064
rect 376998 284008 379530 284064
rect 376937 284006 379530 284008
rect 376937 284003 377003 284006
rect 379470 283996 379530 284006
rect 219390 283936 220064 283996
rect 379470 283936 380052 283996
rect 216673 282434 216739 282437
rect 216673 282432 219450 282434
rect 216673 282376 216678 282432
rect 216734 282376 219450 282432
rect 216673 282374 219450 282376
rect 216673 282371 216739 282374
rect 219390 282364 219450 282374
rect 59494 282304 60032 282364
rect 219390 282304 220064 282364
rect 379470 282304 380052 282364
rect 57513 282298 57579 282301
rect 59494 282298 59554 282304
rect 57513 282296 59554 282298
rect 57513 282240 57518 282296
rect 57574 282240 59554 282296
rect 57513 282238 59554 282240
rect 376937 282298 377003 282301
rect 379470 282298 379530 282304
rect 376937 282296 379530 282298
rect 376937 282240 376942 282296
rect 376998 282240 379530 282296
rect 376937 282238 379530 282240
rect 57513 282235 57579 282238
rect 376937 282235 377003 282238
rect 216765 282162 216831 282165
rect 376753 282162 376819 282165
rect 216765 282160 219450 282162
rect 216765 282104 216770 282160
rect 216826 282104 219450 282160
rect 216765 282102 219450 282104
rect 216765 282099 216831 282102
rect 219390 282092 219450 282102
rect 376753 282160 379530 282162
rect 376753 282104 376758 282160
rect 376814 282104 379530 282160
rect 376753 282102 379530 282104
rect 376753 282099 376819 282102
rect 379470 282092 379530 282102
rect 58801 282026 58867 282029
rect 60002 282026 60062 282062
rect 219390 282032 220064 282092
rect 379470 282032 380052 282092
rect 58801 282024 60062 282026
rect 58801 281968 58806 282024
rect 58862 281968 60062 282024
rect 58801 281966 60062 281968
rect 58801 281963 58867 281966
rect -960 279972 480 280212
rect 375005 274682 375071 274685
rect 376886 274682 376892 274684
rect 375005 274680 376892 274682
rect 375005 274624 375010 274680
rect 375066 274624 376892 274680
rect 375005 274622 376892 274624
rect 375005 274619 375071 274622
rect 376886 274620 376892 274622
rect 376956 274620 376962 274684
rect 95969 273868 96035 273869
rect 95904 273804 95910 273868
rect 95974 273866 96035 273868
rect 95974 273864 96066 273866
rect 96030 273808 96066 273864
rect 95974 273806 96066 273808
rect 95974 273804 96035 273806
rect 95969 273803 96035 273804
rect 266353 273732 266419 273733
rect 278037 273732 278103 273733
rect 266353 273730 266382 273732
rect 266290 273728 266382 273730
rect 266290 273672 266358 273728
rect 266290 273670 266382 273672
rect 266353 273668 266382 273670
rect 266446 273668 266452 273732
rect 278037 273730 278078 273732
rect 277986 273728 278078 273730
rect 277986 273672 278042 273728
rect 277986 273670 278078 273672
rect 278037 273668 278078 273670
rect 278142 273668 278148 273732
rect 266353 273667 266419 273668
rect 278037 273667 278103 273668
rect 110965 273596 111031 273597
rect 133413 273596 133479 273597
rect 135897 273596 135963 273597
rect 138473 273596 138539 273597
rect 140865 273596 140931 273597
rect 250713 273596 250779 273597
rect 273345 273596 273411 273597
rect 110965 273594 111006 273596
rect 110914 273592 111006 273594
rect 110914 273536 110970 273592
rect 110914 273534 111006 273536
rect 110965 273532 111006 273534
rect 111070 273532 111076 273596
rect 133413 273594 133446 273596
rect 133354 273592 133446 273594
rect 133354 273536 133418 273592
rect 133354 273534 133446 273536
rect 133413 273532 133446 273534
rect 133510 273532 133516 273596
rect 135888 273532 135894 273596
rect 135958 273594 135964 273596
rect 138472 273594 138478 273596
rect 135958 273534 136050 273594
rect 138386 273534 138478 273594
rect 135958 273532 135964 273534
rect 138472 273532 138478 273534
rect 138542 273532 138548 273596
rect 140865 273594 140926 273596
rect 140834 273592 140926 273594
rect 140834 273536 140870 273592
rect 140834 273534 140926 273536
rect 140865 273532 140926 273534
rect 140990 273532 140996 273596
rect 250713 273594 250742 273596
rect 250650 273592 250742 273594
rect 250650 273536 250718 273592
rect 250650 273534 250742 273536
rect 250713 273532 250742 273534
rect 250806 273532 250812 273596
rect 273312 273532 273318 273596
rect 273382 273594 273411 273596
rect 275737 273596 275803 273597
rect 283465 273596 283531 273597
rect 421097 273596 421163 273597
rect 450997 273596 451063 273597
rect 275737 273594 275766 273596
rect 273382 273592 273474 273594
rect 273406 273536 273474 273592
rect 273382 273534 273474 273536
rect 275674 273592 275766 273594
rect 275674 273536 275742 273592
rect 275674 273534 275766 273536
rect 273382 273532 273411 273534
rect 110965 273531 111031 273532
rect 133413 273531 133479 273532
rect 135897 273531 135963 273532
rect 138473 273531 138539 273532
rect 140865 273531 140931 273532
rect 250713 273531 250779 273532
rect 273345 273531 273411 273532
rect 275737 273532 275766 273534
rect 275830 273532 275836 273596
rect 283465 273594 283518 273596
rect 283426 273592 283518 273594
rect 283426 273536 283470 273592
rect 283426 273534 283518 273536
rect 283465 273532 283518 273534
rect 283582 273532 283588 273596
rect 421072 273532 421078 273596
rect 421142 273594 421163 273596
rect 450992 273594 450998 273596
rect 421142 273592 421234 273594
rect 421158 273536 421234 273592
rect 421142 273534 421234 273536
rect 450906 273534 450998 273594
rect 421142 273532 421163 273534
rect 450992 273532 450998 273534
rect 451062 273532 451068 273596
rect 275737 273531 275803 273532
rect 283465 273531 283531 273532
rect 421097 273531 421163 273532
rect 450997 273531 451063 273532
rect 376886 273396 376892 273460
rect 376956 273458 376962 273460
rect 422886 273458 422892 273460
rect 376956 273398 422892 273458
rect 376956 273396 376962 273398
rect 422886 273396 422892 273398
rect 422956 273396 422962 273460
rect 430982 273458 430988 273460
rect 423078 273398 430988 273458
rect 218421 273322 218487 273325
rect 285949 273324 286015 273325
rect 218830 273322 218836 273324
rect 218421 273320 218836 273322
rect 218421 273264 218426 273320
rect 218482 273264 218836 273320
rect 218421 273262 218836 273264
rect 218421 273259 218487 273262
rect 218830 273260 218836 273262
rect 218900 273260 218906 273324
rect 285949 273322 285996 273324
rect 285904 273320 285996 273322
rect 285904 273264 285954 273320
rect 285904 273262 285996 273264
rect 285949 273260 285996 273262
rect 286060 273260 286066 273324
rect 359406 273260 359412 273324
rect 359476 273322 359482 273324
rect 423078 273322 423138 273398
rect 430982 273396 430988 273398
rect 431052 273396 431058 273460
rect 423397 273324 423463 273325
rect 423765 273324 423831 273325
rect 426433 273324 426499 273325
rect 423397 273322 423444 273324
rect 359476 273262 423138 273322
rect 423352 273320 423444 273322
rect 423352 273264 423402 273320
rect 423352 273262 423444 273264
rect 359476 273260 359482 273262
rect 423397 273260 423444 273262
rect 423508 273260 423514 273324
rect 423765 273322 423812 273324
rect 423720 273320 423812 273322
rect 423720 273264 423770 273320
rect 423720 273262 423812 273264
rect 423765 273260 423812 273262
rect 423876 273260 423882 273324
rect 426382 273260 426388 273324
rect 426452 273322 426499 273324
rect 426452 273320 426544 273322
rect 426494 273264 426544 273320
rect 426452 273262 426544 273264
rect 426452 273260 426499 273262
rect 285949 273259 286015 273260
rect 423397 273259 423463 273260
rect 423765 273259 423831 273260
rect 426433 273259 426499 273260
rect 58801 273186 58867 273189
rect 100753 273188 100819 273189
rect 58801 273184 84210 273186
rect 58801 273128 58806 273184
rect 58862 273128 84210 273184
rect 58801 273126 84210 273128
rect 58801 273123 58867 273126
rect 84150 273050 84210 273126
rect 100702 273124 100708 273188
rect 100772 273186 100819 273188
rect 100772 273184 100864 273186
rect 100814 273128 100864 273184
rect 100772 273126 100864 273128
rect 100772 273124 100819 273126
rect 199326 273124 199332 273188
rect 199396 273186 199402 273188
rect 318374 273186 318380 273188
rect 199396 273126 318380 273186
rect 199396 273124 199402 273126
rect 318374 273124 318380 273126
rect 318444 273124 318450 273188
rect 359590 273124 359596 273188
rect 359660 273186 359666 273188
rect 485998 273186 486004 273188
rect 359660 273126 486004 273186
rect 359660 273124 359666 273126
rect 485998 273124 486004 273126
rect 486068 273124 486074 273188
rect 100753 273123 100819 273124
rect 102726 273050 102732 273052
rect 84150 272990 102732 273050
rect 102726 272988 102732 272990
rect 102796 272988 102802 273052
rect 196566 272988 196572 273052
rect 196636 273050 196642 273052
rect 311014 273050 311020 273052
rect 196636 272990 311020 273050
rect 196636 272988 196642 272990
rect 311014 272988 311020 272990
rect 311084 272988 311090 273052
rect 361113 273050 361179 273053
rect 483238 273050 483244 273052
rect 361113 273048 483244 273050
rect 361113 272992 361118 273048
rect 361174 272992 483244 273048
rect 361113 272990 483244 272992
rect 361113 272987 361179 272990
rect 483238 272988 483244 272990
rect 483308 272988 483314 273052
rect 76005 272916 76071 272917
rect 90725 272916 90791 272917
rect 93669 272916 93735 272917
rect 95877 272916 95943 272917
rect 98453 272916 98519 272917
rect 99373 272916 99439 272917
rect 76005 272914 76052 272916
rect 75960 272912 76052 272914
rect 75960 272856 76010 272912
rect 75960 272854 76052 272856
rect 76005 272852 76052 272854
rect 76116 272852 76122 272916
rect 90725 272914 90772 272916
rect 90680 272912 90772 272914
rect 90680 272856 90730 272912
rect 90680 272854 90772 272856
rect 90725 272852 90772 272854
rect 90836 272852 90842 272916
rect 93669 272914 93716 272916
rect 93624 272912 93716 272914
rect 93624 272856 93674 272912
rect 93624 272854 93716 272856
rect 93669 272852 93716 272854
rect 93780 272852 93786 272916
rect 95877 272914 95924 272916
rect 95832 272912 95924 272914
rect 95832 272856 95882 272912
rect 95832 272854 95924 272856
rect 95877 272852 95924 272854
rect 95988 272852 95994 272916
rect 98453 272914 98500 272916
rect 98408 272912 98500 272914
rect 98408 272856 98458 272912
rect 98408 272854 98500 272856
rect 98453 272852 98500 272854
rect 98564 272852 98570 272916
rect 99373 272914 99420 272916
rect 99328 272912 99420 272914
rect 99328 272856 99378 272912
rect 99328 272854 99420 272856
rect 99373 272852 99420 272854
rect 99484 272852 99490 272916
rect 199510 272852 199516 272916
rect 199580 272914 199586 272916
rect 287973 272914 288039 272917
rect 288157 272916 288223 272917
rect 290917 272916 290983 272917
rect 293309 272916 293375 272917
rect 300853 272916 300919 272917
rect 288157 272914 288204 272916
rect 199580 272912 288039 272914
rect 199580 272856 287978 272912
rect 288034 272856 288039 272912
rect 199580 272854 288039 272856
rect 288112 272912 288204 272914
rect 288112 272856 288162 272912
rect 288112 272854 288204 272856
rect 199580 272852 199586 272854
rect 76005 272851 76071 272852
rect 90725 272851 90791 272852
rect 93669 272851 93735 272852
rect 95877 272851 95943 272852
rect 98453 272851 98519 272852
rect 99373 272851 99439 272852
rect 287973 272851 288039 272854
rect 288157 272852 288204 272854
rect 288268 272852 288274 272916
rect 290917 272914 290964 272916
rect 290872 272912 290964 272914
rect 290872 272856 290922 272912
rect 290872 272854 290964 272856
rect 290917 272852 290964 272854
rect 291028 272852 291034 272916
rect 293309 272914 293356 272916
rect 293264 272912 293356 272914
rect 293264 272856 293314 272912
rect 293264 272854 293356 272856
rect 293309 272852 293356 272854
rect 293420 272852 293426 272916
rect 300853 272914 300900 272916
rect 300808 272912 300900 272914
rect 300808 272856 300858 272912
rect 300808 272854 300900 272856
rect 300853 272852 300900 272854
rect 300964 272852 300970 272916
rect 371601 272914 371667 272917
rect 480846 272914 480852 272916
rect 371601 272912 480852 272914
rect 371601 272856 371606 272912
rect 371662 272856 480852 272912
rect 371601 272854 480852 272856
rect 288157 272851 288223 272852
rect 290917 272851 290983 272852
rect 293309 272851 293375 272852
rect 300853 272851 300919 272852
rect 371601 272851 371667 272854
rect 480846 272852 480852 272854
rect 480916 272852 480922 272916
rect 60825 272778 60891 272781
rect 61009 272778 61075 272781
rect 298461 272780 298527 272781
rect 425973 272780 426039 272781
rect 428181 272780 428247 272781
rect 431125 272780 431191 272781
rect 468477 272780 468543 272781
rect 470869 272780 470935 272781
rect 473445 272780 473511 272781
rect 103830 272778 103836 272780
rect 60825 272776 103836 272778
rect 60825 272720 60830 272776
rect 60886 272720 61014 272776
rect 61070 272720 103836 272776
rect 60825 272718 103836 272720
rect 60825 272715 60891 272718
rect 61009 272715 61075 272718
rect 103830 272716 103836 272718
rect 103900 272716 103906 272780
rect 217358 272716 217364 272780
rect 217428 272778 217434 272780
rect 298461 272778 298508 272780
rect 217428 272718 296730 272778
rect 298416 272776 298508 272778
rect 298416 272720 298466 272776
rect 298416 272718 298508 272720
rect 217428 272716 217434 272718
rect 61745 272642 61811 272645
rect 143533 272644 143599 272645
rect 117998 272642 118004 272644
rect 61745 272640 118004 272642
rect 61745 272584 61750 272640
rect 61806 272584 118004 272640
rect 61745 272582 118004 272584
rect 61745 272579 61811 272582
rect 117998 272580 118004 272582
rect 118068 272580 118074 272644
rect 143533 272642 143580 272644
rect 143488 272640 143580 272642
rect 143488 272584 143538 272640
rect 143488 272582 143580 272584
rect 143533 272580 143580 272582
rect 143644 272580 143650 272644
rect 287973 272642 288039 272645
rect 295926 272642 295932 272644
rect 287973 272640 295932 272642
rect 287973 272584 287978 272640
rect 288034 272584 295932 272640
rect 287973 272582 295932 272584
rect 143533 272579 143599 272580
rect 287973 272579 288039 272582
rect 295926 272580 295932 272582
rect 295996 272580 296002 272644
rect 296670 272642 296730 272718
rect 298461 272716 298508 272718
rect 298572 272716 298578 272780
rect 425973 272778 426020 272780
rect 425928 272776 426020 272778
rect 425928 272720 425978 272776
rect 425928 272718 426020 272720
rect 425973 272716 426020 272718
rect 426084 272716 426090 272780
rect 428181 272778 428228 272780
rect 428136 272776 428228 272778
rect 428136 272720 428186 272776
rect 428136 272718 428228 272720
rect 428181 272716 428228 272718
rect 428292 272716 428298 272780
rect 431125 272778 431172 272780
rect 431080 272776 431172 272778
rect 431080 272720 431130 272776
rect 431080 272718 431172 272720
rect 431125 272716 431172 272718
rect 431236 272716 431242 272780
rect 468477 272778 468524 272780
rect 468432 272776 468524 272778
rect 468432 272720 468482 272776
rect 468432 272718 468524 272720
rect 468477 272716 468524 272718
rect 468588 272716 468594 272780
rect 470869 272778 470916 272780
rect 470824 272776 470916 272778
rect 470824 272720 470874 272776
rect 470824 272718 470916 272720
rect 470869 272716 470916 272718
rect 470980 272716 470986 272780
rect 473445 272778 473492 272780
rect 473400 272776 473492 272778
rect 473400 272720 473450 272776
rect 473400 272718 473492 272720
rect 473445 272716 473492 272718
rect 473556 272716 473562 272780
rect 298461 272715 298527 272716
rect 425973 272715 426039 272716
rect 428181 272715 428247 272716
rect 431125 272715 431191 272716
rect 468477 272715 468543 272716
rect 470869 272715 470935 272716
rect 473445 272715 473511 272716
rect 305821 272644 305887 272645
rect 320909 272644 320975 272645
rect 475837 272644 475903 272645
rect 478413 272644 478479 272645
rect 303470 272642 303476 272644
rect 296670 272582 303476 272642
rect 303470 272580 303476 272582
rect 303540 272580 303546 272644
rect 305821 272642 305868 272644
rect 305776 272640 305868 272642
rect 305776 272584 305826 272640
rect 305776 272582 305868 272584
rect 305821 272580 305868 272582
rect 305932 272580 305938 272644
rect 320909 272642 320956 272644
rect 320864 272640 320956 272642
rect 320864 272584 320914 272640
rect 320864 272582 320956 272584
rect 320909 272580 320956 272582
rect 321020 272580 321026 272644
rect 475837 272642 475884 272644
rect 475792 272640 475884 272642
rect 475792 272584 475842 272640
rect 475792 272582 475884 272584
rect 475837 272580 475884 272582
rect 475948 272580 475954 272644
rect 478413 272642 478460 272644
rect 478368 272640 478460 272642
rect 478368 272584 478418 272640
rect 478368 272582 478460 272584
rect 478413 272580 478460 272582
rect 478524 272580 478530 272644
rect 305821 272579 305887 272580
rect 320909 272579 320975 272580
rect 475837 272579 475903 272580
rect 478413 272579 478479 272580
rect 61469 272506 61535 272509
rect 119102 272506 119108 272508
rect 61469 272504 119108 272506
rect 61469 272448 61474 272504
rect 61530 272448 119108 272504
rect 61469 272446 119108 272448
rect 61469 272443 61535 272446
rect 119102 272444 119108 272446
rect 119172 272444 119178 272508
rect 96981 272372 97047 272373
rect 96981 272370 97028 272372
rect 96936 272368 97028 272370
rect 96936 272312 96986 272368
rect 96936 272310 97028 272312
rect 96981 272308 97028 272310
rect 97092 272308 97098 272372
rect 96981 272307 97047 272308
rect 113541 272236 113607 272237
rect 235993 272236 236059 272237
rect 113541 272234 113588 272236
rect 113496 272232 113588 272234
rect 113496 272176 113546 272232
rect 113496 272174 113588 272176
rect 113541 272172 113588 272174
rect 113652 272172 113658 272236
rect 235942 272172 235948 272236
rect 236012 272234 236059 272236
rect 265157 272236 265223 272237
rect 401685 272236 401751 272237
rect 416037 272236 416103 272237
rect 437933 272236 437999 272237
rect 455781 272236 455847 272237
rect 265157 272234 265204 272236
rect 236012 272232 236104 272234
rect 236054 272176 236104 272232
rect 236012 272174 236104 272176
rect 265112 272232 265204 272234
rect 265112 272176 265162 272232
rect 265112 272174 265204 272176
rect 236012 272172 236059 272174
rect 113541 272171 113607 272172
rect 235993 272171 236059 272172
rect 265157 272172 265204 272174
rect 265268 272172 265274 272236
rect 401685 272234 401732 272236
rect 401640 272232 401732 272234
rect 401640 272176 401690 272232
rect 401640 272174 401732 272176
rect 401685 272172 401732 272174
rect 401796 272172 401802 272236
rect 416037 272234 416084 272236
rect 415992 272232 416084 272234
rect 415992 272176 416042 272232
rect 415992 272174 416084 272176
rect 416037 272172 416084 272174
rect 416148 272172 416154 272236
rect 437933 272234 437980 272236
rect 437888 272232 437980 272234
rect 437888 272176 437938 272232
rect 437888 272174 437980 272176
rect 437933 272172 437980 272174
rect 438044 272172 438050 272236
rect 455781 272234 455828 272236
rect 455736 272232 455828 272234
rect 455736 272176 455786 272232
rect 455736 272174 455828 272176
rect 455781 272172 455828 272174
rect 455892 272172 455898 272236
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 265157 272171 265223 272172
rect 401685 272171 401751 272172
rect 416037 272171 416103 272172
rect 437933 272171 437999 272172
rect 455781 272171 455847 272172
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 49049 271826 49115 271829
rect 49233 271826 49299 271829
rect 75913 271826 75979 271829
rect 77150 271826 77156 271828
rect 49049 271824 55230 271826
rect 49049 271768 49054 271824
rect 49110 271768 49238 271824
rect 49294 271768 55230 271824
rect 49049 271766 55230 271768
rect 49049 271763 49115 271766
rect 49233 271763 49299 271766
rect 55170 271690 55230 271766
rect 75913 271824 77156 271826
rect 75913 271768 75918 271824
rect 75974 271768 77156 271824
rect 75913 271766 77156 271768
rect 75913 271763 75979 271766
rect 77150 271764 77156 271766
rect 77220 271764 77226 271828
rect 82813 271826 82879 271829
rect 83038 271826 83044 271828
rect 82813 271824 83044 271826
rect 82813 271768 82818 271824
rect 82874 271768 83044 271824
rect 82813 271766 83044 271768
rect 82813 271763 82879 271766
rect 83038 271764 83044 271766
rect 83108 271764 83114 271828
rect 83958 271764 83964 271828
rect 84028 271826 84034 271828
rect 84193 271826 84259 271829
rect 84028 271824 84259 271826
rect 84028 271768 84198 271824
rect 84254 271768 84259 271824
rect 84028 271766 84259 271768
rect 84028 271764 84034 271766
rect 84193 271763 84259 271766
rect 86953 271826 87019 271829
rect 87638 271826 87644 271828
rect 86953 271824 87644 271826
rect 86953 271768 86958 271824
rect 87014 271768 87644 271824
rect 86953 271766 87644 271768
rect 86953 271763 87019 271766
rect 87638 271764 87644 271766
rect 87708 271764 87714 271828
rect 94221 271826 94287 271829
rect 94446 271826 94452 271828
rect 94221 271824 94452 271826
rect 94221 271768 94226 271824
rect 94282 271768 94452 271824
rect 94221 271766 94452 271768
rect 94221 271763 94287 271766
rect 94446 271764 94452 271766
rect 94516 271764 94522 271828
rect 97993 271826 98059 271829
rect 98126 271826 98132 271828
rect 97993 271824 98132 271826
rect 97993 271768 97998 271824
rect 98054 271768 98132 271824
rect 97993 271766 98132 271768
rect 97993 271763 98059 271766
rect 98126 271764 98132 271766
rect 98196 271764 98202 271828
rect 100753 271826 100819 271829
rect 114461 271828 114527 271829
rect 101806 271826 101812 271828
rect 100753 271824 101812 271826
rect 100753 271768 100758 271824
rect 100814 271768 101812 271824
rect 100753 271766 101812 271768
rect 100753 271763 100819 271766
rect 101806 271764 101812 271766
rect 101876 271764 101882 271828
rect 114461 271826 114508 271828
rect 114416 271824 114508 271826
rect 114416 271768 114466 271824
rect 114416 271766 114508 271768
rect 114461 271764 114508 271766
rect 114572 271764 114578 271828
rect 123201 271826 123267 271829
rect 123518 271826 123524 271828
rect 123201 271824 123524 271826
rect 123201 271768 123206 271824
rect 123262 271768 123524 271824
rect 123201 271766 123524 271768
rect 114461 271763 114527 271764
rect 123201 271763 123267 271766
rect 123518 271764 123524 271766
rect 123588 271764 123594 271828
rect 128353 271826 128419 271829
rect 128670 271826 128676 271828
rect 128353 271824 128676 271826
rect 128353 271768 128358 271824
rect 128414 271768 128676 271824
rect 128353 271766 128676 271768
rect 128353 271763 128419 271766
rect 128670 271764 128676 271766
rect 128740 271764 128746 271828
rect 129733 271826 129799 271829
rect 130878 271826 130884 271828
rect 129733 271824 130884 271826
rect 129733 271768 129738 271824
rect 129794 271768 130884 271824
rect 129733 271766 130884 271768
rect 129733 271763 129799 271766
rect 130878 271764 130884 271766
rect 130948 271764 130954 271828
rect 150934 271764 150940 271828
rect 151004 271826 151010 271828
rect 151353 271826 151419 271829
rect 151004 271824 151419 271826
rect 151004 271768 151358 271824
rect 151414 271768 151419 271824
rect 151004 271766 151419 271768
rect 151004 271764 151010 271766
rect 151353 271763 151419 271766
rect 154062 271764 154068 271828
rect 154132 271826 154138 271828
rect 154481 271826 154547 271829
rect 154132 271824 154547 271826
rect 154132 271768 154486 271824
rect 154542 271768 154547 271824
rect 154132 271766 154547 271768
rect 154132 271764 154138 271766
rect 154481 271763 154547 271766
rect 155902 271764 155908 271828
rect 155972 271826 155978 271828
rect 157241 271826 157307 271829
rect 155972 271824 157307 271826
rect 155972 271768 157246 271824
rect 157302 271768 157307 271824
rect 155972 271766 157307 271768
rect 155972 271764 155978 271766
rect 157241 271763 157307 271766
rect 196617 271826 196683 271829
rect 196750 271826 196756 271828
rect 196617 271824 196756 271826
rect 196617 271768 196622 271824
rect 196678 271768 196756 271824
rect 196617 271766 196756 271768
rect 196617 271763 196683 271766
rect 196750 271764 196756 271766
rect 196820 271764 196826 271828
rect 268193 271826 268259 271829
rect 268694 271826 268700 271828
rect 268193 271824 268700 271826
rect 268193 271768 268198 271824
rect 268254 271768 268700 271824
rect 268193 271766 268700 271768
rect 268193 271763 268259 271766
rect 268694 271764 268700 271766
rect 268764 271764 268770 271828
rect 270493 271826 270559 271829
rect 270902 271826 270908 271828
rect 270493 271824 270908 271826
rect 270493 271768 270498 271824
rect 270554 271768 270908 271824
rect 270493 271766 270908 271768
rect 270493 271763 270559 271766
rect 270902 271764 270908 271766
rect 270972 271764 270978 271828
rect 276013 271826 276079 271829
rect 276238 271826 276244 271828
rect 276013 271824 276244 271826
rect 276013 271768 276018 271824
rect 276074 271768 276244 271824
rect 276013 271766 276244 271768
rect 276013 271763 276079 271766
rect 276238 271764 276244 271766
rect 276308 271764 276314 271828
rect 280153 271826 280219 271829
rect 280838 271826 280844 271828
rect 280153 271824 280844 271826
rect 280153 271768 280158 271824
rect 280214 271768 280844 271824
rect 280153 271766 280844 271768
rect 280153 271763 280219 271766
rect 280838 271764 280844 271766
rect 280908 271764 280914 271828
rect 307753 271826 307819 271829
rect 308622 271826 308628 271828
rect 307753 271824 308628 271826
rect 307753 271768 307758 271824
rect 307814 271768 308628 271824
rect 307753 271766 308628 271768
rect 307753 271763 307819 271766
rect 308622 271764 308628 271766
rect 308692 271764 308698 271828
rect 313273 271826 313339 271829
rect 313406 271826 313412 271828
rect 313273 271824 313412 271826
rect 313273 271768 313278 271824
rect 313334 271768 313412 271824
rect 313273 271766 313412 271768
rect 313273 271763 313339 271766
rect 313406 271764 313412 271766
rect 313476 271764 313482 271828
rect 343398 271764 343404 271828
rect 343468 271826 343474 271828
rect 343541 271826 343607 271829
rect 343468 271824 343607 271826
rect 343468 271768 343546 271824
rect 343602 271768 343607 271824
rect 343468 271766 343607 271768
rect 343468 271764 343474 271766
rect 343541 271763 343607 271766
rect 402973 271828 403039 271829
rect 402973 271824 403020 271828
rect 403084 271826 403090 271828
rect 412817 271826 412883 271829
rect 418470 271826 418476 271828
rect 402973 271768 402978 271824
rect 402973 271764 403020 271768
rect 403084 271766 403130 271826
rect 412817 271824 418476 271826
rect 412817 271768 412822 271824
rect 412878 271768 418476 271824
rect 412817 271766 418476 271768
rect 403084 271764 403090 271766
rect 402973 271763 403039 271764
rect 412817 271763 412883 271766
rect 418470 271764 418476 271766
rect 418540 271764 418546 271828
rect 433333 271826 433399 271829
rect 433558 271826 433564 271828
rect 433333 271824 433564 271826
rect 433333 271768 433338 271824
rect 433394 271768 433564 271824
rect 433333 271766 433564 271768
rect 433333 271763 433399 271766
rect 433558 271764 433564 271766
rect 433628 271764 433634 271828
rect 434713 271826 434779 271829
rect 435950 271826 435956 271828
rect 434713 271824 435956 271826
rect 434713 271768 434718 271824
rect 434774 271768 435956 271824
rect 434713 271766 435956 271768
rect 434713 271763 434779 271766
rect 435950 271764 435956 271766
rect 436020 271764 436026 271828
rect 437473 271826 437539 271829
rect 438526 271826 438532 271828
rect 437473 271824 438532 271826
rect 437473 271768 437478 271824
rect 437534 271768 438532 271824
rect 437473 271766 438532 271768
rect 437473 271763 437539 271766
rect 438526 271764 438532 271766
rect 438596 271764 438602 271828
rect 445753 271826 445819 271829
rect 445886 271826 445892 271828
rect 445753 271824 445892 271826
rect 445753 271768 445758 271824
rect 445814 271768 445892 271824
rect 445753 271766 445892 271768
rect 445753 271763 445819 271766
rect 445886 271764 445892 271766
rect 445956 271764 445962 271828
rect 447133 271826 447199 271829
rect 448278 271826 448284 271828
rect 447133 271824 448284 271826
rect 447133 271768 447138 271824
rect 447194 271768 448284 271824
rect 447133 271766 448284 271768
rect 447133 271763 447199 271766
rect 448278 271764 448284 271766
rect 448348 271764 448354 271828
rect 452653 271826 452719 271829
rect 453430 271826 453436 271828
rect 452653 271824 453436 271826
rect 452653 271768 452658 271824
rect 452714 271768 453436 271824
rect 452653 271766 453436 271768
rect 452653 271763 452719 271766
rect 453430 271764 453436 271766
rect 453500 271764 453506 271828
rect 458173 271826 458239 271829
rect 458398 271826 458404 271828
rect 458173 271824 458404 271826
rect 458173 271768 458178 271824
rect 458234 271768 458404 271824
rect 458173 271766 458404 271768
rect 458173 271763 458239 271766
rect 458398 271764 458404 271766
rect 458468 271764 458474 271828
rect 84653 271692 84719 271693
rect 81934 271690 81940 271692
rect 55170 271630 81940 271690
rect 81934 271628 81940 271630
rect 82004 271628 82010 271692
rect 84653 271690 84700 271692
rect 84608 271688 84700 271690
rect 84608 271632 84658 271688
rect 84608 271630 84700 271632
rect 84653 271628 84700 271630
rect 84764 271628 84770 271692
rect 103513 271690 103579 271693
rect 103830 271690 103836 271692
rect 103513 271688 103836 271690
rect 103513 271632 103518 271688
rect 103574 271632 103836 271688
rect 103513 271630 103836 271632
rect 84653 271627 84719 271628
rect 103513 271627 103579 271630
rect 103830 271628 103836 271630
rect 103900 271628 103906 271692
rect 120073 271690 120139 271693
rect 120758 271690 120764 271692
rect 120073 271688 120764 271690
rect 120073 271632 120078 271688
rect 120134 271632 120764 271688
rect 120073 271630 120764 271632
rect 120073 271627 120139 271630
rect 120758 271628 120764 271630
rect 120828 271628 120834 271692
rect 125593 271690 125659 271693
rect 125910 271690 125916 271692
rect 125593 271688 125916 271690
rect 125593 271632 125598 271688
rect 125654 271632 125916 271688
rect 125593 271630 125916 271632
rect 125593 271627 125659 271630
rect 125910 271628 125916 271630
rect 125980 271628 125986 271692
rect 158478 271628 158484 271692
rect 158548 271690 158554 271692
rect 158621 271690 158687 271693
rect 158548 271688 158687 271690
rect 158548 271632 158626 271688
rect 158682 271632 158687 271688
rect 158548 271630 158687 271632
rect 158548 271628 158554 271630
rect 158621 271627 158687 271630
rect 160870 271628 160876 271692
rect 160940 271690 160946 271692
rect 161289 271690 161355 271693
rect 160940 271688 161355 271690
rect 160940 271632 161294 271688
rect 161350 271632 161355 271688
rect 160940 271630 161355 271632
rect 160940 271628 160946 271630
rect 161289 271627 161355 271630
rect 163446 271628 163452 271692
rect 163516 271690 163522 271692
rect 164141 271690 164207 271693
rect 163516 271688 164207 271690
rect 163516 271632 164146 271688
rect 164202 271632 164207 271688
rect 163516 271630 164207 271632
rect 163516 271628 163522 271630
rect 164141 271627 164207 271630
rect 166022 271628 166028 271692
rect 166092 271690 166098 271692
rect 198774 271690 198780 271692
rect 166092 271630 198780 271690
rect 166092 271628 166098 271630
rect 198774 271628 198780 271630
rect 198844 271628 198850 271692
rect 216029 271690 216095 271693
rect 315062 271690 315068 271692
rect 216029 271688 315068 271690
rect 216029 271632 216034 271688
rect 216090 271632 315068 271688
rect 216029 271630 315068 271632
rect 216029 271627 216095 271630
rect 315062 271628 315068 271630
rect 315132 271628 315138 271692
rect 376385 271690 376451 271693
rect 465942 271690 465948 271692
rect 376385 271688 465948 271690
rect 376385 271632 376390 271688
rect 376446 271632 465948 271688
rect 376385 271630 465948 271632
rect 376385 271627 376451 271630
rect 465942 271628 465948 271630
rect 466012 271628 466018 271692
rect 503110 271628 503116 271692
rect 503180 271690 503186 271692
rect 503621 271690 503687 271693
rect 503180 271688 503687 271690
rect 503180 271632 503626 271688
rect 503682 271632 503687 271688
rect 503180 271630 503687 271632
rect 503180 271628 503186 271630
rect 503621 271627 503687 271630
rect 46933 271554 46999 271557
rect 115933 271556 115999 271557
rect 80462 271554 80468 271556
rect 46933 271552 80468 271554
rect 46933 271496 46938 271552
rect 46994 271496 80468 271552
rect 46933 271494 80468 271496
rect 46933 271491 46999 271494
rect 80462 271492 80468 271494
rect 80532 271492 80538 271556
rect 115933 271554 115980 271556
rect 115888 271552 115980 271554
rect 115888 271496 115938 271552
rect 115888 271494 115980 271496
rect 115933 271492 115980 271494
rect 116044 271492 116050 271556
rect 117313 271554 117379 271557
rect 118366 271554 118372 271556
rect 117313 271552 118372 271554
rect 117313 271496 117318 271552
rect 117374 271496 118372 271552
rect 117313 271494 118372 271496
rect 115933 271491 115999 271492
rect 117313 271491 117379 271494
rect 118366 271492 118372 271494
rect 118436 271492 118442 271556
rect 127617 271554 127683 271557
rect 196617 271554 196683 271557
rect 127617 271552 196683 271554
rect 127617 271496 127622 271552
rect 127678 271496 196622 271552
rect 196678 271496 196683 271552
rect 127617 271494 196683 271496
rect 127617 271491 127683 271494
rect 196617 271491 196683 271494
rect 217174 271492 217180 271556
rect 217244 271554 217250 271556
rect 258257 271554 258323 271557
rect 263593 271556 263659 271557
rect 258390 271554 258396 271556
rect 217244 271494 258090 271554
rect 217244 271492 217250 271494
rect 51901 271418 51967 271421
rect 52361 271418 52427 271421
rect 65333 271418 65399 271421
rect 51901 271416 65399 271418
rect 51901 271360 51906 271416
rect 51962 271360 52366 271416
rect 52422 271360 65338 271416
rect 65394 271360 65399 271416
rect 51901 271358 65399 271360
rect 51901 271355 51967 271358
rect 52361 271355 52427 271358
rect 65333 271355 65399 271358
rect 100753 271418 100819 271421
rect 101070 271418 101076 271420
rect 100753 271416 101076 271418
rect 100753 271360 100758 271416
rect 100814 271360 101076 271416
rect 100753 271358 101076 271360
rect 100753 271355 100819 271358
rect 101070 271356 101076 271358
rect 101140 271356 101146 271420
rect 104893 271418 104959 271421
rect 105854 271418 105860 271420
rect 104893 271416 105860 271418
rect 104893 271360 104898 271416
rect 104954 271360 105860 271416
rect 104893 271358 105860 271360
rect 104893 271355 104959 271358
rect 105854 271356 105860 271358
rect 105924 271356 105930 271420
rect 183134 271356 183140 271420
rect 183204 271418 183210 271420
rect 183461 271418 183527 271421
rect 183204 271416 183527 271418
rect 183204 271360 183466 271416
rect 183522 271360 183527 271416
rect 183204 271358 183527 271360
rect 183204 271356 183210 271358
rect 183461 271355 183527 271358
rect 216397 271418 216463 271421
rect 216581 271418 216647 271421
rect 237046 271418 237052 271420
rect 216397 271416 237052 271418
rect 216397 271360 216402 271416
rect 216458 271360 216586 271416
rect 216642 271360 237052 271416
rect 216397 271358 237052 271360
rect 216397 271355 216463 271358
rect 216581 271355 216647 271358
rect 237046 271356 237052 271358
rect 237116 271356 237122 271420
rect 258030 271418 258090 271494
rect 258257 271552 258396 271554
rect 258257 271496 258262 271552
rect 258318 271496 258396 271552
rect 258257 271494 258396 271496
rect 258257 271491 258323 271494
rect 258390 271492 258396 271494
rect 258460 271492 258466 271556
rect 263542 271492 263548 271556
rect 263612 271554 263659 271556
rect 264973 271554 265039 271557
rect 265934 271554 265940 271556
rect 263612 271552 263704 271554
rect 263654 271496 263704 271552
rect 263612 271494 263704 271496
rect 264973 271552 265940 271554
rect 264973 271496 264978 271552
rect 265034 271496 265940 271552
rect 264973 271494 265940 271496
rect 263612 271492 263659 271494
rect 263593 271491 263659 271492
rect 264973 271491 265039 271494
rect 265934 271492 265940 271494
rect 266004 271492 266010 271556
rect 268009 271554 268075 271557
rect 268326 271554 268332 271556
rect 268009 271552 268332 271554
rect 268009 271496 268014 271552
rect 268070 271496 268332 271552
rect 268009 271494 268332 271496
rect 268009 271491 268075 271494
rect 268326 271492 268332 271494
rect 268396 271492 268402 271556
rect 271873 271554 271939 271557
rect 272558 271554 272564 271556
rect 271873 271552 272564 271554
rect 271873 271496 271878 271552
rect 271934 271496 272564 271552
rect 271873 271494 272564 271496
rect 271873 271491 271939 271494
rect 272558 271492 272564 271494
rect 272628 271492 272634 271556
rect 276974 271492 276980 271556
rect 277044 271554 277050 271556
rect 277117 271554 277183 271557
rect 277044 271552 277183 271554
rect 277044 271496 277122 271552
rect 277178 271496 277183 271552
rect 277044 271494 277183 271496
rect 277044 271492 277050 271494
rect 277117 271491 277183 271494
rect 343214 271492 343220 271556
rect 343284 271554 343290 271556
rect 343541 271554 343607 271557
rect 343284 271552 343607 271554
rect 343284 271496 343546 271552
rect 343602 271496 343607 271552
rect 343284 271494 343607 271496
rect 343284 271492 343290 271494
rect 343541 271491 343607 271494
rect 376201 271554 376267 271557
rect 460974 271554 460980 271556
rect 376201 271552 460980 271554
rect 376201 271496 376206 271552
rect 376262 271496 460980 271552
rect 376201 271494 460980 271496
rect 376201 271491 376267 271494
rect 460974 271492 460980 271494
rect 461044 271492 461050 271556
rect 273478 271418 273484 271420
rect 258030 271358 273484 271418
rect 273478 271356 273484 271358
rect 273548 271356 273554 271420
rect 277669 271418 277735 271421
rect 278446 271418 278452 271420
rect 277669 271416 278452 271418
rect 277669 271360 277674 271416
rect 277730 271360 278452 271416
rect 277669 271358 278452 271360
rect 277669 271355 277735 271358
rect 278446 271356 278452 271358
rect 278516 271356 278522 271420
rect 377806 271356 377812 271420
rect 377876 271418 377882 271420
rect 412817 271418 412883 271421
rect 415526 271418 415532 271420
rect 377876 271416 412883 271418
rect 377876 271360 412822 271416
rect 412878 271360 412883 271416
rect 377876 271358 412883 271360
rect 377876 271356 377882 271358
rect 412817 271355 412883 271358
rect 412958 271358 415532 271418
rect 45921 271282 45987 271285
rect 59629 271282 59695 271285
rect 45921 271280 59695 271282
rect 45921 271224 45926 271280
rect 45982 271224 59634 271280
rect 59690 271224 59695 271280
rect 45921 271222 59695 271224
rect 45921 271219 45987 271222
rect 59629 271219 59695 271222
rect 252553 271282 252619 271285
rect 253606 271282 253612 271284
rect 252553 271280 253612 271282
rect 252553 271224 252558 271280
rect 252614 271224 253612 271280
rect 252553 271222 253612 271224
rect 252553 271219 252619 271222
rect 253606 271220 253612 271222
rect 253676 271220 253682 271284
rect 260833 271282 260899 271285
rect 260966 271282 260972 271284
rect 260833 271280 260972 271282
rect 260833 271224 260838 271280
rect 260894 271224 260972 271280
rect 260833 271222 260972 271224
rect 260833 271219 260899 271222
rect 260966 271220 260972 271222
rect 261036 271220 261042 271284
rect 396022 271282 396028 271284
rect 383610 271222 396028 271282
rect 52453 271146 52519 271149
rect 52821 271146 52887 271149
rect 67357 271146 67423 271149
rect 52453 271144 67423 271146
rect 52453 271088 52458 271144
rect 52514 271088 52826 271144
rect 52882 271088 67362 271144
rect 67418 271088 67423 271144
rect 52453 271086 67423 271088
rect 52453 271083 52519 271086
rect 52821 271083 52887 271086
rect 67357 271083 67423 271086
rect 77293 271146 77359 271149
rect 88333 271148 88399 271149
rect 183461 271148 183527 271149
rect 78254 271146 78260 271148
rect 77293 271144 78260 271146
rect 77293 271088 77298 271144
rect 77354 271088 78260 271144
rect 77293 271086 78260 271088
rect 77293 271083 77359 271086
rect 78254 271084 78260 271086
rect 78324 271084 78330 271148
rect 88333 271146 88380 271148
rect 88288 271144 88380 271146
rect 88288 271088 88338 271144
rect 88288 271086 88380 271088
rect 88333 271084 88380 271086
rect 88444 271084 88450 271148
rect 183461 271146 183508 271148
rect 183416 271144 183508 271146
rect 183416 271088 183466 271144
rect 183416 271086 183508 271088
rect 183461 271084 183508 271086
rect 183572 271084 183578 271148
rect 247033 271146 247099 271149
rect 248270 271146 248276 271148
rect 247033 271144 248276 271146
rect 247033 271088 247038 271144
rect 247094 271088 248276 271144
rect 247033 271086 248276 271088
rect 88333 271083 88399 271084
rect 183461 271083 183527 271084
rect 247033 271083 247099 271086
rect 248270 271084 248276 271086
rect 248340 271084 248346 271148
rect 255313 271146 255379 271149
rect 256182 271146 256188 271148
rect 255313 271144 256188 271146
rect 255313 271088 255318 271144
rect 255374 271088 256188 271144
rect 255313 271086 256188 271088
rect 255313 271083 255379 271086
rect 256182 271084 256188 271086
rect 256252 271084 256258 271148
rect 78673 271010 78739 271013
rect 79542 271010 79548 271012
rect 78673 271008 79548 271010
rect 78673 270952 78678 271008
rect 78734 270952 79548 271008
rect 78673 270950 79548 270952
rect 78673 270947 78739 270950
rect 79542 270948 79548 270950
rect 79612 270948 79618 271012
rect 88333 271010 88399 271013
rect 88742 271010 88748 271012
rect 88333 271008 88748 271010
rect 88333 270952 88338 271008
rect 88394 270952 88748 271008
rect 88333 270950 88748 270952
rect 88333 270947 88399 270950
rect 88742 270948 88748 270950
rect 88812 270948 88818 271012
rect 89713 271010 89779 271013
rect 90030 271010 90036 271012
rect 89713 271008 90036 271010
rect 89713 270952 89718 271008
rect 89774 270952 90036 271008
rect 89713 270950 90036 270952
rect 89713 270947 89779 270950
rect 90030 270948 90036 270950
rect 90100 270948 90106 271012
rect 106365 271010 106431 271013
rect 107510 271010 107516 271012
rect 106365 271008 107516 271010
rect 106365 270952 106370 271008
rect 106426 270952 107516 271008
rect 106365 270950 107516 270952
rect 106365 270947 106431 270950
rect 107510 270948 107516 270950
rect 107580 270948 107586 271012
rect 107653 271010 107719 271013
rect 108614 271010 108620 271012
rect 107653 271008 108620 271010
rect 107653 270952 107658 271008
rect 107714 270952 108620 271008
rect 107653 270950 108620 270952
rect 107653 270947 107719 270950
rect 108614 270948 108620 270950
rect 108684 270948 108690 271012
rect 111793 271010 111859 271013
rect 112110 271010 112116 271012
rect 111793 271008 112116 271010
rect 111793 270952 111798 271008
rect 111854 270952 112116 271008
rect 111793 270950 112116 270952
rect 111793 270947 111859 270950
rect 112110 270948 112116 270950
rect 112180 270948 112186 271012
rect 207749 271010 207815 271013
rect 325550 271010 325556 271012
rect 207749 271008 325556 271010
rect 207749 270952 207754 271008
rect 207810 270952 325556 271008
rect 207749 270950 325556 270952
rect 207749 270947 207815 270950
rect 325550 270948 325556 270950
rect 325620 270948 325626 271012
rect 374545 271010 374611 271013
rect 374913 271010 374979 271013
rect 383610 271010 383670 271222
rect 396022 271220 396028 271222
rect 396092 271220 396098 271284
rect 396717 271282 396783 271285
rect 412958 271282 413018 271358
rect 415526 271356 415532 271358
rect 415596 271356 415602 271420
rect 440233 271418 440299 271421
rect 440918 271418 440924 271420
rect 440233 271416 440924 271418
rect 440233 271360 440238 271416
rect 440294 271360 440924 271416
rect 440233 271358 440924 271360
rect 440233 271355 440299 271358
rect 440918 271356 440924 271358
rect 440988 271356 440994 271420
rect 396717 271280 413018 271282
rect 396717 271224 396722 271280
rect 396778 271224 413018 271280
rect 396717 271222 413018 271224
rect 413093 271282 413159 271285
rect 413686 271282 413692 271284
rect 413093 271280 413692 271282
rect 413093 271224 413098 271280
rect 413154 271224 413692 271280
rect 413093 271222 413692 271224
rect 396717 271219 396783 271222
rect 413093 271219 413159 271222
rect 413686 271220 413692 271222
rect 413756 271220 413762 271284
rect 439262 271220 439268 271284
rect 439332 271282 439338 271284
rect 440141 271282 440207 271285
rect 439332 271280 440207 271282
rect 439332 271224 440146 271280
rect 440202 271224 440207 271280
rect 439332 271222 440207 271224
rect 439332 271220 439338 271222
rect 440141 271219 440207 271222
rect 442993 271282 443059 271285
rect 443494 271282 443500 271284
rect 442993 271280 443500 271282
rect 442993 271224 442998 271280
rect 443054 271224 443500 271280
rect 442993 271222 443500 271224
rect 442993 271219 443059 271222
rect 443494 271220 443500 271222
rect 443564 271220 443570 271284
rect 503478 271220 503484 271284
rect 503548 271282 503554 271284
rect 503621 271282 503687 271285
rect 503548 271280 503687 271282
rect 503548 271224 503626 271280
rect 503682 271224 503687 271280
rect 503548 271222 503687 271224
rect 503548 271220 503554 271222
rect 503621 271219 503687 271222
rect 409873 271146 409939 271149
rect 410742 271146 410748 271148
rect 409873 271144 410748 271146
rect 409873 271088 409878 271144
rect 409934 271088 410748 271144
rect 409873 271086 410748 271088
rect 409873 271083 409939 271086
rect 410742 271084 410748 271086
rect 410812 271084 410818 271148
rect 414013 271146 414079 271149
rect 414422 271146 414428 271148
rect 414013 271144 414428 271146
rect 414013 271088 414018 271144
rect 414074 271088 414428 271144
rect 414013 271086 414428 271088
rect 414013 271083 414079 271086
rect 414422 271084 414428 271086
rect 414492 271084 414498 271148
rect 416773 271146 416839 271149
rect 416998 271146 417004 271148
rect 416773 271144 417004 271146
rect 416773 271088 416778 271144
rect 416834 271088 417004 271144
rect 416773 271086 417004 271088
rect 416773 271083 416839 271086
rect 416998 271084 417004 271086
rect 417068 271084 417074 271148
rect 433333 271146 433399 271149
rect 434662 271146 434668 271148
rect 433333 271144 434668 271146
rect 433333 271088 433338 271144
rect 433394 271088 434668 271144
rect 433333 271086 434668 271088
rect 433333 271083 433399 271086
rect 434662 271084 434668 271086
rect 434732 271084 434738 271148
rect 374545 271008 383670 271010
rect 374545 270952 374550 271008
rect 374606 270952 374918 271008
rect 374974 270952 383670 271008
rect 374545 270950 383670 270952
rect 404353 271010 404419 271013
rect 405038 271010 405044 271012
rect 404353 271008 405044 271010
rect 404353 270952 404358 271008
rect 404414 270952 405044 271008
rect 404353 270950 405044 270952
rect 374545 270947 374611 270950
rect 374913 270947 374979 270950
rect 404353 270947 404419 270950
rect 405038 270948 405044 270950
rect 405108 270948 405114 271012
rect 407113 271010 407179 271013
rect 408166 271010 408172 271012
rect 407113 271008 408172 271010
rect 407113 270952 407118 271008
rect 407174 270952 408172 271008
rect 407113 270950 408172 270952
rect 407113 270947 407179 270950
rect 408166 270948 408172 270950
rect 408236 270948 408242 271012
rect 411253 271010 411319 271013
rect 412398 271010 412404 271012
rect 411253 271008 412404 271010
rect 411253 270952 411258 271008
rect 411314 270952 412404 271008
rect 411253 270950 412404 270952
rect 411253 270947 411319 270950
rect 412398 270948 412404 270950
rect 412468 270948 412474 271012
rect 427077 271010 427143 271013
rect 428590 271010 428596 271012
rect 427077 271008 428596 271010
rect 427077 270952 427082 271008
rect 427138 270952 428596 271008
rect 427077 270950 428596 270952
rect 427077 270947 427143 270950
rect 428590 270948 428596 270950
rect 428660 270948 428666 271012
rect 429193 271010 429259 271013
rect 429694 271010 429700 271012
rect 429193 271008 429700 271010
rect 429193 270952 429198 271008
rect 429254 270952 429700 271008
rect 429193 270950 429700 270952
rect 429193 270947 429259 270950
rect 429694 270948 429700 270950
rect 429764 270948 429770 271012
rect 433374 270948 433380 271012
rect 433444 271010 433450 271012
rect 434713 271010 434779 271013
rect 433444 271008 434779 271010
rect 433444 270952 434718 271008
rect 434774 270952 434779 271008
rect 433444 270950 434779 270952
rect 433444 270948 433450 270950
rect 434713 270947 434779 270950
rect 435766 270948 435772 271012
rect 435836 271010 435842 271012
rect 436093 271010 436159 271013
rect 435836 271008 436159 271010
rect 435836 270952 436098 271008
rect 436154 270952 436159 271008
rect 435836 270950 436159 270952
rect 435836 270948 435842 270950
rect 436093 270947 436159 270950
rect 85573 270874 85639 270877
rect 86534 270874 86540 270876
rect 85573 270872 86540 270874
rect 85573 270816 85578 270872
rect 85634 270816 86540 270872
rect 85573 270814 86540 270816
rect 85573 270811 85639 270814
rect 86534 270812 86540 270814
rect 86604 270812 86610 270876
rect 92473 270874 92539 270877
rect 93342 270874 93348 270876
rect 92473 270872 93348 270874
rect 92473 270816 92478 270872
rect 92534 270816 93348 270872
rect 92473 270814 93348 270816
rect 92473 270811 92539 270814
rect 93342 270812 93348 270814
rect 93412 270812 93418 270876
rect 104893 270874 104959 270877
rect 105302 270874 105308 270876
rect 104893 270872 105308 270874
rect 104893 270816 104898 270872
rect 104954 270816 105308 270872
rect 104893 270814 105308 270816
rect 104893 270811 104959 270814
rect 105302 270812 105308 270814
rect 105372 270812 105378 270876
rect 106273 270874 106339 270877
rect 106406 270874 106412 270876
rect 106273 270872 106412 270874
rect 106273 270816 106278 270872
rect 106334 270816 106412 270872
rect 106273 270814 106412 270816
rect 106273 270811 106339 270814
rect 106406 270812 106412 270814
rect 106476 270812 106482 270876
rect 253933 270874 253999 270877
rect 254526 270874 254532 270876
rect 253933 270872 254532 270874
rect 253933 270816 253938 270872
rect 253994 270816 254532 270872
rect 253933 270814 254532 270816
rect 253933 270811 253999 270814
rect 254526 270812 254532 270814
rect 254596 270812 254602 270876
rect 278998 270812 279004 270876
rect 279068 270874 279074 270876
rect 280061 270874 280127 270877
rect 279068 270872 280127 270874
rect 279068 270816 280066 270872
rect 280122 270816 280127 270872
rect 279068 270814 280127 270816
rect 279068 270812 279074 270814
rect 280061 270811 280127 270814
rect 372245 270874 372311 270877
rect 462630 270874 462636 270876
rect 372245 270872 462636 270874
rect 372245 270816 372250 270872
rect 372306 270816 462636 270872
rect 372245 270814 462636 270816
rect 372245 270811 372311 270814
rect 462630 270812 462636 270814
rect 462700 270812 462706 270876
rect 110413 270738 110479 270741
rect 111190 270738 111196 270740
rect 110413 270736 111196 270738
rect 110413 270680 110418 270736
rect 110474 270680 111196 270736
rect 110413 270678 111196 270680
rect 110413 270675 110479 270678
rect 111190 270676 111196 270678
rect 111260 270676 111266 270740
rect 244222 270676 244228 270740
rect 244292 270738 244298 270740
rect 244365 270738 244431 270741
rect 244292 270736 244431 270738
rect 244292 270680 244370 270736
rect 244426 270680 244431 270736
rect 244292 270678 244431 270680
rect 244292 270676 244298 270678
rect 244365 270675 244431 270678
rect 251265 270738 251331 270741
rect 252318 270738 252324 270740
rect 251265 270736 252324 270738
rect 251265 270680 251270 270736
rect 251326 270680 252324 270736
rect 251265 270678 252324 270680
rect 251265 270675 251331 270678
rect 252318 270676 252324 270678
rect 252388 270676 252394 270740
rect 255313 270738 255379 270741
rect 255814 270738 255820 270740
rect 255313 270736 255820 270738
rect 255313 270680 255318 270736
rect 255374 270680 255820 270736
rect 255313 270678 255820 270680
rect 255313 270675 255379 270678
rect 255814 270676 255820 270678
rect 255884 270676 255890 270740
rect 259545 270738 259611 270741
rect 260598 270738 260604 270740
rect 259545 270736 260604 270738
rect 259545 270680 259550 270736
rect 259606 270680 260604 270736
rect 259545 270678 260604 270680
rect 259545 270675 259611 270678
rect 260598 270676 260604 270678
rect 260668 270676 260674 270740
rect 412909 270738 412975 270741
rect 413318 270738 413324 270740
rect 412909 270736 413324 270738
rect 412909 270680 412914 270736
rect 412970 270680 413324 270736
rect 412909 270678 413324 270680
rect 412909 270675 412975 270678
rect 413318 270676 413324 270678
rect 413388 270676 413394 270740
rect 418245 270738 418311 270741
rect 419206 270738 419212 270740
rect 418245 270736 419212 270738
rect 418245 270680 418250 270736
rect 418306 270680 419212 270736
rect 418245 270678 419212 270680
rect 418245 270675 418311 270678
rect 419206 270676 419212 270678
rect 419276 270676 419282 270740
rect 425697 270738 425763 270741
rect 427670 270738 427676 270740
rect 425697 270736 427676 270738
rect 425697 270680 425702 270736
rect 425758 270680 427676 270736
rect 425697 270678 427676 270680
rect 425697 270675 425763 270678
rect 427670 270676 427676 270678
rect 427740 270676 427746 270740
rect 59629 270602 59695 270605
rect 60825 270602 60891 270605
rect 59629 270600 60891 270602
rect 59629 270544 59634 270600
rect 59690 270544 60830 270600
rect 60886 270544 60891 270600
rect 59629 270542 60891 270544
rect 59629 270539 59695 270542
rect 60825 270539 60891 270542
rect 91093 270602 91159 270605
rect 91318 270602 91324 270604
rect 91093 270600 91324 270602
rect 91093 270544 91098 270600
rect 91154 270544 91324 270600
rect 91093 270542 91324 270544
rect 91093 270539 91159 270542
rect 91318 270540 91324 270542
rect 91388 270540 91394 270604
rect 107745 270602 107811 270605
rect 108246 270602 108252 270604
rect 107745 270600 108252 270602
rect 107745 270544 107750 270600
rect 107806 270544 108252 270600
rect 107745 270542 108252 270544
rect 107745 270539 107811 270542
rect 108246 270540 108252 270542
rect 108316 270540 108322 270604
rect 109033 270602 109099 270605
rect 113173 270604 113239 270605
rect 115841 270604 115907 270605
rect 109534 270602 109540 270604
rect 109033 270600 109540 270602
rect 109033 270544 109038 270600
rect 109094 270544 109540 270600
rect 109033 270542 109540 270544
rect 109033 270539 109099 270542
rect 109534 270540 109540 270542
rect 109604 270540 109610 270604
rect 113173 270600 113220 270604
rect 113284 270602 113290 270604
rect 113173 270544 113178 270600
rect 113173 270540 113220 270544
rect 113284 270542 113330 270602
rect 113284 270540 113290 270542
rect 115790 270540 115796 270604
rect 115860 270602 115907 270604
rect 115860 270600 115952 270602
rect 115902 270544 115952 270600
rect 115860 270542 115952 270544
rect 115860 270540 115907 270542
rect 117078 270540 117084 270604
rect 117148 270602 117154 270604
rect 117221 270602 117287 270605
rect 117148 270600 117287 270602
rect 117148 270544 117226 270600
rect 117282 270544 117287 270600
rect 117148 270542 117287 270544
rect 117148 270540 117154 270542
rect 113173 270539 113239 270540
rect 115841 270539 115907 270540
rect 117221 270539 117287 270542
rect 144913 270602 144979 270605
rect 145598 270602 145604 270604
rect 144913 270600 145604 270602
rect 144913 270544 144918 270600
rect 144974 270544 145604 270600
rect 144913 270542 145604 270544
rect 144913 270539 144979 270542
rect 145598 270540 145604 270542
rect 145668 270540 145674 270604
rect 147673 270602 147739 270605
rect 148542 270602 148548 270604
rect 147673 270600 148548 270602
rect 147673 270544 147678 270600
rect 147734 270544 148548 270600
rect 147673 270542 148548 270544
rect 147673 270539 147739 270542
rect 148542 270540 148548 270542
rect 148612 270540 148618 270604
rect 239121 270602 239187 270605
rect 242893 270604 242959 270605
rect 239254 270602 239260 270604
rect 239121 270600 239260 270602
rect 239121 270544 239126 270600
rect 239182 270544 239260 270600
rect 239121 270542 239260 270544
rect 239121 270539 239187 270542
rect 239254 270540 239260 270542
rect 239324 270540 239330 270604
rect 242893 270602 242940 270604
rect 242848 270600 242940 270602
rect 242848 270544 242898 270600
rect 242848 270542 242940 270544
rect 242893 270540 242940 270542
rect 243004 270540 243010 270604
rect 244273 270602 244339 270605
rect 245326 270602 245332 270604
rect 244273 270600 245332 270602
rect 244273 270544 244278 270600
rect 244334 270544 245332 270600
rect 244273 270542 245332 270544
rect 242893 270539 242959 270540
rect 244273 270539 244339 270542
rect 245326 270540 245332 270542
rect 245396 270540 245402 270604
rect 245653 270602 245719 270605
rect 246430 270602 246436 270604
rect 245653 270600 246436 270602
rect 245653 270544 245658 270600
rect 245714 270544 246436 270600
rect 245653 270542 246436 270544
rect 245653 270539 245719 270542
rect 246430 270540 246436 270542
rect 246500 270540 246506 270604
rect 247033 270602 247099 270605
rect 247718 270602 247724 270604
rect 247033 270600 247724 270602
rect 247033 270544 247038 270600
rect 247094 270544 247724 270600
rect 247033 270542 247724 270544
rect 247033 270539 247099 270542
rect 247718 270540 247724 270542
rect 247788 270540 247794 270604
rect 248505 270602 248571 270605
rect 248638 270602 248644 270604
rect 248505 270600 248644 270602
rect 248505 270544 248510 270600
rect 248566 270544 248644 270600
rect 248505 270542 248644 270544
rect 248505 270539 248571 270542
rect 248638 270540 248644 270542
rect 248708 270540 248714 270604
rect 249793 270602 249859 270605
rect 251173 270604 251239 270605
rect 250110 270602 250116 270604
rect 249793 270600 250116 270602
rect 249793 270544 249798 270600
rect 249854 270544 250116 270600
rect 249793 270542 250116 270544
rect 249793 270539 249859 270542
rect 250110 270540 250116 270542
rect 250180 270540 250186 270604
rect 251173 270602 251220 270604
rect 251128 270600 251220 270602
rect 251128 270544 251178 270600
rect 251128 270542 251220 270544
rect 251173 270540 251220 270542
rect 251284 270540 251290 270604
rect 252553 270602 252619 270605
rect 253422 270602 253428 270604
rect 252553 270600 253428 270602
rect 252553 270544 252558 270600
rect 252614 270544 253428 270600
rect 252553 270542 253428 270544
rect 251173 270539 251239 270540
rect 252553 270539 252619 270542
rect 253422 270540 253428 270542
rect 253492 270540 253498 270604
rect 256693 270602 256759 270605
rect 256918 270602 256924 270604
rect 256693 270600 256924 270602
rect 256693 270544 256698 270600
rect 256754 270544 256924 270600
rect 256693 270542 256924 270544
rect 256693 270539 256759 270542
rect 256918 270540 256924 270542
rect 256988 270540 256994 270604
rect 258073 270602 258139 270605
rect 259453 270604 259519 270605
rect 258390 270602 258396 270604
rect 258073 270600 258396 270602
rect 258073 270544 258078 270600
rect 258134 270544 258396 270600
rect 258073 270542 258396 270544
rect 258073 270539 258139 270542
rect 258390 270540 258396 270542
rect 258460 270540 258466 270604
rect 259453 270602 259500 270604
rect 259408 270600 259500 270602
rect 259408 270544 259458 270600
rect 259408 270542 259500 270544
rect 259453 270540 259500 270542
rect 259564 270540 259570 270604
rect 260833 270602 260899 270605
rect 262070 270602 262076 270604
rect 260833 270600 262076 270602
rect 260833 270544 260838 270600
rect 260894 270544 262076 270600
rect 260833 270542 262076 270544
rect 259453 270539 259519 270540
rect 260833 270539 260899 270542
rect 262070 270540 262076 270542
rect 262140 270540 262146 270604
rect 262213 270602 262279 270605
rect 262806 270602 262812 270604
rect 262213 270600 262812 270602
rect 262213 270544 262218 270600
rect 262274 270544 262812 270600
rect 262213 270542 262812 270544
rect 262213 270539 262279 270542
rect 262806 270540 262812 270542
rect 262876 270540 262882 270604
rect 263593 270602 263659 270605
rect 263910 270602 263916 270604
rect 263593 270600 263916 270602
rect 263593 270544 263598 270600
rect 263654 270544 263916 270600
rect 263593 270542 263916 270544
rect 263593 270539 263659 270542
rect 263910 270540 263916 270542
rect 263980 270540 263986 270604
rect 266353 270602 266419 270605
rect 267590 270602 267596 270604
rect 266353 270600 267596 270602
rect 266353 270544 266358 270600
rect 266414 270544 267596 270600
rect 266353 270542 267596 270544
rect 266353 270539 266419 270542
rect 267590 270540 267596 270542
rect 267660 270540 267666 270604
rect 269113 270602 269179 270605
rect 269798 270602 269804 270604
rect 269113 270600 269804 270602
rect 269113 270544 269118 270600
rect 269174 270544 269804 270600
rect 269113 270542 269804 270544
rect 269113 270539 269179 270542
rect 269798 270540 269804 270542
rect 269868 270540 269874 270604
rect 270493 270602 270559 270605
rect 271270 270602 271276 270604
rect 270493 270600 271276 270602
rect 270493 270544 270498 270600
rect 270554 270544 271276 270600
rect 270493 270542 271276 270544
rect 270493 270539 270559 270542
rect 271270 270540 271276 270542
rect 271340 270540 271346 270604
rect 273161 270602 273227 270605
rect 274398 270602 274404 270604
rect 273161 270600 274404 270602
rect 273161 270544 273166 270600
rect 273222 270544 274404 270600
rect 273161 270542 274404 270544
rect 273161 270539 273227 270542
rect 274398 270540 274404 270542
rect 274468 270540 274474 270604
rect 396073 270602 396139 270605
rect 397453 270604 397519 270605
rect 397126 270602 397132 270604
rect 396073 270600 397132 270602
rect 396073 270544 396078 270600
rect 396134 270544 397132 270600
rect 396073 270542 397132 270544
rect 396073 270539 396139 270542
rect 397126 270540 397132 270542
rect 397196 270540 397202 270604
rect 397453 270602 397500 270604
rect 397408 270600 397500 270602
rect 397408 270544 397458 270600
rect 397408 270542 397500 270544
rect 397453 270540 397500 270542
rect 397564 270540 397570 270604
rect 398833 270602 398899 270605
rect 399518 270602 399524 270604
rect 398833 270600 399524 270602
rect 398833 270544 398838 270600
rect 398894 270544 399524 270600
rect 398833 270542 399524 270544
rect 397453 270539 397519 270540
rect 398833 270539 398899 270542
rect 399518 270540 399524 270542
rect 399588 270540 399594 270604
rect 400213 270602 400279 270605
rect 400438 270602 400444 270604
rect 400213 270600 400444 270602
rect 400213 270544 400218 270600
rect 400274 270544 400444 270600
rect 400213 270542 400444 270544
rect 400213 270539 400279 270542
rect 400438 270540 400444 270542
rect 400508 270540 400514 270604
rect 403525 270602 403591 270605
rect 404118 270602 404124 270604
rect 403525 270600 404124 270602
rect 403525 270544 403530 270600
rect 403586 270544 404124 270600
rect 403525 270542 404124 270544
rect 403525 270539 403591 270542
rect 404118 270540 404124 270542
rect 404188 270540 404194 270604
rect 405733 270602 405799 270605
rect 406510 270602 406516 270604
rect 405733 270600 406516 270602
rect 405733 270544 405738 270600
rect 405794 270544 406516 270600
rect 405733 270542 406516 270544
rect 405733 270539 405799 270542
rect 406510 270540 406516 270542
rect 406580 270540 406586 270604
rect 407113 270602 407179 270605
rect 407614 270602 407620 270604
rect 407113 270600 407620 270602
rect 407113 270544 407118 270600
rect 407174 270544 407620 270600
rect 407113 270542 407620 270544
rect 407113 270539 407179 270542
rect 407614 270540 407620 270542
rect 407684 270540 407690 270604
rect 408493 270602 408559 270605
rect 408718 270602 408724 270604
rect 408493 270600 408724 270602
rect 408493 270544 408498 270600
rect 408554 270544 408724 270600
rect 408493 270542 408724 270544
rect 408493 270539 408559 270542
rect 408718 270540 408724 270542
rect 408788 270540 408794 270604
rect 409873 270602 409939 270605
rect 411345 270604 411411 270605
rect 418153 270604 418219 270605
rect 410006 270602 410012 270604
rect 409873 270600 410012 270602
rect 409873 270544 409878 270600
rect 409934 270544 410012 270600
rect 409873 270542 410012 270544
rect 409873 270539 409939 270542
rect 410006 270540 410012 270542
rect 410076 270540 410082 270604
rect 411294 270540 411300 270604
rect 411364 270602 411411 270604
rect 411364 270600 411456 270602
rect 411406 270544 411456 270600
rect 411364 270542 411456 270544
rect 411364 270540 411411 270542
rect 418102 270540 418108 270604
rect 418172 270602 418219 270604
rect 419533 270602 419599 270605
rect 420678 270602 420684 270604
rect 418172 270600 418264 270602
rect 418214 270544 418264 270600
rect 418172 270542 418264 270544
rect 419533 270600 420684 270602
rect 419533 270544 419538 270600
rect 419594 270544 420684 270600
rect 419533 270542 420684 270544
rect 418172 270540 418219 270542
rect 411345 270539 411411 270540
rect 418153 270539 418219 270540
rect 419533 270539 419599 270542
rect 420678 270540 420684 270542
rect 420748 270540 420754 270604
rect 420913 270602 420979 270605
rect 421782 270602 421788 270604
rect 420913 270600 421788 270602
rect 420913 270544 420918 270600
rect 420974 270544 421788 270600
rect 420913 270542 421788 270544
rect 420913 270539 420979 270542
rect 421782 270540 421788 270542
rect 421852 270540 421858 270604
rect 436185 270602 436251 270605
rect 436870 270602 436876 270604
rect 436185 270600 436876 270602
rect 436185 270544 436190 270600
rect 436246 270544 436876 270600
rect 436185 270542 436876 270544
rect 436185 270539 436251 270542
rect 436870 270540 436876 270542
rect 436940 270540 436946 270604
rect 91502 270466 91508 270468
rect 64830 270406 91508 270466
rect 51901 270330 51967 270333
rect 57462 270330 57468 270332
rect 51901 270328 57468 270330
rect 51901 270272 51906 270328
rect 51962 270272 57468 270328
rect 51901 270270 57468 270272
rect 51901 270267 51967 270270
rect 57462 270268 57468 270270
rect 57532 270330 57538 270332
rect 64830 270330 64890 270406
rect 91502 270404 91508 270406
rect 91572 270404 91578 270468
rect 206645 270466 206711 270469
rect 323342 270466 323348 270468
rect 206645 270464 323348 270466
rect 206645 270408 206650 270464
rect 206706 270408 323348 270464
rect 206645 270406 323348 270408
rect 206645 270403 206711 270406
rect 323342 270404 323348 270406
rect 323412 270404 323418 270468
rect 374361 270466 374427 270469
rect 432270 270466 432276 270468
rect 373950 270464 432276 270466
rect 373950 270408 374366 270464
rect 374422 270408 432276 270464
rect 373950 270406 432276 270408
rect 57532 270270 64890 270330
rect 214373 270330 214439 270333
rect 214925 270330 214991 270333
rect 216857 270330 216923 270333
rect 241646 270330 241652 270332
rect 214373 270328 216322 270330
rect 214373 270272 214378 270328
rect 214434 270272 214930 270328
rect 214986 270272 216322 270328
rect 214373 270270 216322 270272
rect 57532 270268 57538 270270
rect 214373 270267 214439 270270
rect 214925 270267 214991 270270
rect 216262 270194 216322 270270
rect 216857 270328 241652 270330
rect 216857 270272 216862 270328
rect 216918 270272 241652 270328
rect 216857 270270 241652 270272
rect 216857 270267 216923 270270
rect 241646 270268 241652 270270
rect 241716 270268 241722 270332
rect 240542 270194 240548 270196
rect 216262 270134 240548 270194
rect 240542 270132 240548 270134
rect 240612 270132 240618 270196
rect 212257 270058 212323 270061
rect 215569 270058 215635 270061
rect 216857 270058 216923 270061
rect 212257 270056 216923 270058
rect 212257 270000 212262 270056
rect 212318 270000 215574 270056
rect 215630 270000 216862 270056
rect 216918 270000 216923 270056
rect 212257 269998 216923 270000
rect 212257 269995 212323 269998
rect 215569 269995 215635 269998
rect 216857 269995 216923 269998
rect 373165 270058 373231 270061
rect 373950 270058 374010 270406
rect 374361 270403 374427 270406
rect 432270 270404 432276 270406
rect 432340 270404 432346 270468
rect 378685 270330 378751 270333
rect 425278 270330 425284 270332
rect 378685 270328 425284 270330
rect 378685 270272 378690 270328
rect 378746 270272 425284 270328
rect 378685 270270 425284 270272
rect 378685 270267 378751 270270
rect 425278 270268 425284 270270
rect 425348 270268 425354 270332
rect 373165 270056 374010 270058
rect 373165 270000 373170 270056
rect 373226 270000 374010 270056
rect 373165 269998 374010 270000
rect 373165 269995 373231 269998
rect 208025 269786 208091 269789
rect 209313 269786 209379 269789
rect 238150 269786 238156 269788
rect 208025 269784 238156 269786
rect 208025 269728 208030 269784
rect 208086 269728 209318 269784
rect 209374 269728 238156 269784
rect 208025 269726 238156 269728
rect 208025 269723 208091 269726
rect 209313 269723 209379 269726
rect 238150 269724 238156 269726
rect 238220 269724 238226 269788
rect 372981 269786 373047 269789
rect 389265 269786 389331 269789
rect 372981 269784 389331 269786
rect 372981 269728 372986 269784
rect 373042 269728 389270 269784
rect 389326 269728 389331 269784
rect 372981 269726 389331 269728
rect 372981 269723 373047 269726
rect 389265 269723 389331 269726
rect 375414 269044 375420 269108
rect 375484 269106 375490 269108
rect 376661 269106 376727 269109
rect 375484 269104 376727 269106
rect 375484 269048 376666 269104
rect 376722 269048 376727 269104
rect 375484 269046 376727 269048
rect 375484 269044 375490 269046
rect 376661 269043 376727 269046
rect 44766 268364 44772 268428
rect 44836 268426 44842 268428
rect 46565 268426 46631 268429
rect 77845 268426 77911 268429
rect 44836 268424 77911 268426
rect 44836 268368 46570 268424
rect 46626 268368 77850 268424
rect 77906 268368 77911 268424
rect 44836 268366 77911 268368
rect 44836 268364 44842 268366
rect 46565 268363 46631 268366
rect 77845 268363 77911 268366
rect 217542 268364 217548 268428
rect 217612 268426 217618 268428
rect 229185 268426 229251 268429
rect 217612 268424 229251 268426
rect 217612 268368 229190 268424
rect 229246 268368 229251 268424
rect 217612 268366 229251 268368
rect 217612 268364 217618 268366
rect 229185 268363 229251 268366
rect 46606 267684 46612 267748
rect 46676 267746 46682 267748
rect 53097 267746 53163 267749
rect 46676 267744 53163 267746
rect 46676 267688 53102 267744
rect 53158 267688 53163 267744
rect 46676 267686 53163 267688
rect 46676 267684 46682 267686
rect 53097 267683 53163 267686
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 53046 254010 53052 254012
rect 6870 253950 53052 254010
rect 53046 253948 53052 253950
rect 53116 253948 53122 254012
rect 190862 253676 190868 253740
rect 190932 253738 190938 253740
rect 191741 253738 191807 253741
rect 190932 253736 191807 253738
rect 190932 253680 191746 253736
rect 191802 253680 191807 253736
rect 190932 253678 191807 253680
rect 190932 253676 190938 253678
rect 191741 253675 191807 253678
rect 339718 253404 339724 253468
rect 339788 253466 339794 253468
rect 340781 253466 340847 253469
rect 339788 253464 340847 253466
rect 339788 253408 340786 253464
rect 340842 253408 340847 253464
rect 339788 253406 340847 253408
rect 339788 253404 339794 253406
rect 340781 253403 340847 253406
rect 499798 253268 499804 253332
rect 499868 253330 499874 253332
rect 500861 253330 500927 253333
rect 499868 253328 500927 253330
rect 499868 253272 500866 253328
rect 500922 253272 500927 253328
rect 499868 253270 500927 253272
rect 499868 253268 499874 253270
rect 500861 253267 500927 253270
rect 178534 253132 178540 253196
rect 178604 253194 178610 253196
rect 179321 253194 179387 253197
rect 178604 253192 179387 253194
rect 178604 253136 179326 253192
rect 179382 253136 179387 253192
rect 178604 253134 179387 253136
rect 178604 253132 178610 253134
rect 179321 253131 179387 253134
rect 179638 253132 179644 253196
rect 179708 253194 179714 253196
rect 180517 253194 180583 253197
rect 179708 253192 180583 253194
rect 179708 253136 180522 253192
rect 180578 253136 180583 253192
rect 179708 253134 180583 253136
rect 179708 253132 179714 253134
rect 180517 253131 180583 253134
rect 350942 253132 350948 253196
rect 351012 253194 351018 253196
rect 351821 253194 351887 253197
rect 351012 253192 351887 253194
rect 351012 253136 351826 253192
rect 351882 253136 351887 253192
rect 351012 253134 351887 253136
rect 351012 253132 351018 253134
rect 351821 253131 351887 253134
rect 338430 252996 338436 253060
rect 338500 253058 338506 253060
rect 339401 253058 339467 253061
rect 338500 253056 339467 253058
rect 338500 253000 339406 253056
rect 339462 253000 339467 253056
rect 338500 252998 339467 253000
rect 338500 252996 338506 252998
rect 339401 252995 339467 252998
rect 498510 252724 498516 252788
rect 498580 252786 498586 252788
rect 499205 252786 499271 252789
rect 498580 252784 499271 252786
rect 498580 252728 499210 252784
rect 499266 252728 499271 252784
rect 498580 252726 499271 252728
rect 498580 252724 498586 252726
rect 499205 252723 499271 252726
rect 510889 252652 510955 252653
rect 510838 252650 510844 252652
rect 510798 252590 510844 252650
rect 510908 252648 510955 252652
rect 510950 252592 510955 252648
rect 510838 252588 510844 252590
rect 510908 252588 510955 252592
rect 510889 252587 510955 252588
rect 56685 252514 56751 252517
rect 57462 252514 57468 252516
rect 56685 252512 57468 252514
rect 56685 252456 56690 252512
rect 56746 252456 57468 252512
rect 56685 252454 57468 252456
rect 56685 252451 56751 252454
rect 57462 252452 57468 252454
rect 57532 252452 57538 252516
rect 57278 252316 57284 252380
rect 57348 252378 57354 252380
rect 60917 252378 60983 252381
rect 57348 252376 60983 252378
rect 57348 252320 60922 252376
rect 60978 252320 60983 252376
rect 57348 252318 60983 252320
rect 57348 252316 57354 252318
rect 60917 252315 60983 252318
rect 217542 251772 217548 251836
rect 217612 251834 217618 251836
rect 231853 251834 231919 251837
rect 217612 251832 231919 251834
rect 217612 251776 231858 251832
rect 231914 251776 231919 251832
rect 217612 251774 231919 251776
rect 217612 251772 217618 251774
rect 231853 251771 231919 251774
rect 377990 251772 377996 251836
rect 378060 251834 378066 251836
rect 396717 251834 396783 251837
rect 378060 251832 396783 251834
rect 378060 251776 396722 251832
rect 396778 251776 396783 251832
rect 378060 251774 396783 251776
rect 378060 251772 378066 251774
rect 396717 251771 396783 251774
rect 46790 251092 46796 251156
rect 46860 251154 46866 251156
rect 58617 251154 58683 251157
rect 46860 251152 58683 251154
rect 46860 251096 58622 251152
rect 58678 251096 58683 251152
rect 46860 251094 58683 251096
rect 46860 251092 46866 251094
rect 58617 251091 58683 251094
rect 198825 246258 198891 246261
rect 358905 246258 358971 246261
rect 519261 246258 519327 246261
rect 196558 246256 198891 246258
rect 196558 246200 198830 246256
rect 198886 246200 198891 246256
rect 196558 246198 198891 246200
rect 196558 246190 196618 246198
rect 198825 246195 198891 246198
rect 356562 246256 358971 246258
rect 356562 246200 358910 246256
rect 358966 246200 358971 246256
rect 356562 246198 358971 246200
rect 356562 246190 356622 246198
rect 358905 246195 358971 246198
rect 516558 246256 519327 246258
rect 516558 246200 519266 246256
rect 519322 246200 519327 246256
rect 516558 246198 519327 246200
rect 516558 246190 516618 246198
rect 519261 246195 519327 246198
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 57145 204234 57211 204237
rect 57513 204234 57579 204237
rect 376753 204234 376819 204237
rect 377213 204234 377279 204237
rect 57145 204232 60062 204234
rect 57145 204176 57150 204232
rect 57206 204176 57518 204232
rect 57574 204176 60062 204232
rect 57145 204174 60062 204176
rect 57145 204171 57211 204174
rect 57513 204171 57579 204174
rect 60002 203894 60062 204174
rect 376753 204232 377279 204234
rect 376753 204176 376758 204232
rect 376814 204176 377218 204232
rect 377274 204176 377279 204232
rect 376753 204174 377279 204176
rect 376753 204171 376819 204174
rect 377213 204171 377279 204174
rect 216857 203962 216923 203965
rect 217501 203962 217567 203965
rect 376937 203962 377003 203965
rect 216857 203960 219450 203962
rect 216857 203904 216862 203960
rect 216918 203904 217506 203960
rect 217562 203924 219450 203960
rect 376937 203960 379530 203962
rect 217562 203904 220064 203924
rect 216857 203902 220064 203904
rect 216857 203899 216923 203902
rect 217501 203899 217567 203902
rect 219390 203864 220064 203902
rect 376937 203904 376942 203960
rect 376998 203924 379530 203960
rect 376998 203904 380052 203924
rect 376937 203902 380052 203904
rect 376937 203899 377003 203902
rect 379470 203864 380052 203902
rect 56593 203010 56659 203013
rect 216949 203010 217015 203013
rect 376753 203010 376819 203013
rect 56593 203008 60062 203010
rect 56593 202952 56598 203008
rect 56654 202952 60062 203008
rect 56593 202950 60062 202952
rect 56593 202947 56659 202950
rect 60002 202942 60062 202950
rect 216949 203008 219450 203010
rect 216949 202952 216954 203008
rect 217010 202972 219450 203008
rect 376753 203008 379530 203010
rect 217010 202952 220064 202972
rect 216949 202950 220064 202952
rect 216949 202947 217015 202950
rect 219390 202912 220064 202950
rect 376753 202952 376758 203008
rect 376814 202972 379530 203008
rect 376814 202952 380052 202972
rect 376753 202950 380052 202952
rect 376753 202947 376819 202950
rect 379470 202912 380052 202950
rect -960 201922 480 202012
rect -960 201862 6930 201922
rect -960 201772 480 201862
rect 6870 201514 6930 201862
rect 51574 201514 51580 201516
rect 6870 201454 51580 201514
rect 51574 201452 51580 201454
rect 51644 201452 51650 201516
rect 56777 201378 56843 201381
rect 57881 201378 57947 201381
rect 376845 201378 376911 201381
rect 377673 201378 377739 201381
rect 56777 201376 60062 201378
rect 56777 201320 56782 201376
rect 56838 201320 57886 201376
rect 57942 201320 60062 201376
rect 56777 201318 60062 201320
rect 56777 201315 56843 201318
rect 57881 201315 57947 201318
rect 60002 200766 60062 201318
rect 376845 201376 377739 201378
rect 376845 201320 376850 201376
rect 376906 201320 377678 201376
rect 377734 201320 377739 201376
rect 376845 201318 377739 201320
rect 376845 201315 376911 201318
rect 377673 201315 377739 201318
rect 217685 200834 217751 200837
rect 377673 200834 377739 200837
rect 217685 200832 219450 200834
rect 217685 200776 217690 200832
rect 217746 200796 219450 200832
rect 377673 200832 379530 200834
rect 217746 200776 220064 200796
rect 217685 200774 220064 200776
rect 217685 200771 217751 200774
rect 219390 200736 220064 200774
rect 377673 200776 377678 200832
rect 377734 200796 379530 200832
rect 377734 200776 380052 200796
rect 377673 200774 380052 200776
rect 377673 200771 377739 200774
rect 379470 200736 380052 200774
rect 57697 199882 57763 199885
rect 217409 199882 217475 199885
rect 377949 199882 378015 199885
rect 57697 199880 60062 199882
rect 57697 199824 57702 199880
rect 57758 199824 60062 199880
rect 57697 199822 60062 199824
rect 57697 199819 57763 199822
rect 60002 199814 60062 199822
rect 217409 199880 219450 199882
rect 217409 199824 217414 199880
rect 217470 199844 219450 199880
rect 377949 199880 379530 199882
rect 217470 199824 220064 199844
rect 217409 199822 220064 199824
rect 217409 199819 217475 199822
rect 219390 199784 220064 199822
rect 377949 199824 377954 199880
rect 378010 199844 379530 199880
rect 378010 199824 380052 199844
rect 377949 199822 380052 199824
rect 377949 199819 378015 199822
rect 379470 199784 380052 199822
rect 57329 198794 57395 198797
rect 57697 198794 57763 198797
rect 57329 198792 57763 198794
rect 57329 198736 57334 198792
rect 57390 198736 57702 198792
rect 57758 198736 57763 198792
rect 57329 198734 57763 198736
rect 57329 198731 57395 198734
rect 57697 198731 57763 198734
rect 376937 198794 377003 198797
rect 377949 198794 378015 198797
rect 376937 198792 378015 198794
rect 376937 198736 376942 198792
rect 376998 198736 377954 198792
rect 378010 198736 378015 198792
rect 376937 198734 378015 198736
rect 376937 198731 377003 198734
rect 377949 198731 378015 198734
rect 57789 198114 57855 198117
rect 217777 198114 217843 198117
rect 377581 198114 377647 198117
rect 57789 198112 60062 198114
rect 57789 198056 57794 198112
rect 57850 198056 60062 198112
rect 57789 198054 60062 198056
rect 57789 198051 57855 198054
rect 60002 198046 60062 198054
rect 217777 198112 219450 198114
rect 217777 198056 217782 198112
rect 217838 198076 219450 198112
rect 377581 198112 379530 198114
rect 217838 198056 220064 198076
rect 217777 198054 220064 198056
rect 217777 198051 217843 198054
rect 219390 198016 220064 198054
rect 377581 198056 377586 198112
rect 377642 198076 379530 198112
rect 377642 198056 380052 198076
rect 377581 198054 380052 198056
rect 377581 198051 377647 198054
rect 379470 198016 380052 198054
rect 217501 197434 217567 197437
rect 217777 197434 217843 197437
rect 217501 197432 217843 197434
rect 217501 197376 217506 197432
rect 217562 197376 217782 197432
rect 217838 197376 217843 197432
rect 217501 197374 217843 197376
rect 217501 197371 217567 197374
rect 217777 197371 217843 197374
rect 217225 197026 217291 197029
rect 217593 197026 217659 197029
rect 377305 197026 377371 197029
rect 377857 197026 377923 197029
rect 217225 197024 219450 197026
rect 217225 196968 217230 197024
rect 217286 196968 217598 197024
rect 217654 196988 219450 197024
rect 377305 197024 379530 197026
rect 217654 196968 220064 196988
rect 217225 196966 220064 196968
rect 217225 196963 217291 196966
rect 217593 196963 217659 196966
rect 57421 196346 57487 196349
rect 60002 196346 60062 196958
rect 219390 196928 220064 196966
rect 377305 196968 377310 197024
rect 377366 196968 377862 197024
rect 377918 196988 379530 197024
rect 377918 196968 380052 196988
rect 377305 196966 380052 196968
rect 377305 196963 377371 196966
rect 377857 196963 377923 196966
rect 379470 196928 380052 196966
rect 57421 196344 60062 196346
rect 57421 196288 57426 196344
rect 57482 196288 60062 196344
rect 57421 196286 60062 196288
rect 57421 196283 57487 196286
rect 56961 195258 57027 195261
rect 57789 195258 57855 195261
rect 217133 195258 217199 195261
rect 217593 195258 217659 195261
rect 377397 195258 377463 195261
rect 377949 195258 378015 195261
rect 56961 195256 60062 195258
rect 56961 195200 56966 195256
rect 57022 195200 57794 195256
rect 57850 195200 60062 195256
rect 56961 195198 60062 195200
rect 56961 195195 57027 195198
rect 57789 195195 57855 195198
rect 60002 195190 60062 195198
rect 217133 195256 219450 195258
rect 217133 195200 217138 195256
rect 217194 195200 217598 195256
rect 217654 195220 219450 195256
rect 377397 195256 379530 195258
rect 217654 195200 220064 195220
rect 217133 195198 220064 195200
rect 217133 195195 217199 195198
rect 217593 195195 217659 195198
rect 219390 195160 220064 195198
rect 377397 195200 377402 195256
rect 377458 195200 377954 195256
rect 378010 195220 379530 195256
rect 378010 195200 380052 195220
rect 377397 195198 380052 195200
rect 377397 195195 377463 195198
rect 377949 195195 378015 195198
rect 379470 195160 380052 195198
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 199377 186418 199443 186421
rect 359365 186418 359431 186421
rect 518893 186418 518959 186421
rect 519353 186418 519419 186421
rect 196558 186416 199443 186418
rect 196558 186360 199382 186416
rect 199438 186360 199443 186416
rect 196558 186358 199443 186360
rect 196558 186350 196618 186358
rect 199377 186355 199443 186358
rect 356562 186416 359431 186418
rect 356562 186360 359370 186416
rect 359426 186360 359431 186416
rect 356562 186358 359431 186360
rect 356562 186350 356622 186358
rect 359365 186355 359431 186358
rect 516558 186416 519419 186418
rect 516558 186360 518898 186416
rect 518954 186360 519358 186416
rect 519414 186360 519419 186416
rect 516558 186358 519419 186360
rect 516558 186350 516618 186358
rect 518893 186355 518959 186358
rect 519353 186355 519419 186358
rect 198733 184922 198799 184925
rect 199285 184922 199351 184925
rect 359089 184922 359155 184925
rect 196558 184920 199351 184922
rect 196558 184864 198738 184920
rect 198794 184864 199290 184920
rect 199346 184864 199351 184920
rect 196558 184862 199351 184864
rect 196558 184718 196618 184862
rect 198733 184859 198799 184862
rect 199285 184859 199351 184862
rect 356562 184920 359155 184922
rect 356562 184864 359094 184920
rect 359150 184864 359155 184920
rect 356562 184862 359155 184864
rect 356562 184718 356622 184862
rect 359089 184859 359155 184862
rect 519537 184786 519603 184789
rect 520181 184786 520247 184789
rect 516558 184784 520247 184786
rect 516558 184728 519542 184784
rect 519598 184728 520186 184784
rect 520242 184728 520247 184784
rect 516558 184726 520247 184728
rect 516558 184718 516618 184726
rect 519537 184723 519603 184726
rect 520181 184723 520247 184726
rect 359273 183562 359339 183565
rect 359549 183562 359615 183565
rect 356562 183560 359615 183562
rect 356562 183504 359278 183560
rect 359334 183504 359554 183560
rect 359610 183504 359615 183560
rect 356562 183502 359615 183504
rect 199101 183426 199167 183429
rect 196558 183424 199167 183426
rect 196558 183368 199106 183424
rect 199162 183368 199167 183424
rect 196558 183366 199167 183368
rect 196558 183358 196618 183366
rect 199101 183363 199167 183366
rect 356562 183358 356622 183502
rect 359273 183499 359339 183502
rect 359549 183499 359615 183502
rect 519077 183426 519143 183429
rect 520089 183426 520155 183429
rect 516558 183424 520155 183426
rect 516558 183368 519082 183424
rect 519138 183368 520094 183424
rect 520150 183368 520155 183424
rect 516558 183366 520155 183368
rect 516558 183358 516618 183366
rect 519077 183363 519143 183366
rect 520089 183363 520155 183366
rect 198733 182066 198799 182069
rect 198917 182066 198983 182069
rect 358813 182066 358879 182069
rect 359181 182066 359247 182069
rect 196558 182064 198983 182066
rect 196558 182008 198738 182064
rect 198794 182008 198922 182064
rect 198978 182008 198983 182064
rect 196558 182006 198983 182008
rect 196558 181862 196618 182006
rect 198733 182003 198799 182006
rect 198917 182003 198983 182006
rect 356562 182064 359247 182066
rect 356562 182008 358818 182064
rect 358874 182008 359186 182064
rect 359242 182008 359247 182064
rect 356562 182006 359247 182008
rect 356562 181862 356622 182006
rect 358813 182003 358879 182006
rect 359181 182003 359247 182006
rect 519169 181930 519235 181933
rect 519353 181930 519419 181933
rect 516558 181928 519419 181930
rect 516558 181872 519174 181928
rect 519230 181872 519358 181928
rect 519414 181872 519419 181928
rect 516558 181870 519419 181872
rect 516558 181862 516618 181870
rect 519169 181867 519235 181870
rect 519353 181867 519419 181870
rect 199009 180706 199075 180709
rect 358997 180706 359063 180709
rect 518985 180706 519051 180709
rect 196558 180704 199075 180706
rect 196558 180648 199014 180704
rect 199070 180648 199075 180704
rect 196558 180646 199075 180648
rect 196558 180638 196618 180646
rect 199009 180643 199075 180646
rect 356562 180704 359063 180706
rect 356562 180648 359002 180704
rect 359058 180648 359063 180704
rect 356562 180646 359063 180648
rect 356562 180638 356622 180646
rect 358997 180643 359063 180646
rect 516558 180704 519051 180706
rect 516558 180648 518990 180704
rect 519046 180648 519051 180704
rect 516558 180646 519051 180648
rect 516558 180638 516618 180646
rect 518985 180643 519051 180646
rect 199009 179482 199075 179485
rect 199193 179482 199259 179485
rect 199009 179480 199259 179482
rect 199009 179424 199014 179480
rect 199070 179424 199198 179480
rect 199254 179424 199259 179480
rect 199009 179422 199259 179424
rect 199009 179419 199075 179422
rect 199193 179419 199259 179422
rect 583520 179060 584960 179300
rect 59077 177578 59143 177581
rect 59077 177576 60062 177578
rect 59077 177520 59082 177576
rect 59138 177520 60062 177576
rect 59077 177518 60062 177520
rect 59077 177515 59143 177518
rect 60002 176966 60062 177518
rect 217041 177034 217107 177037
rect 377029 177034 377095 177037
rect 217041 177032 219450 177034
rect 217041 176976 217046 177032
rect 217102 176996 219450 177032
rect 377029 177032 379530 177034
rect 217102 176976 220064 176996
rect 217041 176974 220064 176976
rect 217041 176971 217107 176974
rect 219390 176936 220064 176974
rect 377029 176976 377034 177032
rect 377090 176996 379530 177032
rect 377090 176976 380052 176996
rect 377029 176974 380052 176976
rect 377029 176971 377095 176974
rect 379470 176936 380052 176974
rect -960 175796 480 176036
rect 57237 175402 57303 175405
rect 57881 175402 57947 175405
rect 216673 175402 216739 175405
rect 376937 175402 377003 175405
rect 57237 175400 60062 175402
rect 57237 175344 57242 175400
rect 57298 175344 57886 175400
rect 57942 175344 60062 175400
rect 57237 175342 60062 175344
rect 57237 175339 57303 175342
rect 57881 175339 57947 175342
rect 60002 175334 60062 175342
rect 216673 175400 219450 175402
rect 216673 175344 216678 175400
rect 216734 175364 219450 175400
rect 376937 175400 379530 175402
rect 216734 175344 220064 175364
rect 216673 175342 220064 175344
rect 216673 175339 216739 175342
rect 219390 175304 220064 175342
rect 376937 175344 376942 175400
rect 376998 175364 379530 175400
rect 376998 175344 380052 175364
rect 376937 175342 380052 175344
rect 376937 175339 377003 175342
rect 379470 175304 380052 175342
rect 57646 175068 57652 175132
rect 57716 175130 57722 175132
rect 217133 175130 217199 175133
rect 377397 175130 377463 175133
rect 57716 175092 59554 175130
rect 217133 175128 219450 175130
rect 57716 175070 60032 175092
rect 57716 175068 57722 175070
rect 59494 175032 60032 175070
rect 217133 175072 217138 175128
rect 217194 175092 219450 175128
rect 377397 175128 379530 175130
rect 217194 175072 220064 175092
rect 217133 175070 220064 175072
rect 217133 175067 217199 175070
rect 219390 175032 220064 175070
rect 377397 175072 377402 175128
rect 377458 175092 379530 175128
rect 377458 175072 380052 175092
rect 377397 175070 380052 175072
rect 377397 175067 377463 175070
rect 379470 175032 380052 175070
rect 57830 166908 57836 166972
rect 57900 166970 57906 166972
rect 57900 166910 143572 166970
rect 57900 166908 57906 166910
rect 101029 166836 101095 166837
rect 103513 166836 103579 166837
rect 108297 166836 108363 166837
rect 138473 166836 138539 166837
rect 140865 166836 140931 166837
rect 143512 166836 143572 166910
rect 198222 166908 198228 166972
rect 198292 166970 198298 166972
rect 198292 166910 313500 166970
rect 198292 166908 198298 166910
rect 145925 166836 145991 166837
rect 313440 166836 313500 166910
rect 418429 166836 418495 166837
rect 421005 166836 421071 166837
rect 423397 166836 423463 166837
rect 445845 166836 445911 166837
rect 470961 166836 471027 166837
rect 473445 166836 473511 166837
rect 101029 166832 101078 166836
rect 101142 166834 101148 166836
rect 101029 166776 101034 166832
rect 101029 166772 101078 166776
rect 101142 166774 101186 166834
rect 103513 166832 103526 166836
rect 103590 166834 103596 166836
rect 108280 166834 108286 166836
rect 103513 166776 103518 166832
rect 101142 166772 101148 166774
rect 103513 166772 103526 166776
rect 103590 166774 103670 166834
rect 108206 166774 108286 166834
rect 108350 166832 108363 166836
rect 108358 166776 108363 166832
rect 103590 166772 103596 166774
rect 108280 166772 108286 166774
rect 108350 166772 108363 166776
rect 138472 166772 138478 166836
rect 138542 166834 138548 166836
rect 138542 166774 138630 166834
rect 140865 166832 140926 166836
rect 140865 166776 140870 166832
rect 138542 166772 138548 166774
rect 140865 166772 140926 166776
rect 140990 166834 140996 166836
rect 140990 166774 141022 166834
rect 140990 166772 140996 166774
rect 143504 166772 143510 166836
rect 143574 166772 143580 166836
rect 145925 166832 145958 166836
rect 146022 166834 146028 166836
rect 145925 166776 145930 166832
rect 145925 166772 145958 166776
rect 146022 166774 146082 166834
rect 146022 166772 146028 166774
rect 213494 166772 213500 166836
rect 213564 166834 213570 166836
rect 303504 166834 303510 166836
rect 213564 166774 303510 166834
rect 213564 166772 213570 166774
rect 303504 166772 303510 166774
rect 303574 166772 303580 166836
rect 313432 166772 313438 166836
rect 313502 166772 313508 166836
rect 418429 166834 418476 166836
rect 418384 166832 418476 166834
rect 418384 166776 418434 166832
rect 418384 166774 418476 166776
rect 418429 166772 418476 166774
rect 418540 166772 418546 166836
rect 421005 166834 421052 166836
rect 420960 166832 421052 166834
rect 420960 166776 421010 166832
rect 420960 166774 421052 166776
rect 421005 166772 421052 166774
rect 421116 166772 421122 166836
rect 423397 166834 423444 166836
rect 423352 166832 423444 166834
rect 423352 166776 423402 166832
rect 423352 166774 423444 166776
rect 423397 166772 423444 166774
rect 423508 166772 423514 166836
rect 445845 166834 445892 166836
rect 445800 166832 445892 166834
rect 445800 166776 445850 166832
rect 445800 166774 445892 166776
rect 445845 166772 445892 166774
rect 445956 166772 445962 166836
rect 470961 166832 470990 166836
rect 471054 166834 471060 166836
rect 473432 166834 473438 166836
rect 470961 166776 470966 166832
rect 470961 166772 470990 166776
rect 471054 166774 471118 166834
rect 473354 166774 473438 166834
rect 473502 166832 473511 166836
rect 473506 166776 473511 166832
rect 471054 166772 471060 166774
rect 473432 166772 473438 166774
rect 473502 166772 473511 166776
rect 101029 166771 101095 166772
rect 103513 166771 103579 166772
rect 108297 166771 108363 166772
rect 138473 166771 138539 166772
rect 140865 166771 140931 166772
rect 145925 166771 145991 166772
rect 418429 166771 418495 166772
rect 421005 166771 421071 166772
rect 423397 166771 423463 166772
rect 445845 166771 445911 166772
rect 470961 166771 471027 166772
rect 473445 166771 473511 166772
rect 475837 166836 475903 166837
rect 478413 166836 478479 166837
rect 480897 166836 480963 166837
rect 475837 166832 475886 166836
rect 475950 166834 475956 166836
rect 475837 166776 475842 166832
rect 475837 166772 475886 166776
rect 475950 166774 475994 166834
rect 478413 166832 478470 166836
rect 478534 166834 478540 166836
rect 478413 166776 478418 166832
rect 475950 166772 475956 166774
rect 478413 166772 478470 166776
rect 478534 166774 478570 166834
rect 480897 166832 480918 166836
rect 480982 166834 480988 166836
rect 480897 166776 480902 166832
rect 478534 166772 478540 166774
rect 480897 166772 480918 166776
rect 480982 166774 481054 166834
rect 480982 166772 480988 166774
rect 475837 166771 475903 166772
rect 478413 166771 478479 166772
rect 480897 166771 480963 166772
rect 148501 166700 148567 166701
rect 163313 166700 163379 166701
rect 165889 166700 165955 166701
rect 285949 166700 286015 166701
rect 291009 166700 291075 166701
rect 148501 166698 148548 166700
rect 148456 166696 148548 166698
rect 148456 166640 148506 166696
rect 148456 166638 148548 166640
rect 148501 166636 148548 166638
rect 148612 166636 148618 166700
rect 163313 166696 163366 166700
rect 163430 166698 163436 166700
rect 163313 166640 163318 166696
rect 163313 166636 163366 166640
rect 163430 166638 163470 166698
rect 165889 166696 165950 166700
rect 165889 166640 165894 166696
rect 163430 166636 163436 166638
rect 165889 166636 165950 166640
rect 166014 166698 166020 166700
rect 166014 166638 166046 166698
rect 166014 166636 166020 166638
rect 205214 166636 205220 166700
rect 205284 166698 205290 166700
rect 205284 166638 273270 166698
rect 205284 166636 205290 166638
rect 148501 166635 148567 166636
rect 163313 166635 163379 166636
rect 165889 166635 165955 166636
rect 107653 166564 107719 166565
rect 107600 166562 107606 166564
rect 107562 166502 107606 166562
rect 107670 166560 107719 166564
rect 150893 166564 150959 166565
rect 153285 166564 153351 166565
rect 183277 166564 183343 166565
rect 150893 166562 150940 166564
rect 107714 166504 107719 166560
rect 107600 166500 107606 166502
rect 107670 166500 107719 166504
rect 150848 166560 150940 166562
rect 150848 166504 150898 166560
rect 150848 166502 150940 166504
rect 107653 166499 107719 166500
rect 150893 166500 150940 166502
rect 151004 166500 151010 166564
rect 153285 166562 153332 166564
rect 153240 166560 153332 166562
rect 153240 166504 153290 166560
rect 153240 166502 153332 166504
rect 153285 166500 153332 166502
rect 153396 166500 153402 166564
rect 183216 166562 183222 166564
rect 183186 166502 183222 166562
rect 183286 166560 183343 166564
rect 260925 166564 260991 166565
rect 265893 166564 265959 166565
rect 270861 166564 270927 166565
rect 260925 166562 260972 166564
rect 183338 166504 183343 166560
rect 183216 166500 183222 166502
rect 183286 166500 183343 166504
rect 260880 166560 260972 166562
rect 260880 166504 260930 166560
rect 260880 166502 260972 166504
rect 150893 166499 150959 166500
rect 153285 166499 153351 166500
rect 183277 166499 183343 166500
rect 260925 166500 260972 166502
rect 261036 166500 261042 166564
rect 265893 166562 265940 166564
rect 265848 166560 265940 166562
rect 265848 166504 265898 166560
rect 265848 166502 265940 166504
rect 265893 166500 265940 166502
rect 266004 166500 266010 166564
rect 270861 166562 270908 166564
rect 270816 166560 270908 166562
rect 270816 166504 270866 166560
rect 270816 166502 270908 166504
rect 270861 166500 270908 166502
rect 270972 166500 270978 166564
rect 273210 166562 273270 166638
rect 285949 166696 285966 166700
rect 286030 166698 286036 166700
rect 290992 166698 290998 166700
rect 285949 166640 285954 166696
rect 285949 166636 285966 166640
rect 286030 166638 286106 166698
rect 290918 166638 290998 166698
rect 291062 166696 291075 166700
rect 291070 166640 291075 166696
rect 286030 166636 286036 166638
rect 290992 166636 290998 166638
rect 291062 166636 291075 166640
rect 285949 166635 286015 166636
rect 291009 166635 291075 166636
rect 293401 166700 293467 166701
rect 295885 166700 295951 166701
rect 298461 166700 298527 166701
rect 305913 166700 305979 166701
rect 483381 166700 483447 166701
rect 485957 166700 486023 166701
rect 293401 166696 293446 166700
rect 293510 166698 293516 166700
rect 293401 166640 293406 166696
rect 293401 166636 293446 166640
rect 293510 166638 293558 166698
rect 295885 166696 295894 166700
rect 295958 166698 295964 166700
rect 295885 166640 295890 166696
rect 293510 166636 293516 166638
rect 295885 166636 295894 166640
rect 295958 166638 296042 166698
rect 298461 166696 298478 166700
rect 298542 166698 298548 166700
rect 298461 166640 298466 166696
rect 295958 166636 295964 166638
rect 298461 166636 298478 166640
rect 298542 166638 298618 166698
rect 305913 166696 305958 166700
rect 306022 166698 306028 166700
rect 483360 166698 483366 166700
rect 305913 166640 305918 166696
rect 298542 166636 298548 166638
rect 305913 166636 305958 166640
rect 306022 166638 306070 166698
rect 483290 166638 483366 166698
rect 483430 166696 483447 166700
rect 485944 166698 485950 166700
rect 483442 166640 483447 166696
rect 306022 166636 306028 166638
rect 483360 166636 483366 166638
rect 483430 166636 483447 166640
rect 485866 166638 485950 166698
rect 486014 166696 486023 166700
rect 486018 166640 486023 166696
rect 485944 166636 485950 166638
rect 486014 166636 486023 166640
rect 293401 166635 293467 166636
rect 295885 166635 295951 166636
rect 298461 166635 298527 166636
rect 305913 166635 305979 166636
rect 483381 166635 483447 166636
rect 485957 166635 486023 166636
rect 503253 166564 503319 166565
rect 288272 166562 288278 166564
rect 273210 166502 288278 166562
rect 288272 166500 288278 166502
rect 288342 166500 288348 166564
rect 503216 166562 503222 166564
rect 503162 166502 503222 166562
rect 503286 166560 503319 166564
rect 503314 166504 503319 166560
rect 503216 166500 503222 166502
rect 503286 166500 503319 166504
rect 260925 166499 260991 166500
rect 265893 166499 265959 166500
rect 270861 166499 270927 166500
rect 503253 166499 503319 166500
rect 96061 166292 96127 166293
rect 98453 166292 98519 166293
rect 428181 166292 428247 166293
rect 430941 166292 431007 166293
rect 96061 166290 96108 166292
rect 96016 166288 96108 166290
rect 96016 166232 96066 166288
rect 96016 166230 96108 166232
rect 96061 166228 96108 166230
rect 96172 166228 96178 166292
rect 98453 166290 98500 166292
rect 98408 166288 98500 166290
rect 98408 166232 98458 166288
rect 98408 166230 98500 166232
rect 98453 166228 98500 166230
rect 98564 166228 98570 166292
rect 428181 166290 428228 166292
rect 428136 166288 428228 166290
rect 428136 166232 428186 166288
rect 428136 166230 428228 166232
rect 428181 166228 428228 166230
rect 428292 166228 428298 166292
rect 430941 166290 430988 166292
rect 430896 166288 430988 166290
rect 430896 166232 430946 166288
rect 430896 166230 430988 166232
rect 430941 166228 430988 166230
rect 431052 166228 431058 166292
rect 96061 166227 96127 166228
rect 98453 166227 98519 166228
rect 428181 166227 428247 166228
rect 430941 166227 431007 166228
rect 583520 165732 584960 165972
rect 81433 165610 81499 165613
rect 81750 165610 81756 165612
rect 81433 165608 81756 165610
rect 81433 165552 81438 165608
rect 81494 165552 81756 165608
rect 81433 165550 81756 165552
rect 81433 165547 81499 165550
rect 81750 165548 81756 165550
rect 81820 165548 81826 165612
rect 84285 165610 84351 165613
rect 85430 165610 85436 165612
rect 84285 165608 85436 165610
rect 84285 165552 84290 165608
rect 84346 165552 85436 165608
rect 84285 165550 85436 165552
rect 84285 165547 84351 165550
rect 85430 165548 85436 165550
rect 85500 165548 85506 165612
rect 91185 165610 91251 165613
rect 92422 165610 92428 165612
rect 91185 165608 92428 165610
rect 91185 165552 91190 165608
rect 91246 165552 92428 165608
rect 91185 165550 92428 165552
rect 91185 165547 91251 165550
rect 92422 165548 92428 165550
rect 92492 165548 92498 165612
rect 95233 165610 95299 165613
rect 99373 165612 99439 165613
rect 95734 165610 95740 165612
rect 95233 165608 95740 165610
rect 95233 165552 95238 165608
rect 95294 165552 95740 165608
rect 95233 165550 95740 165552
rect 95233 165547 95299 165550
rect 95734 165548 95740 165550
rect 95804 165548 95810 165612
rect 99373 165608 99420 165612
rect 99484 165610 99490 165612
rect 99373 165552 99378 165608
rect 99373 165548 99420 165552
rect 99484 165550 99530 165610
rect 99484 165548 99490 165550
rect 100702 165548 100708 165612
rect 100772 165610 100778 165612
rect 100845 165610 100911 165613
rect 100772 165608 100911 165610
rect 100772 165552 100850 165608
rect 100906 165552 100911 165608
rect 100772 165550 100911 165552
rect 100772 165548 100778 165550
rect 99373 165547 99439 165548
rect 100845 165547 100911 165550
rect 105169 165610 105235 165613
rect 105302 165610 105308 165612
rect 105169 165608 105308 165610
rect 105169 165552 105174 165608
rect 105230 165552 105308 165608
rect 105169 165550 105308 165552
rect 105169 165547 105235 165550
rect 105302 165548 105308 165550
rect 105372 165548 105378 165612
rect 105721 165610 105787 165613
rect 106365 165612 106431 165613
rect 105854 165610 105860 165612
rect 105721 165608 105860 165610
rect 105721 165552 105726 165608
rect 105782 165552 105860 165608
rect 105721 165550 105860 165552
rect 105721 165547 105787 165550
rect 105854 165548 105860 165550
rect 105924 165548 105930 165612
rect 106365 165608 106412 165612
rect 106476 165610 106482 165612
rect 108297 165610 108363 165613
rect 109677 165612 109743 165613
rect 110965 165612 111031 165613
rect 108614 165610 108620 165612
rect 106365 165552 106370 165608
rect 106365 165548 106412 165552
rect 106476 165550 106522 165610
rect 108297 165608 108620 165610
rect 108297 165552 108302 165608
rect 108358 165552 108620 165608
rect 108297 165550 108620 165552
rect 106476 165548 106482 165550
rect 106365 165547 106431 165548
rect 108297 165547 108363 165550
rect 108614 165548 108620 165550
rect 108684 165548 108690 165612
rect 109677 165608 109724 165612
rect 109788 165610 109794 165612
rect 109677 165552 109682 165608
rect 109677 165548 109724 165552
rect 109788 165550 109834 165610
rect 110965 165608 111012 165612
rect 111076 165610 111082 165612
rect 111885 165610 111951 165613
rect 113541 165612 113607 165613
rect 115933 165612 115999 165613
rect 112110 165610 112116 165612
rect 110965 165552 110970 165608
rect 109788 165548 109794 165550
rect 110965 165548 111012 165552
rect 111076 165550 111122 165610
rect 111885 165608 112116 165610
rect 111885 165552 111890 165608
rect 111946 165552 112116 165608
rect 111885 165550 112116 165552
rect 111076 165548 111082 165550
rect 109677 165547 109743 165548
rect 110965 165547 111031 165548
rect 111885 165547 111951 165550
rect 112110 165548 112116 165550
rect 112180 165548 112186 165612
rect 113541 165608 113588 165612
rect 113652 165610 113658 165612
rect 113541 165552 113546 165608
rect 113541 165548 113588 165552
rect 113652 165550 113698 165610
rect 115933 165608 115980 165612
rect 116044 165610 116050 165612
rect 117865 165610 117931 165613
rect 118325 165612 118391 165613
rect 119061 165612 119127 165613
rect 120901 165612 120967 165613
rect 123477 165612 123543 165613
rect 125869 165612 125935 165613
rect 117998 165610 118004 165612
rect 115933 165552 115938 165608
rect 113652 165548 113658 165550
rect 115933 165548 115980 165552
rect 116044 165550 116090 165610
rect 117865 165608 118004 165610
rect 117865 165552 117870 165608
rect 117926 165552 118004 165608
rect 117865 165550 118004 165552
rect 116044 165548 116050 165550
rect 113541 165547 113607 165548
rect 115933 165547 115999 165548
rect 117865 165547 117931 165550
rect 117998 165548 118004 165550
rect 118068 165548 118074 165612
rect 118325 165608 118372 165612
rect 118436 165610 118442 165612
rect 118325 165552 118330 165608
rect 118325 165548 118372 165552
rect 118436 165550 118482 165610
rect 119061 165608 119108 165612
rect 119172 165610 119178 165612
rect 119061 165552 119066 165608
rect 118436 165548 118442 165550
rect 119061 165548 119108 165552
rect 119172 165550 119218 165610
rect 120901 165608 120948 165612
rect 121012 165610 121018 165612
rect 120901 165552 120906 165608
rect 119172 165548 119178 165550
rect 120901 165548 120948 165552
rect 121012 165550 121058 165610
rect 123477 165608 123524 165612
rect 123588 165610 123594 165612
rect 123477 165552 123482 165608
rect 121012 165548 121018 165550
rect 123477 165548 123524 165552
rect 123588 165550 123634 165610
rect 125869 165608 125916 165612
rect 125980 165610 125986 165612
rect 128353 165610 128419 165613
rect 128486 165610 128492 165612
rect 125869 165552 125874 165608
rect 123588 165548 123594 165550
rect 125869 165548 125916 165552
rect 125980 165550 126026 165610
rect 128353 165608 128492 165610
rect 128353 165552 128358 165608
rect 128414 165552 128492 165608
rect 128353 165550 128492 165552
rect 125980 165548 125986 165550
rect 118325 165547 118391 165548
rect 119061 165547 119127 165548
rect 120901 165547 120967 165548
rect 123477 165547 123543 165548
rect 125869 165547 125935 165548
rect 128353 165547 128419 165550
rect 128486 165548 128492 165550
rect 128556 165548 128562 165612
rect 129733 165610 129799 165613
rect 130878 165610 130884 165612
rect 129733 165608 130884 165610
rect 129733 165552 129738 165608
rect 129794 165552 130884 165608
rect 129733 165550 130884 165552
rect 129733 165547 129799 165550
rect 130878 165548 130884 165550
rect 130948 165548 130954 165612
rect 132493 165610 132559 165613
rect 183369 165612 183435 165613
rect 235993 165612 236059 165613
rect 133454 165610 133460 165612
rect 132493 165608 133460 165610
rect 132493 165552 132498 165608
rect 132554 165552 133460 165608
rect 132493 165550 133460 165552
rect 132493 165547 132559 165550
rect 133454 165548 133460 165550
rect 133524 165548 133530 165612
rect 183318 165548 183324 165612
rect 183388 165610 183435 165612
rect 183388 165608 183480 165610
rect 183430 165552 183480 165608
rect 183388 165550 183480 165552
rect 183388 165548 183435 165550
rect 235942 165548 235948 165612
rect 236012 165610 236059 165612
rect 238753 165610 238819 165613
rect 239622 165610 239628 165612
rect 236012 165608 236104 165610
rect 236054 165552 236104 165608
rect 236012 165550 236104 165552
rect 238753 165608 239628 165610
rect 238753 165552 238758 165608
rect 238814 165552 239628 165608
rect 238753 165550 239628 165552
rect 236012 165548 236059 165550
rect 183369 165547 183435 165548
rect 235993 165547 236059 165548
rect 238753 165547 238819 165550
rect 239622 165548 239628 165550
rect 239692 165548 239698 165612
rect 242893 165610 242959 165613
rect 243118 165610 243124 165612
rect 242893 165608 243124 165610
rect 242893 165552 242898 165608
rect 242954 165552 243124 165608
rect 242893 165550 243124 165552
rect 242893 165547 242959 165550
rect 243118 165548 243124 165550
rect 243188 165548 243194 165612
rect 247033 165610 247099 165613
rect 247534 165610 247540 165612
rect 247033 165608 247540 165610
rect 247033 165552 247038 165608
rect 247094 165552 247540 165608
rect 247033 165550 247540 165552
rect 247033 165547 247099 165550
rect 247534 165548 247540 165550
rect 247604 165548 247610 165612
rect 247677 165610 247743 165613
rect 248270 165610 248276 165612
rect 247677 165608 248276 165610
rect 247677 165552 247682 165608
rect 247738 165552 248276 165608
rect 247677 165550 248276 165552
rect 247677 165547 247743 165550
rect 248270 165548 248276 165550
rect 248340 165548 248346 165612
rect 249793 165610 249859 165613
rect 250662 165610 250668 165612
rect 249793 165608 250668 165610
rect 249793 165552 249798 165608
rect 249854 165552 250668 165608
rect 249793 165550 250668 165552
rect 249793 165547 249859 165550
rect 250662 165548 250668 165550
rect 250732 165548 250738 165612
rect 252553 165610 252619 165613
rect 253606 165610 253612 165612
rect 252553 165608 253612 165610
rect 252553 165552 252558 165608
rect 252614 165552 253612 165608
rect 252553 165550 253612 165552
rect 252553 165547 252619 165550
rect 253606 165548 253612 165550
rect 253676 165548 253682 165612
rect 258073 165610 258139 165613
rect 258390 165610 258396 165612
rect 258073 165608 258396 165610
rect 258073 165552 258078 165608
rect 258134 165552 258396 165608
rect 258073 165550 258396 165552
rect 258073 165547 258139 165550
rect 258390 165548 258396 165550
rect 258460 165548 258466 165612
rect 260833 165610 260899 165613
rect 261702 165610 261708 165612
rect 260833 165608 261708 165610
rect 260833 165552 260838 165608
rect 260894 165552 261708 165608
rect 260833 165550 261708 165552
rect 260833 165547 260899 165550
rect 261702 165548 261708 165550
rect 261772 165548 261778 165612
rect 264973 165610 265039 165613
rect 265198 165610 265204 165612
rect 264973 165608 265204 165610
rect 264973 165552 264978 165608
rect 265034 165552 265204 165608
rect 264973 165550 265204 165552
rect 264973 165547 265039 165550
rect 265198 165548 265204 165550
rect 265268 165548 265274 165612
rect 266486 165548 266492 165612
rect 266556 165610 266562 165612
rect 267641 165610 267707 165613
rect 266556 165608 267707 165610
rect 266556 165552 267646 165608
rect 267702 165552 267707 165608
rect 266556 165550 267707 165552
rect 266556 165548 266562 165550
rect 267641 165547 267707 165550
rect 267917 165610 267983 165613
rect 268326 165610 268332 165612
rect 267917 165608 268332 165610
rect 267917 165552 267922 165608
rect 267978 165552 268332 165608
rect 267917 165550 268332 165552
rect 267917 165547 267983 165550
rect 268326 165548 268332 165550
rect 268396 165548 268402 165612
rect 280153 165610 280219 165613
rect 283373 165612 283439 165613
rect 300853 165612 300919 165613
rect 308397 165612 308463 165613
rect 280838 165610 280844 165612
rect 280153 165608 280844 165610
rect 280153 165552 280158 165608
rect 280214 165552 280844 165608
rect 280153 165550 280844 165552
rect 280153 165547 280219 165550
rect 280838 165548 280844 165550
rect 280908 165548 280914 165612
rect 283373 165608 283420 165612
rect 283484 165610 283490 165612
rect 283373 165552 283378 165608
rect 283373 165548 283420 165552
rect 283484 165550 283530 165610
rect 300853 165608 300900 165612
rect 300964 165610 300970 165612
rect 300853 165552 300858 165608
rect 283484 165548 283490 165550
rect 300853 165548 300900 165552
rect 300964 165550 301010 165610
rect 308397 165608 308444 165612
rect 308508 165610 308514 165612
rect 323025 165610 323091 165613
rect 325877 165612 325943 165613
rect 343265 165612 343331 165613
rect 343449 165612 343515 165613
rect 323342 165610 323348 165612
rect 308397 165552 308402 165608
rect 300964 165548 300970 165550
rect 308397 165548 308444 165552
rect 308508 165550 308554 165610
rect 323025 165608 323348 165610
rect 323025 165552 323030 165608
rect 323086 165552 323348 165608
rect 323025 165550 323348 165552
rect 308508 165548 308514 165550
rect 283373 165547 283439 165548
rect 300853 165547 300919 165548
rect 308397 165547 308463 165548
rect 323025 165547 323091 165550
rect 323342 165548 323348 165550
rect 323412 165548 323418 165612
rect 325877 165608 325924 165612
rect 325988 165610 325994 165612
rect 343214 165610 343220 165612
rect 325877 165552 325882 165608
rect 325877 165548 325924 165552
rect 325988 165550 326034 165610
rect 343174 165550 343220 165610
rect 343284 165608 343331 165612
rect 343326 165552 343331 165608
rect 325988 165548 325994 165550
rect 343214 165548 343220 165550
rect 343284 165548 343331 165552
rect 343398 165548 343404 165612
rect 343468 165610 343515 165612
rect 397453 165610 397519 165613
rect 398230 165610 398236 165612
rect 343468 165608 343560 165610
rect 343510 165552 343560 165608
rect 343468 165550 343560 165552
rect 397453 165608 398236 165610
rect 397453 165552 397458 165608
rect 397514 165552 398236 165608
rect 397453 165550 398236 165552
rect 343468 165548 343515 165550
rect 325877 165547 325943 165548
rect 343265 165547 343331 165548
rect 343449 165547 343515 165548
rect 397453 165547 397519 165550
rect 398230 165548 398236 165550
rect 398300 165548 398306 165612
rect 401593 165610 401659 165613
rect 401726 165610 401732 165612
rect 401593 165608 401732 165610
rect 401593 165552 401598 165608
rect 401654 165552 401732 165608
rect 401593 165550 401732 165552
rect 401593 165547 401659 165550
rect 401726 165548 401732 165550
rect 401796 165548 401802 165612
rect 404353 165610 404419 165613
rect 405406 165610 405412 165612
rect 404353 165608 405412 165610
rect 404353 165552 404358 165608
rect 404414 165552 405412 165608
rect 404353 165550 405412 165552
rect 404353 165547 404419 165550
rect 405406 165548 405412 165550
rect 405476 165548 405482 165612
rect 407113 165610 407179 165613
rect 408166 165610 408172 165612
rect 407113 165608 408172 165610
rect 407113 165552 407118 165608
rect 407174 165552 408172 165608
rect 407113 165550 408172 165552
rect 407113 165547 407179 165550
rect 408166 165548 408172 165550
rect 408236 165548 408242 165612
rect 409873 165610 409939 165613
rect 410742 165610 410748 165612
rect 409873 165608 410748 165610
rect 409873 165552 409878 165608
rect 409934 165552 410748 165608
rect 409873 165550 410748 165552
rect 409873 165547 409939 165550
rect 410742 165548 410748 165550
rect 410812 165548 410818 165612
rect 415393 165610 415459 165613
rect 416037 165612 416103 165613
rect 415894 165610 415900 165612
rect 415393 165608 415900 165610
rect 415393 165552 415398 165608
rect 415454 165552 415900 165608
rect 415393 165550 415900 165552
rect 415393 165547 415459 165550
rect 415894 165548 415900 165550
rect 415964 165548 415970 165612
rect 416037 165608 416084 165612
rect 416148 165610 416154 165612
rect 418613 165610 418679 165613
rect 419390 165610 419396 165612
rect 416037 165552 416042 165608
rect 416037 165548 416084 165552
rect 416148 165550 416194 165610
rect 418613 165608 419396 165610
rect 418613 165552 418618 165608
rect 418674 165552 419396 165608
rect 418613 165550 419396 165552
rect 416148 165548 416154 165550
rect 416037 165547 416103 165548
rect 418613 165547 418679 165550
rect 419390 165548 419396 165550
rect 419460 165548 419466 165612
rect 423673 165610 423739 165613
rect 423806 165610 423812 165612
rect 423673 165608 423812 165610
rect 423673 165552 423678 165608
rect 423734 165552 423812 165608
rect 423673 165550 423812 165552
rect 423673 165547 423739 165550
rect 423806 165548 423812 165550
rect 423876 165548 423882 165612
rect 426382 165548 426388 165612
rect 426452 165610 426458 165612
rect 427629 165610 427695 165613
rect 433333 165612 433399 165613
rect 433333 165610 433380 165612
rect 426452 165608 427695 165610
rect 426452 165552 427634 165608
rect 427690 165552 427695 165608
rect 426452 165550 427695 165552
rect 433288 165608 433380 165610
rect 433288 165552 433338 165608
rect 433288 165550 433380 165552
rect 426452 165548 426458 165550
rect 427629 165547 427695 165550
rect 433333 165548 433380 165550
rect 433444 165548 433450 165612
rect 433517 165610 433583 165613
rect 434294 165610 434300 165612
rect 433517 165608 434300 165610
rect 433517 165552 433522 165608
rect 433578 165552 434300 165608
rect 433517 165550 434300 165552
rect 433333 165547 433399 165548
rect 433517 165547 433583 165550
rect 434294 165548 434300 165550
rect 434364 165548 434370 165612
rect 434713 165610 434779 165613
rect 437749 165612 437815 165613
rect 435950 165610 435956 165612
rect 434713 165608 435956 165610
rect 434713 165552 434718 165608
rect 434774 165552 435956 165608
rect 434713 165550 435956 165552
rect 434713 165547 434779 165550
rect 435950 165548 435956 165550
rect 436020 165548 436026 165612
rect 437749 165610 437796 165612
rect 437704 165608 437796 165610
rect 437704 165552 437754 165608
rect 437704 165550 437796 165552
rect 437749 165548 437796 165550
rect 437860 165548 437866 165612
rect 438025 165610 438091 165613
rect 438526 165610 438532 165612
rect 438025 165608 438532 165610
rect 438025 165552 438030 165608
rect 438086 165552 438532 165608
rect 438025 165550 438532 165552
rect 437749 165547 437815 165548
rect 438025 165547 438091 165550
rect 438526 165548 438532 165550
rect 438596 165548 438602 165612
rect 442993 165610 443059 165613
rect 443494 165610 443500 165612
rect 442993 165608 443500 165610
rect 442993 165552 442998 165608
rect 443054 165552 443500 165608
rect 442993 165550 443500 165552
rect 442993 165547 443059 165550
rect 443494 165548 443500 165550
rect 443564 165548 443570 165612
rect 447317 165610 447383 165613
rect 448278 165610 448284 165612
rect 447317 165608 448284 165610
rect 447317 165552 447322 165608
rect 447378 165552 448284 165608
rect 447317 165550 448284 165552
rect 447317 165547 447383 165550
rect 448278 165548 448284 165550
rect 448348 165548 448354 165612
rect 449893 165610 449959 165613
rect 451038 165610 451044 165612
rect 449893 165608 451044 165610
rect 449893 165552 449898 165608
rect 449954 165552 451044 165608
rect 449893 165550 451044 165552
rect 449893 165547 449959 165550
rect 451038 165548 451044 165550
rect 451108 165548 451114 165612
rect 452653 165610 452719 165613
rect 453430 165610 453436 165612
rect 452653 165608 453436 165610
rect 452653 165552 452658 165608
rect 452714 165552 453436 165608
rect 452653 165550 453436 165552
rect 452653 165547 452719 165550
rect 453430 165548 453436 165550
rect 453500 165548 453506 165612
rect 455413 165610 455479 165613
rect 458357 165612 458423 165613
rect 503345 165612 503411 165613
rect 455822 165610 455828 165612
rect 455413 165608 455828 165610
rect 455413 165552 455418 165608
rect 455474 165552 455828 165608
rect 455413 165550 455828 165552
rect 455413 165547 455479 165550
rect 455822 165548 455828 165550
rect 455892 165548 455898 165612
rect 458357 165608 458404 165612
rect 458468 165610 458474 165612
rect 458357 165552 458362 165608
rect 458357 165548 458404 165552
rect 458468 165550 458514 165610
rect 458468 165548 458474 165550
rect 503294 165548 503300 165612
rect 503364 165610 503411 165612
rect 503364 165608 503456 165610
rect 503406 165552 503456 165608
rect 503364 165550 503456 165552
rect 503364 165548 503411 165550
rect 458357 165547 458423 165548
rect 503345 165547 503411 165548
rect 50613 165474 50679 165477
rect 155902 165474 155908 165476
rect 50613 165472 155908 165474
rect 50613 165416 50618 165472
rect 50674 165416 155908 165472
rect 50613 165414 155908 165416
rect 50613 165411 50679 165414
rect 155902 165412 155908 165414
rect 155972 165412 155978 165476
rect 213126 165412 213132 165476
rect 213196 165474 213202 165476
rect 320950 165474 320956 165476
rect 213196 165414 320956 165474
rect 213196 165412 213202 165414
rect 320950 165412 320956 165414
rect 321020 165412 321026 165476
rect 378777 165474 378843 165477
rect 468518 165474 468524 165476
rect 378777 165472 468524 165474
rect 378777 165416 378782 165472
rect 378838 165416 468524 165472
rect 378777 165414 468524 165416
rect 378777 165411 378843 165414
rect 468518 165412 468524 165414
rect 468588 165412 468594 165476
rect 53465 165338 53531 165341
rect 158478 165338 158484 165340
rect 53465 165336 158484 165338
rect 53465 165280 53470 165336
rect 53526 165280 158484 165336
rect 53465 165278 158484 165280
rect 53465 165275 53531 165278
rect 158478 165276 158484 165278
rect 158548 165276 158554 165340
rect 206134 165276 206140 165340
rect 206204 165338 206210 165340
rect 311014 165338 311020 165340
rect 206204 165278 311020 165338
rect 206204 165276 206210 165278
rect 311014 165276 311020 165278
rect 311084 165276 311090 165340
rect 376017 165338 376083 165341
rect 465942 165338 465948 165340
rect 376017 165336 465948 165338
rect 376017 165280 376022 165336
rect 376078 165280 465948 165336
rect 376017 165278 465948 165280
rect 376017 165275 376083 165278
rect 465942 165276 465948 165278
rect 466012 165276 466018 165340
rect 56133 165202 56199 165205
rect 135846 165202 135852 165204
rect 56133 165200 135852 165202
rect 56133 165144 56138 165200
rect 56194 165144 135852 165200
rect 56133 165142 135852 165144
rect 56133 165139 56199 165142
rect 135846 165140 135852 165142
rect 135916 165140 135922 165204
rect 213310 165140 213316 165204
rect 213380 165202 213386 165204
rect 271873 165202 271939 165205
rect 275921 165204 275987 165205
rect 272190 165202 272196 165204
rect 213380 165142 268578 165202
rect 213380 165140 213386 165142
rect 90265 165066 90331 165069
rect 113173 165068 113239 165069
rect 90766 165066 90772 165068
rect 90265 165064 90772 165066
rect 90265 165008 90270 165064
rect 90326 165008 90772 165064
rect 90265 165006 90772 165008
rect 90265 165003 90331 165006
rect 90766 165004 90772 165006
rect 90836 165004 90842 165068
rect 113173 165064 113220 165068
rect 113284 165066 113290 165068
rect 113173 165008 113178 165064
rect 113173 165004 113220 165008
rect 113284 165006 113330 165066
rect 113284 165004 113290 165006
rect 216254 165004 216260 165068
rect 216324 165066 216330 165068
rect 268518 165066 268578 165142
rect 271873 165200 272196 165202
rect 271873 165144 271878 165200
rect 271934 165144 272196 165200
rect 271873 165142 272196 165144
rect 271873 165139 271939 165142
rect 272190 165140 272196 165142
rect 272260 165140 272266 165204
rect 275870 165202 275876 165204
rect 275830 165142 275876 165202
rect 275940 165200 275987 165204
rect 275982 165144 275987 165200
rect 275870 165140 275876 165142
rect 275940 165140 275987 165144
rect 276054 165140 276060 165204
rect 276124 165140 276130 165204
rect 277393 165202 277459 165205
rect 278446 165202 278452 165204
rect 277393 165200 278452 165202
rect 277393 165144 277398 165200
rect 277454 165144 278452 165200
rect 277393 165142 278452 165144
rect 275921 165139 275987 165140
rect 273478 165066 273484 165068
rect 216324 165006 268394 165066
rect 268518 165006 273484 165066
rect 216324 165004 216330 165006
rect 113173 165003 113239 165004
rect 78673 164930 78739 164933
rect 88333 164932 88399 164933
rect 79542 164930 79548 164932
rect 78673 164928 79548 164930
rect 78673 164872 78678 164928
rect 78734 164872 79548 164928
rect 78673 164870 79548 164872
rect 78673 164867 78739 164870
rect 79542 164868 79548 164870
rect 79612 164868 79618 164932
rect 88333 164930 88380 164932
rect 88288 164928 88380 164930
rect 88288 164872 88338 164928
rect 88288 164870 88380 164872
rect 88333 164868 88380 164870
rect 88444 164868 88450 164932
rect 92473 164930 92539 164933
rect 114461 164932 114527 164933
rect 93710 164930 93716 164932
rect 92473 164928 93716 164930
rect 92473 164872 92478 164928
rect 92534 164872 93716 164928
rect 92473 164870 93716 164872
rect 88333 164867 88399 164868
rect 92473 164867 92539 164870
rect 93710 164868 93716 164870
rect 93780 164868 93786 164932
rect 114461 164928 114508 164932
rect 114572 164930 114578 164932
rect 114461 164872 114466 164928
rect 114461 164868 114508 164872
rect 114572 164870 114618 164930
rect 114572 164868 114578 164870
rect 207974 164868 207980 164932
rect 208044 164930 208050 164932
rect 263726 164930 263732 164932
rect 208044 164870 263732 164930
rect 208044 164868 208050 164870
rect 263726 164868 263732 164870
rect 263796 164868 263802 164932
rect 268334 164930 268394 165006
rect 273478 165004 273484 165006
rect 273548 165004 273554 165068
rect 276062 164930 276122 165140
rect 277393 165139 277459 165142
rect 278446 165140 278452 165142
rect 278516 165140 278522 165204
rect 279182 165140 279188 165204
rect 279252 165202 279258 165204
rect 280061 165202 280127 165205
rect 279252 165200 280127 165202
rect 279252 165144 280066 165200
rect 280122 165144 280127 165200
rect 279252 165142 280127 165144
rect 279252 165140 279258 165142
rect 280061 165139 280127 165142
rect 374862 165140 374868 165204
rect 374932 165202 374938 165204
rect 463550 165202 463556 165204
rect 374932 165142 463556 165202
rect 374932 165140 374938 165142
rect 463550 165140 463556 165142
rect 463620 165140 463626 165204
rect 379462 165004 379468 165068
rect 379532 165066 379538 165068
rect 426014 165066 426020 165068
rect 379532 165006 426020 165066
rect 379532 165004 379538 165006
rect 426014 165004 426020 165006
rect 426084 165004 426090 165068
rect 433333 165066 433399 165069
rect 433558 165066 433564 165068
rect 433333 165064 433564 165066
rect 433333 165008 433338 165064
rect 433394 165008 433564 165064
rect 433333 165006 433564 165008
rect 433333 165003 433399 165006
rect 433558 165004 433564 165006
rect 433628 165004 433634 165068
rect 268334 164870 276122 164930
rect 440325 164930 440391 164933
rect 440918 164930 440924 164932
rect 440325 164928 440924 164930
rect 440325 164872 440330 164928
rect 440386 164872 440924 164928
rect 440325 164870 440924 164872
rect 114461 164867 114527 164868
rect 440325 164867 440391 164870
rect 440918 164868 440924 164870
rect 440988 164868 440994 164932
rect 49417 164794 49483 164797
rect 160870 164794 160876 164796
rect 49417 164792 160876 164794
rect 49417 164736 49422 164792
rect 49478 164736 160876 164792
rect 49417 164734 160876 164736
rect 49417 164731 49483 164734
rect 160870 164732 160876 164734
rect 160940 164732 160946 164796
rect 200798 164732 200804 164796
rect 200868 164794 200874 164796
rect 256182 164794 256188 164796
rect 200868 164734 256188 164794
rect 200868 164732 200874 164734
rect 256182 164732 256188 164734
rect 256252 164732 256258 164796
rect 412633 164794 412699 164797
rect 413686 164794 413692 164796
rect 412633 164792 413692 164794
rect 412633 164736 412638 164792
rect 412694 164736 413692 164792
rect 412633 164734 413692 164736
rect 412633 164731 412699 164734
rect 413686 164732 413692 164734
rect 413756 164732 413762 164796
rect 420913 164794 420979 164797
rect 421782 164794 421788 164796
rect 420913 164792 421788 164794
rect 420913 164736 420918 164792
rect 420974 164736 421788 164792
rect 420913 164734 421788 164736
rect 420913 164731 420979 164734
rect 421782 164732 421788 164734
rect 421852 164732 421858 164796
rect 111149 164660 111215 164661
rect 111149 164656 111196 164660
rect 111260 164658 111266 164660
rect 366541 164658 366607 164661
rect 460974 164658 460980 164660
rect 111149 164600 111154 164656
rect 111149 164596 111196 164600
rect 111260 164598 111306 164658
rect 366541 164656 460980 164658
rect 366541 164600 366546 164656
rect 366602 164600 460980 164656
rect 366541 164598 460980 164600
rect 111260 164596 111266 164598
rect 111149 164595 111215 164596
rect 366541 164595 366607 164598
rect 460974 164596 460980 164598
rect 461044 164596 461050 164660
rect 115790 164460 115796 164524
rect 115860 164522 115866 164524
rect 115933 164522 115999 164525
rect 115860 164520 115999 164522
rect 115860 164464 115938 164520
rect 115994 164464 115999 164520
rect 115860 164462 115999 164464
rect 115860 164460 115866 164462
rect 115933 164459 115999 164462
rect 117078 164460 117084 164524
rect 117148 164522 117154 164524
rect 117313 164522 117379 164525
rect 117148 164520 117379 164522
rect 117148 164464 117318 164520
rect 117374 164464 117379 164520
rect 117148 164462 117379 164464
rect 117148 164460 117154 164462
rect 117313 164459 117379 164462
rect 244273 164522 244339 164525
rect 244406 164522 244412 164524
rect 244273 164520 244412 164522
rect 244273 164464 244278 164520
rect 244334 164464 244412 164520
rect 244273 164462 244412 164464
rect 244273 164459 244339 164462
rect 244406 164460 244412 164462
rect 244476 164460 244482 164524
rect 251265 164522 251331 164525
rect 252318 164522 252324 164524
rect 251265 164520 252324 164522
rect 251265 164464 251270 164520
rect 251326 164464 252324 164520
rect 251265 164462 252324 164464
rect 251265 164459 251331 164462
rect 252318 164460 252324 164462
rect 252388 164460 252394 164524
rect 259545 164522 259611 164525
rect 260598 164522 260604 164524
rect 259545 164520 260604 164522
rect 259545 164464 259550 164520
rect 259606 164464 260604 164520
rect 259545 164462 260604 164464
rect 259545 164459 259611 164462
rect 260598 164460 260604 164462
rect 260668 164460 260674 164524
rect 266353 164522 266419 164525
rect 267590 164522 267596 164524
rect 266353 164520 267596 164522
rect 266353 164464 266358 164520
rect 266414 164464 267596 164520
rect 266353 164462 267596 164464
rect 266353 164459 266419 164462
rect 267590 164460 267596 164462
rect 267660 164460 267666 164524
rect 273294 164460 273300 164524
rect 273364 164522 273370 164524
rect 274449 164522 274515 164525
rect 273364 164520 274515 164522
rect 273364 164464 274454 164520
rect 274510 164464 274515 164520
rect 273364 164462 274515 164464
rect 273364 164460 273370 164462
rect 274449 164459 274515 164462
rect 436093 164522 436159 164525
rect 436870 164522 436876 164524
rect 436093 164520 436876 164522
rect 436093 164464 436098 164520
rect 436154 164464 436876 164520
rect 436093 164462 436876 164464
rect 436093 164459 436159 164462
rect 436870 164460 436876 164462
rect 436940 164460 436946 164524
rect 76005 164386 76071 164389
rect 77150 164386 77156 164388
rect 76005 164384 77156 164386
rect 76005 164328 76010 164384
rect 76066 164328 77156 164384
rect 76005 164326 77156 164328
rect 76005 164323 76071 164326
rect 77150 164324 77156 164326
rect 77220 164324 77226 164388
rect 203006 164324 203012 164388
rect 203076 164386 203082 164388
rect 315062 164386 315068 164388
rect 203076 164326 315068 164386
rect 203076 164324 203082 164326
rect 315062 164324 315068 164326
rect 315132 164324 315138 164388
rect 396073 164386 396139 164389
rect 397126 164386 397132 164388
rect 396073 164384 397132 164386
rect 396073 164328 396078 164384
rect 396134 164328 397132 164384
rect 396073 164326 397132 164328
rect 396073 164323 396139 164326
rect 397126 164324 397132 164326
rect 397196 164324 397202 164388
rect 402973 164386 403039 164389
rect 404118 164386 404124 164388
rect 402973 164384 404124 164386
rect 402973 164328 402978 164384
rect 403034 164328 404124 164384
rect 402973 164326 404124 164328
rect 402973 164323 403039 164326
rect 404118 164324 404124 164326
rect 404188 164324 404194 164388
rect 411345 164386 411411 164389
rect 412398 164386 412404 164388
rect 411345 164384 412404 164386
rect 411345 164328 411350 164384
rect 411406 164328 412404 164384
rect 411345 164326 412404 164328
rect 411345 164323 411411 164326
rect 412398 164324 412404 164326
rect 412468 164324 412474 164388
rect 429285 164386 429351 164389
rect 429694 164386 429700 164388
rect 429285 164384 429700 164386
rect 429285 164328 429290 164384
rect 429346 164328 429700 164384
rect 429285 164326 429700 164328
rect 429285 164323 429351 164326
rect 429694 164324 429700 164326
rect 429764 164324 429770 164388
rect 57278 164188 57284 164252
rect 57348 164250 57354 164252
rect 59353 164250 59419 164253
rect 57348 164248 59419 164250
rect 57348 164192 59358 164248
rect 59414 164192 59419 164248
rect 57348 164190 59419 164192
rect 57348 164188 57354 164190
rect 59353 164187 59419 164190
rect 75913 164250 75979 164253
rect 76046 164250 76052 164252
rect 75913 164248 76052 164250
rect 75913 164192 75918 164248
rect 75974 164192 76052 164248
rect 75913 164190 76052 164192
rect 75913 164187 75979 164190
rect 76046 164188 76052 164190
rect 76116 164188 76122 164252
rect 77293 164250 77359 164253
rect 78254 164250 78260 164252
rect 77293 164248 78260 164250
rect 77293 164192 77298 164248
rect 77354 164192 78260 164248
rect 77293 164190 78260 164192
rect 77293 164187 77359 164190
rect 78254 164188 78260 164190
rect 78324 164188 78330 164252
rect 80053 164250 80119 164253
rect 80462 164250 80468 164252
rect 80053 164248 80468 164250
rect 80053 164192 80058 164248
rect 80114 164192 80468 164248
rect 80053 164190 80468 164192
rect 80053 164187 80119 164190
rect 80462 164188 80468 164190
rect 80532 164188 80538 164252
rect 82813 164250 82879 164253
rect 84193 164252 84259 164253
rect 83038 164250 83044 164252
rect 82813 164248 83044 164250
rect 82813 164192 82818 164248
rect 82874 164192 83044 164248
rect 82813 164190 83044 164192
rect 82813 164187 82879 164190
rect 83038 164188 83044 164190
rect 83108 164188 83114 164252
rect 84142 164188 84148 164252
rect 84212 164250 84259 164252
rect 85573 164250 85639 164253
rect 86534 164250 86540 164252
rect 84212 164248 84304 164250
rect 84254 164192 84304 164248
rect 84212 164190 84304 164192
rect 85573 164248 86540 164250
rect 85573 164192 85578 164248
rect 85634 164192 86540 164248
rect 85573 164190 86540 164192
rect 84212 164188 84259 164190
rect 84193 164187 84259 164188
rect 85573 164187 85639 164190
rect 86534 164188 86540 164190
rect 86604 164188 86610 164252
rect 86953 164250 87019 164253
rect 87638 164250 87644 164252
rect 86953 164248 87644 164250
rect 86953 164192 86958 164248
rect 87014 164192 87644 164248
rect 86953 164190 87644 164192
rect 86953 164187 87019 164190
rect 87638 164188 87644 164190
rect 87708 164188 87714 164252
rect 88425 164250 88491 164253
rect 88742 164250 88748 164252
rect 88425 164248 88748 164250
rect 88425 164192 88430 164248
rect 88486 164192 88748 164248
rect 88425 164190 88748 164192
rect 88425 164187 88491 164190
rect 88742 164188 88748 164190
rect 88812 164188 88818 164252
rect 89897 164250 89963 164253
rect 90030 164250 90036 164252
rect 89897 164248 90036 164250
rect 89897 164192 89902 164248
rect 89958 164192 90036 164248
rect 89897 164190 90036 164192
rect 89897 164187 89963 164190
rect 90030 164188 90036 164190
rect 90100 164188 90106 164252
rect 91093 164250 91159 164253
rect 91318 164250 91324 164252
rect 91093 164248 91324 164250
rect 91093 164192 91098 164248
rect 91154 164192 91324 164248
rect 91093 164190 91324 164192
rect 91093 164187 91159 164190
rect 91318 164188 91324 164190
rect 91388 164188 91394 164252
rect 92565 164250 92631 164253
rect 93342 164250 93348 164252
rect 92565 164248 93348 164250
rect 92565 164192 92570 164248
rect 92626 164192 93348 164248
rect 92565 164190 93348 164192
rect 92565 164187 92631 164190
rect 93342 164188 93348 164190
rect 93412 164188 93418 164252
rect 93853 164250 93919 164253
rect 94446 164250 94452 164252
rect 93853 164248 94452 164250
rect 93853 164192 93858 164248
rect 93914 164192 94452 164248
rect 93853 164190 94452 164192
rect 93853 164187 93919 164190
rect 94446 164188 94452 164190
rect 94516 164188 94522 164252
rect 96613 164250 96679 164253
rect 97022 164250 97028 164252
rect 96613 164248 97028 164250
rect 96613 164192 96618 164248
rect 96674 164192 97028 164248
rect 96613 164190 97028 164192
rect 96613 164187 96679 164190
rect 97022 164188 97028 164190
rect 97092 164188 97098 164252
rect 97993 164250 98059 164253
rect 98126 164250 98132 164252
rect 97993 164248 98132 164250
rect 97993 164192 97998 164248
rect 98054 164192 98132 164248
rect 97993 164190 98132 164192
rect 97993 164187 98059 164190
rect 98126 164188 98132 164190
rect 98196 164188 98202 164252
rect 100753 164250 100819 164253
rect 101806 164250 101812 164252
rect 100753 164248 101812 164250
rect 100753 164192 100758 164248
rect 100814 164192 101812 164248
rect 100753 164190 101812 164192
rect 100753 164187 100819 164190
rect 101806 164188 101812 164190
rect 101876 164188 101882 164252
rect 102133 164250 102199 164253
rect 102726 164250 102732 164252
rect 102133 164248 102732 164250
rect 102133 164192 102138 164248
rect 102194 164192 102732 164248
rect 102133 164190 102732 164192
rect 102133 164187 102199 164190
rect 102726 164188 102732 164190
rect 102796 164188 102802 164252
rect 103513 164250 103579 164253
rect 103830 164250 103836 164252
rect 103513 164248 103836 164250
rect 103513 164192 103518 164248
rect 103574 164192 103836 164248
rect 103513 164190 103836 164192
rect 103513 164187 103579 164190
rect 103830 164188 103836 164190
rect 103900 164188 103906 164252
rect 236085 164250 236151 164253
rect 237046 164250 237052 164252
rect 236085 164248 237052 164250
rect 236085 164192 236090 164248
rect 236146 164192 237052 164248
rect 236085 164190 237052 164192
rect 236085 164187 236151 164190
rect 237046 164188 237052 164190
rect 237116 164188 237122 164252
rect 237373 164250 237439 164253
rect 238150 164250 238156 164252
rect 237373 164248 238156 164250
rect 237373 164192 237378 164248
rect 237434 164192 238156 164248
rect 237373 164190 238156 164192
rect 237373 164187 237439 164190
rect 238150 164188 238156 164190
rect 238220 164188 238226 164252
rect 240133 164250 240199 164253
rect 240542 164250 240548 164252
rect 240133 164248 240548 164250
rect 240133 164192 240138 164248
rect 240194 164192 240548 164248
rect 240133 164190 240548 164192
rect 240133 164187 240199 164190
rect 240542 164188 240548 164190
rect 240612 164188 240618 164252
rect 241513 164250 241579 164253
rect 241646 164250 241652 164252
rect 241513 164248 241652 164250
rect 241513 164192 241518 164248
rect 241574 164192 241652 164248
rect 241513 164190 241652 164192
rect 241513 164187 241579 164190
rect 241646 164188 241652 164190
rect 241716 164188 241722 164252
rect 244365 164250 244431 164253
rect 245326 164250 245332 164252
rect 244365 164248 245332 164250
rect 244365 164192 244370 164248
rect 244426 164192 245332 164248
rect 244365 164190 245332 164192
rect 244365 164187 244431 164190
rect 245326 164188 245332 164190
rect 245396 164188 245402 164252
rect 245653 164250 245719 164253
rect 246430 164250 246436 164252
rect 245653 164248 246436 164250
rect 245653 164192 245658 164248
rect 245714 164192 246436 164248
rect 245653 164190 246436 164192
rect 245653 164187 245719 164190
rect 246430 164188 246436 164190
rect 246500 164188 246506 164252
rect 248413 164250 248479 164253
rect 248638 164250 248644 164252
rect 248413 164248 248644 164250
rect 248413 164192 248418 164248
rect 248474 164192 248644 164248
rect 248413 164190 248644 164192
rect 248413 164187 248479 164190
rect 248638 164188 248644 164190
rect 248708 164188 248714 164252
rect 249793 164250 249859 164253
rect 251173 164252 251239 164253
rect 250110 164250 250116 164252
rect 249793 164248 250116 164250
rect 249793 164192 249798 164248
rect 249854 164192 250116 164248
rect 249793 164190 250116 164192
rect 249793 164187 249859 164190
rect 250110 164188 250116 164190
rect 250180 164188 250186 164252
rect 251173 164250 251220 164252
rect 251128 164248 251220 164250
rect 251128 164192 251178 164248
rect 251128 164190 251220 164192
rect 251173 164188 251220 164190
rect 251284 164188 251290 164252
rect 252553 164250 252619 164253
rect 253422 164250 253428 164252
rect 252553 164248 253428 164250
rect 252553 164192 252558 164248
rect 252614 164192 253428 164248
rect 252553 164190 253428 164192
rect 251173 164187 251239 164188
rect 252553 164187 252619 164190
rect 253422 164188 253428 164190
rect 253492 164188 253498 164252
rect 253933 164250 253999 164253
rect 254526 164250 254532 164252
rect 253933 164248 254532 164250
rect 253933 164192 253938 164248
rect 253994 164192 254532 164248
rect 253933 164190 254532 164192
rect 253933 164187 253999 164190
rect 254526 164188 254532 164190
rect 254596 164188 254602 164252
rect 255313 164250 255379 164253
rect 255814 164250 255820 164252
rect 255313 164248 255820 164250
rect 255313 164192 255318 164248
rect 255374 164192 255820 164248
rect 255313 164190 255820 164192
rect 255313 164187 255379 164190
rect 255814 164188 255820 164190
rect 255884 164188 255890 164252
rect 256693 164250 256759 164253
rect 256918 164250 256924 164252
rect 256693 164248 256924 164250
rect 256693 164192 256698 164248
rect 256754 164192 256924 164248
rect 256693 164190 256924 164192
rect 256693 164187 256759 164190
rect 256918 164188 256924 164190
rect 256988 164188 256994 164252
rect 258073 164250 258139 164253
rect 259453 164252 259519 164253
rect 258390 164250 258396 164252
rect 258073 164248 258396 164250
rect 258073 164192 258078 164248
rect 258134 164192 258396 164248
rect 258073 164190 258396 164192
rect 258073 164187 258139 164190
rect 258390 164188 258396 164190
rect 258460 164188 258466 164252
rect 259453 164250 259500 164252
rect 259408 164248 259500 164250
rect 259408 164192 259458 164248
rect 259408 164190 259500 164192
rect 259453 164188 259500 164190
rect 259564 164188 259570 164252
rect 262806 164188 262812 164252
rect 262876 164250 262882 164252
rect 263501 164250 263567 164253
rect 262876 164248 263567 164250
rect 262876 164192 263506 164248
rect 263562 164192 263567 164248
rect 262876 164190 263567 164192
rect 262876 164188 262882 164190
rect 259453 164187 259519 164188
rect 263501 164187 263567 164190
rect 263777 164250 263843 164253
rect 263910 164250 263916 164252
rect 263777 164248 263916 164250
rect 263777 164192 263782 164248
rect 263838 164192 263916 164248
rect 263777 164190 263916 164192
rect 263777 164187 263843 164190
rect 263910 164188 263916 164190
rect 263980 164188 263986 164252
rect 267733 164250 267799 164253
rect 268694 164250 268700 164252
rect 267733 164248 268700 164250
rect 267733 164192 267738 164248
rect 267794 164192 268700 164248
rect 267733 164190 268700 164192
rect 267733 164187 267799 164190
rect 268694 164188 268700 164190
rect 268764 164188 268770 164252
rect 269113 164250 269179 164253
rect 269798 164250 269804 164252
rect 269113 164248 269804 164250
rect 269113 164192 269118 164248
rect 269174 164192 269804 164248
rect 269113 164190 269804 164192
rect 269113 164187 269179 164190
rect 269798 164188 269804 164190
rect 269868 164188 269874 164252
rect 270493 164250 270559 164253
rect 271270 164250 271276 164252
rect 270493 164248 271276 164250
rect 270493 164192 270498 164248
rect 270554 164192 271276 164248
rect 270493 164190 271276 164192
rect 270493 164187 270559 164190
rect 271270 164188 271276 164190
rect 271340 164188 271346 164252
rect 274398 164188 274404 164252
rect 274468 164250 274474 164252
rect 274541 164250 274607 164253
rect 274468 164248 274607 164250
rect 274468 164192 274546 164248
rect 274602 164192 274607 164248
rect 274468 164190 274607 164192
rect 274468 164188 274474 164190
rect 274541 164187 274607 164190
rect 276013 164250 276079 164253
rect 276974 164250 276980 164252
rect 276013 164248 276980 164250
rect 276013 164192 276018 164248
rect 276074 164192 276980 164248
rect 276013 164190 276980 164192
rect 276013 164187 276079 164190
rect 276974 164188 276980 164190
rect 277044 164188 277050 164252
rect 278078 164188 278084 164252
rect 278148 164250 278154 164252
rect 278681 164250 278747 164253
rect 318374 164250 318380 164252
rect 278148 164248 278747 164250
rect 278148 164192 278686 164248
rect 278742 164192 278747 164248
rect 278148 164190 278747 164192
rect 278148 164188 278154 164190
rect 278681 164187 278747 164190
rect 315990 164190 318380 164250
rect 56869 164114 56935 164117
rect 57697 164116 57763 164117
rect 57646 164114 57652 164116
rect 56869 164112 57652 164114
rect 57716 164114 57763 164116
rect 57716 164112 57844 164114
rect 56869 164056 56874 164112
rect 56930 164056 57652 164112
rect 57758 164056 57844 164112
rect 56869 164054 57652 164056
rect 56869 164051 56935 164054
rect 57646 164052 57652 164054
rect 57716 164054 57844 164056
rect 57716 164052 57763 164054
rect 208158 164052 208164 164116
rect 208228 164114 208234 164116
rect 315990 164114 316050 164190
rect 318374 164188 318380 164190
rect 318444 164188 318450 164252
rect 396022 164188 396028 164252
rect 396092 164250 396098 164252
rect 396165 164250 396231 164253
rect 396092 164248 396231 164250
rect 396092 164192 396170 164248
rect 396226 164192 396231 164248
rect 396092 164190 396231 164192
rect 396092 164188 396098 164190
rect 396165 164187 396231 164190
rect 398833 164250 398899 164253
rect 399518 164250 399524 164252
rect 398833 164248 399524 164250
rect 398833 164192 398838 164248
rect 398894 164192 399524 164248
rect 398833 164190 399524 164192
rect 398833 164187 398899 164190
rect 399518 164188 399524 164190
rect 399588 164188 399594 164252
rect 400213 164250 400279 164253
rect 403065 164252 403131 164253
rect 400438 164250 400444 164252
rect 400213 164248 400444 164250
rect 400213 164192 400218 164248
rect 400274 164192 400444 164248
rect 400213 164190 400444 164192
rect 400213 164187 400279 164190
rect 400438 164188 400444 164190
rect 400508 164188 400514 164252
rect 403014 164188 403020 164252
rect 403084 164250 403131 164252
rect 405733 164250 405799 164253
rect 406510 164250 406516 164252
rect 403084 164248 403176 164250
rect 403126 164192 403176 164248
rect 403084 164190 403176 164192
rect 405733 164248 406516 164250
rect 405733 164192 405738 164248
rect 405794 164192 406516 164248
rect 405733 164190 406516 164192
rect 403084 164188 403131 164190
rect 403065 164187 403131 164188
rect 405733 164187 405799 164190
rect 406510 164188 406516 164190
rect 406580 164188 406586 164252
rect 407205 164250 407271 164253
rect 407614 164250 407620 164252
rect 407205 164248 407620 164250
rect 407205 164192 407210 164248
rect 407266 164192 407620 164248
rect 407205 164190 407620 164192
rect 407205 164187 407271 164190
rect 407614 164188 407620 164190
rect 407684 164188 407690 164252
rect 408493 164250 408559 164253
rect 409965 164252 410031 164253
rect 411253 164252 411319 164253
rect 408718 164250 408724 164252
rect 408493 164248 408724 164250
rect 408493 164192 408498 164248
rect 408554 164192 408724 164248
rect 408493 164190 408724 164192
rect 408493 164187 408559 164190
rect 408718 164188 408724 164190
rect 408788 164188 408794 164252
rect 409965 164250 410012 164252
rect 409920 164248 410012 164250
rect 409920 164192 409970 164248
rect 409920 164190 410012 164192
rect 409965 164188 410012 164190
rect 410076 164188 410082 164252
rect 411253 164250 411300 164252
rect 411208 164248 411300 164250
rect 411208 164192 411258 164248
rect 411208 164190 411300 164192
rect 411253 164188 411300 164190
rect 411364 164188 411370 164252
rect 412725 164250 412791 164253
rect 413318 164250 413324 164252
rect 412725 164248 413324 164250
rect 412725 164192 412730 164248
rect 412786 164192 413324 164248
rect 412725 164190 413324 164192
rect 409965 164187 410031 164188
rect 411253 164187 411319 164188
rect 412725 164187 412791 164190
rect 413318 164188 413324 164190
rect 413388 164188 413394 164252
rect 414013 164250 414079 164253
rect 414422 164250 414428 164252
rect 414013 164248 414428 164250
rect 414013 164192 414018 164248
rect 414074 164192 414428 164248
rect 414013 164190 414428 164192
rect 414013 164187 414079 164190
rect 414422 164188 414428 164190
rect 414492 164188 414498 164252
rect 416773 164250 416839 164253
rect 416998 164250 417004 164252
rect 416773 164248 417004 164250
rect 416773 164192 416778 164248
rect 416834 164192 417004 164248
rect 416773 164190 417004 164192
rect 416773 164187 416839 164190
rect 416998 164188 417004 164190
rect 417068 164188 417074 164252
rect 418153 164250 418219 164253
rect 418286 164250 418292 164252
rect 418153 164248 418292 164250
rect 418153 164192 418158 164248
rect 418214 164192 418292 164248
rect 418153 164190 418292 164192
rect 418153 164187 418219 164190
rect 418286 164188 418292 164190
rect 418356 164188 418362 164252
rect 419533 164250 419599 164253
rect 420678 164250 420684 164252
rect 419533 164248 420684 164250
rect 419533 164192 419538 164248
rect 419594 164192 420684 164248
rect 419533 164190 420684 164192
rect 419533 164187 419599 164190
rect 420678 164188 420684 164190
rect 420748 164188 420754 164252
rect 422293 164250 422359 164253
rect 422886 164250 422892 164252
rect 422293 164248 422892 164250
rect 422293 164192 422298 164248
rect 422354 164192 422892 164248
rect 422293 164190 422892 164192
rect 422293 164187 422359 164190
rect 422886 164188 422892 164190
rect 422956 164188 422962 164252
rect 425278 164188 425284 164252
rect 425348 164250 425354 164252
rect 426341 164250 426407 164253
rect 427721 164252 427787 164253
rect 427670 164250 427676 164252
rect 425348 164248 426407 164250
rect 425348 164192 426346 164248
rect 426402 164192 426407 164248
rect 425348 164190 426407 164192
rect 427630 164190 427676 164250
rect 427740 164248 427787 164252
rect 427782 164192 427787 164248
rect 425348 164188 425354 164190
rect 426341 164187 426407 164190
rect 427670 164188 427676 164190
rect 427740 164188 427787 164192
rect 428774 164188 428780 164252
rect 428844 164250 428850 164252
rect 429101 164250 429167 164253
rect 428844 164248 429167 164250
rect 428844 164192 429106 164248
rect 429162 164192 429167 164248
rect 428844 164190 429167 164192
rect 428844 164188 428850 164190
rect 427721 164187 427787 164188
rect 429101 164187 429167 164190
rect 430573 164250 430639 164253
rect 431166 164250 431172 164252
rect 430573 164248 431172 164250
rect 430573 164192 430578 164248
rect 430634 164192 431172 164248
rect 430573 164190 431172 164192
rect 430573 164187 430639 164190
rect 431166 164188 431172 164190
rect 431236 164188 431242 164252
rect 431953 164250 432019 164253
rect 432270 164250 432276 164252
rect 431953 164248 432276 164250
rect 431953 164192 431958 164248
rect 432014 164192 432276 164248
rect 431953 164190 432276 164192
rect 431953 164187 432019 164190
rect 432270 164188 432276 164190
rect 432340 164188 432346 164252
rect 434713 164250 434779 164253
rect 435766 164250 435772 164252
rect 434713 164248 435772 164250
rect 434713 164192 434718 164248
rect 434774 164192 435772 164248
rect 434713 164190 435772 164192
rect 434713 164187 434779 164190
rect 435766 164188 435772 164190
rect 435836 164188 435842 164252
rect 439262 164188 439268 164252
rect 439332 164250 439338 164252
rect 440141 164250 440207 164253
rect 439332 164248 440207 164250
rect 439332 164192 440146 164248
rect 440202 164192 440207 164248
rect 439332 164190 440207 164192
rect 439332 164188 439338 164190
rect 440141 164187 440207 164190
rect 208228 164054 316050 164114
rect 208228 164052 208234 164054
rect 57697 164051 57763 164052
rect 57513 163978 57579 163981
rect 57830 163978 57836 163980
rect 57513 163976 57836 163978
rect 57513 163920 57518 163976
rect 57574 163920 57836 163976
rect 57513 163918 57836 163920
rect 57513 163915 57579 163918
rect 57830 163916 57836 163918
rect 57900 163916 57906 163980
rect 373533 163434 373599 163437
rect 377397 163434 377463 163437
rect 373533 163432 377463 163434
rect 373533 163376 373538 163432
rect 373594 163376 377402 163432
rect 377458 163376 377463 163432
rect 373533 163374 377463 163376
rect 373533 163371 373599 163374
rect 377397 163371 377463 163374
rect -960 162740 480 162980
rect 377254 162964 377260 163028
rect 377324 163026 377330 163028
rect 377397 163026 377463 163029
rect 377324 163024 377463 163026
rect 377324 162968 377402 163024
rect 377458 162968 377463 163024
rect 377324 162966 377463 162968
rect 377324 162964 377330 162966
rect 377397 162963 377463 162966
rect 217542 162692 217548 162756
rect 217612 162754 217618 162756
rect 217869 162754 217935 162757
rect 217612 162752 217935 162754
rect 217612 162696 217874 162752
rect 217930 162696 217935 162752
rect 217612 162694 217935 162696
rect 217612 162692 217618 162694
rect 217869 162691 217935 162694
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 360878 149154 360884 149156
rect 246 149094 360884 149154
rect 360878 149092 360884 149094
rect 360948 149092 360954 149156
rect 217358 146372 217364 146436
rect 217428 146434 217434 146436
rect 276013 146434 276079 146437
rect 217428 146432 276079 146434
rect 217428 146376 276018 146432
rect 276074 146376 276079 146432
rect 217428 146374 276079 146376
rect 217428 146372 217434 146374
rect 276013 146371 276079 146374
rect 56041 146298 56107 146301
rect 58801 146298 58867 146301
rect 59077 146298 59143 146301
rect 103513 146298 103579 146301
rect 56041 146296 59002 146298
rect 56041 146240 56046 146296
rect 56102 146240 58806 146296
rect 58862 146240 59002 146296
rect 56041 146238 59002 146240
rect 56041 146235 56107 146238
rect 58801 146235 58867 146238
rect 58942 146162 59002 146238
rect 59077 146296 103579 146298
rect 59077 146240 59082 146296
rect 59138 146240 103518 146296
rect 103574 146240 103579 146296
rect 59077 146238 103579 146240
rect 59077 146235 59143 146238
rect 103513 146235 103579 146238
rect 219893 146298 219959 146301
rect 267825 146298 267891 146301
rect 219893 146296 267891 146298
rect 219893 146240 219898 146296
rect 219954 146240 267830 146296
rect 267886 146240 267891 146296
rect 219893 146238 267891 146240
rect 219893 146235 219959 146238
rect 267825 146235 267891 146238
rect 377990 146236 377996 146300
rect 378060 146298 378066 146300
rect 379053 146298 379119 146301
rect 426433 146298 426499 146301
rect 378060 146296 379119 146298
rect 378060 146240 379058 146296
rect 379114 146240 379119 146296
rect 378060 146238 379119 146240
rect 378060 146236 378066 146238
rect 379053 146235 379119 146238
rect 383610 146296 426499 146298
rect 383610 146240 426438 146296
rect 426494 146240 426499 146296
rect 383610 146238 426499 146240
rect 102133 146162 102199 146165
rect 58942 146160 102199 146162
rect 58942 146104 102138 146160
rect 102194 146104 102199 146160
rect 58942 146102 102199 146104
rect 102133 146099 102199 146102
rect 216397 146162 216463 146165
rect 263593 146162 263659 146165
rect 216397 146160 263659 146162
rect 216397 146104 216402 146160
rect 216458 146104 263598 146160
rect 263654 146104 263659 146160
rect 216397 146102 263659 146104
rect 216397 146099 216463 146102
rect 263593 146099 263659 146102
rect 377622 146100 377628 146164
rect 377692 146162 377698 146164
rect 378685 146162 378751 146165
rect 383610 146162 383670 146238
rect 426433 146235 426499 146238
rect 377692 146160 383670 146162
rect 377692 146104 378690 146160
rect 378746 146104 383670 146160
rect 377692 146102 383670 146104
rect 377692 146100 377698 146102
rect 378685 146099 378751 146102
rect 73797 146026 73863 146029
rect 100753 146026 100819 146029
rect 73797 146024 100819 146026
rect 73797 145968 73802 146024
rect 73858 145968 100758 146024
rect 100814 145968 100819 146024
rect 73797 145966 100819 145968
rect 73797 145963 73863 145966
rect 100753 145963 100819 145966
rect 213269 145890 213335 145893
rect 237373 145890 237439 145893
rect 213269 145888 237439 145890
rect 213269 145832 213274 145888
rect 213330 145832 237378 145888
rect 237434 145832 237439 145888
rect 213269 145830 237439 145832
rect 213269 145827 213335 145830
rect 237373 145827 237439 145830
rect 379053 145890 379119 145893
rect 415393 145890 415459 145893
rect 379053 145888 415459 145890
rect 379053 145832 379058 145888
rect 379114 145832 415398 145888
rect 415454 145832 415459 145888
rect 379053 145830 415459 145832
rect 379053 145827 379119 145830
rect 415393 145827 415459 145830
rect 58709 145754 58775 145757
rect 92565 145754 92631 145757
rect 58709 145752 92631 145754
rect 58709 145696 58714 145752
rect 58770 145696 92570 145752
rect 92626 145696 92631 145752
rect 58709 145694 92631 145696
rect 58709 145691 58775 145694
rect 92565 145691 92631 145694
rect 210877 145754 210943 145757
rect 220077 145754 220143 145757
rect 267733 145754 267799 145757
rect 210877 145752 267799 145754
rect 210877 145696 210882 145752
rect 210938 145696 220082 145752
rect 220138 145696 267738 145752
rect 267794 145696 267799 145752
rect 210877 145694 267799 145696
rect 210877 145691 210943 145694
rect 220077 145691 220143 145694
rect 267733 145691 267799 145694
rect 370313 145754 370379 145757
rect 377213 145754 377279 145757
rect 423673 145754 423739 145757
rect 370313 145752 423739 145754
rect 370313 145696 370318 145752
rect 370374 145696 377218 145752
rect 377274 145696 423678 145752
rect 423734 145696 423739 145752
rect 370313 145694 423739 145696
rect 370313 145691 370379 145694
rect 377213 145691 377279 145694
rect 423673 145691 423739 145694
rect 58893 145618 58959 145621
rect 107653 145618 107719 145621
rect 58893 145616 107719 145618
rect 58893 145560 58898 145616
rect 58954 145560 107658 145616
rect 107714 145560 107719 145616
rect 58893 145558 107719 145560
rect 58893 145555 58959 145558
rect 107653 145555 107719 145558
rect 214925 145618 214991 145621
rect 269113 145618 269179 145621
rect 214925 145616 269179 145618
rect 214925 145560 214930 145616
rect 214986 145560 269118 145616
rect 269174 145560 269179 145616
rect 214925 145558 269179 145560
rect 214925 145555 214991 145558
rect 269113 145555 269179 145558
rect 369025 145618 369091 145621
rect 379697 145618 379763 145621
rect 427813 145618 427879 145621
rect 369025 145616 427879 145618
rect 369025 145560 369030 145616
rect 369086 145560 379702 145616
rect 379758 145560 427818 145616
rect 427874 145560 427879 145616
rect 369025 145558 427879 145560
rect 369025 145555 369091 145558
rect 379697 145555 379763 145558
rect 427813 145555 427879 145558
rect 510613 145482 510679 145485
rect 510838 145482 510844 145484
rect 510613 145480 510844 145482
rect 510613 145424 510618 145480
rect 510674 145424 510844 145480
rect 510613 145422 510844 145424
rect 510613 145419 510679 145422
rect 510838 145420 510844 145422
rect 510908 145420 510914 145484
rect 215845 145074 215911 145077
rect 216397 145074 216463 145077
rect 215845 145072 216463 145074
rect 215845 145016 215850 145072
rect 215906 145016 216402 145072
rect 216458 145016 216463 145072
rect 215845 145014 216463 145016
rect 215845 145011 215911 145014
rect 216397 145011 216463 145014
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 190862 144876 190868 144940
rect 190932 144938 190938 144940
rect 191281 144938 191347 144941
rect 190932 144936 191347 144938
rect 190932 144880 191286 144936
rect 191342 144880 191347 144936
rect 190932 144878 191347 144880
rect 190932 144876 190938 144878
rect 179689 144875 179755 144876
rect 191281 144875 191347 144878
rect 219157 144938 219223 144941
rect 219893 144938 219959 144941
rect 338481 144940 338547 144941
rect 338430 144938 338436 144940
rect 219157 144936 219959 144938
rect 219157 144880 219162 144936
rect 219218 144880 219898 144936
rect 219954 144880 219959 144936
rect 219157 144878 219959 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 219157 144875 219223 144878
rect 219893 144875 219959 144878
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144940
rect 499868 144938 499874 144940
rect 500217 144938 500283 144941
rect 499868 144936 500283 144938
rect 499868 144880 500222 144936
rect 500278 144880 500283 144936
rect 499868 144878 500283 144880
rect 499868 144876 499874 144878
rect 500217 144875 500283 144878
rect 377806 144060 377812 144124
rect 377876 144122 377882 144124
rect 440233 144122 440299 144125
rect 377876 144120 440299 144122
rect 377876 144064 440238 144120
rect 440294 144064 440299 144120
rect 377876 144062 440299 144064
rect 377876 144060 377882 144062
rect 440233 144059 440299 144062
rect 57278 140796 57284 140860
rect 57348 140858 57354 140860
rect 59353 140858 59419 140861
rect 57348 140856 59419 140858
rect 57348 140800 59358 140856
rect 59414 140800 59419 140856
rect 57348 140798 59419 140800
rect 57348 140796 57354 140798
rect 59353 140795 59419 140798
rect 358905 139362 358971 139365
rect 519261 139362 519327 139365
rect 356562 139360 358971 139362
rect 356562 139304 358910 139360
rect 358966 139304 358971 139360
rect 356562 139302 358971 139304
rect 198825 139226 198891 139229
rect 197126 139224 198891 139226
rect 197126 139220 198830 139224
rect 196604 139168 198830 139220
rect 198886 139168 198891 139224
rect 356562 139190 356622 139302
rect 358905 139299 358971 139302
rect 516558 139360 519327 139362
rect 516558 139304 519266 139360
rect 519322 139304 519327 139360
rect 516558 139302 519327 139304
rect 516558 139190 516618 139302
rect 519261 139299 519327 139302
rect 583520 139212 584960 139452
rect 196604 139166 198891 139168
rect 196604 139160 197186 139166
rect 198825 139163 198891 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 57145 97474 57211 97477
rect 57145 97472 60062 97474
rect 57145 97416 57150 97472
rect 57206 97416 60062 97472
rect 57145 97414 60062 97416
rect 57145 97411 57211 97414
rect 60002 96894 60062 97414
rect 216857 96930 216923 96933
rect 377029 96930 377095 96933
rect 216857 96928 219450 96930
rect 216857 96872 216862 96928
rect 216918 96924 219450 96928
rect 377029 96928 379530 96930
rect 216918 96872 220064 96924
rect 216857 96870 220064 96872
rect 216857 96867 216923 96870
rect 219390 96864 220064 96870
rect 377029 96872 377034 96928
rect 377090 96924 379530 96928
rect 377090 96872 380052 96924
rect 377029 96870 380052 96872
rect 377029 96867 377095 96870
rect 379470 96864 380052 96870
rect 56593 96522 56659 96525
rect 56593 96520 60062 96522
rect 56593 96464 56598 96520
rect 56654 96464 60062 96520
rect 56593 96462 60062 96464
rect 56593 96459 56659 96462
rect 60002 95942 60062 96462
rect 216949 95978 217015 95981
rect 376753 95978 376819 95981
rect 216949 95976 219450 95978
rect 216949 95920 216954 95976
rect 217010 95972 219450 95976
rect 376753 95976 379530 95978
rect 217010 95920 220064 95972
rect 216949 95918 220064 95920
rect 216949 95915 217015 95918
rect 219390 95912 220064 95918
rect 376753 95920 376758 95976
rect 376814 95972 379530 95976
rect 376814 95920 380052 95972
rect 376753 95918 380052 95920
rect 376753 95915 376819 95918
rect 379470 95912 380052 95918
rect 56777 93802 56843 93805
rect 217685 93802 217751 93805
rect 376845 93802 376911 93805
rect 56777 93800 60062 93802
rect 56777 93744 56782 93800
rect 56838 93744 60062 93800
rect 56777 93742 60062 93744
rect 217685 93800 219450 93802
rect 217685 93744 217690 93800
rect 217746 93796 219450 93800
rect 376845 93800 379530 93802
rect 217746 93744 220064 93796
rect 217685 93742 220064 93744
rect 56777 93739 56843 93742
rect 217685 93739 217751 93742
rect 219390 93736 220064 93742
rect 376845 93744 376850 93800
rect 376906 93796 379530 93800
rect 376906 93744 380052 93796
rect 376845 93742 380052 93744
rect 376845 93739 376911 93742
rect 379470 93736 380052 93742
rect 57329 93394 57395 93397
rect 57329 93392 60062 93394
rect 57329 93336 57334 93392
rect 57390 93336 60062 93392
rect 57329 93334 60062 93336
rect 57329 93331 57395 93334
rect 60002 92814 60062 93334
rect 217409 92850 217475 92853
rect 376937 92850 377003 92853
rect 217409 92848 219450 92850
rect 217409 92792 217414 92848
rect 217470 92844 219450 92848
rect 376937 92848 379530 92850
rect 217470 92792 220064 92844
rect 217409 92790 220064 92792
rect 217409 92787 217475 92790
rect 219390 92784 220064 92790
rect 376937 92792 376942 92848
rect 376998 92844 379530 92848
rect 376998 92792 380052 92844
rect 376937 92790 380052 92792
rect 376937 92787 377003 92790
rect 379470 92784 380052 92790
rect 57605 91082 57671 91085
rect 217501 91082 217567 91085
rect 377765 91082 377831 91085
rect 57605 91080 60062 91082
rect 57605 91024 57610 91080
rect 57666 91024 60062 91080
rect 57605 91022 60062 91024
rect 217501 91080 219450 91082
rect 217501 91024 217506 91080
rect 217562 91076 219450 91080
rect 377765 91080 379530 91082
rect 217562 91024 220064 91076
rect 217501 91022 220064 91024
rect 57605 91019 57671 91022
rect 217501 91019 217567 91022
rect 219390 91016 220064 91022
rect 377765 91024 377770 91080
rect 377826 91076 379530 91080
rect 377826 91024 380052 91076
rect 377765 91022 380052 91024
rect 377765 91019 377831 91022
rect 379470 91016 380052 91022
rect 57421 90538 57487 90541
rect 57421 90536 60062 90538
rect 57421 90480 57426 90536
rect 57482 90480 60062 90536
rect 57421 90478 60062 90480
rect 57421 90475 57487 90478
rect 60002 89958 60062 90478
rect 217225 89994 217291 89997
rect 377305 89994 377371 89997
rect 217225 89992 219450 89994
rect 217225 89936 217230 89992
rect 217286 89988 219450 89992
rect 377305 89992 379530 89994
rect 217286 89936 220064 89988
rect 217225 89934 220064 89936
rect 217225 89931 217291 89934
rect 219390 89928 220064 89934
rect 377305 89936 377310 89992
rect 377366 89988 379530 89992
rect 377366 89936 380052 89988
rect 377305 89934 380052 89936
rect 377305 89931 377371 89934
rect 379470 89928 380052 89934
rect 57789 88226 57855 88229
rect 217593 88226 217659 88229
rect 377949 88226 378015 88229
rect 57789 88224 60062 88226
rect 57789 88168 57794 88224
rect 57850 88168 60062 88224
rect 57789 88166 60062 88168
rect 217593 88224 219450 88226
rect 217593 88168 217598 88224
rect 217654 88220 219450 88224
rect 377949 88224 379530 88226
rect 217654 88168 220064 88220
rect 217593 88166 220064 88168
rect 57789 88163 57855 88166
rect 217593 88163 217659 88166
rect 219390 88160 220064 88166
rect 377949 88168 377954 88224
rect 378010 88220 379530 88224
rect 378010 88168 380052 88220
rect 377949 88166 380052 88168
rect 377949 88163 378015 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 359365 79930 359431 79933
rect 518893 79930 518959 79933
rect 520181 79930 520247 79933
rect 356562 79928 359431 79930
rect 356562 79872 359370 79928
rect 359426 79872 359431 79928
rect 356562 79870 359431 79872
rect 199377 79386 199443 79389
rect 197126 79384 199443 79386
rect 197126 79380 199382 79384
rect 196604 79328 199382 79380
rect 199438 79328 199443 79384
rect 356562 79350 356622 79870
rect 359365 79867 359431 79870
rect 516558 79928 520247 79930
rect 516558 79872 518898 79928
rect 518954 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 518893 79867 518959 79870
rect 520181 79867 520247 79870
rect 196604 79326 199443 79328
rect 196604 79320 197186 79326
rect 199377 79323 199443 79326
rect 359089 78298 359155 78301
rect 519445 78298 519511 78301
rect 356562 78296 359155 78298
rect 356562 78240 359094 78296
rect 359150 78240 359155 78296
rect 356562 78238 359155 78240
rect 199285 77754 199351 77757
rect 197126 77752 199351 77754
rect 197126 77748 199290 77752
rect 196604 77696 199290 77748
rect 199346 77696 199351 77752
rect 356562 77718 356622 78238
rect 359089 78235 359155 78238
rect 516558 78296 519511 78298
rect 516558 78240 519450 78296
rect 519506 78240 519511 78296
rect 516558 78238 519511 78240
rect 516558 77718 516618 78238
rect 519445 78235 519511 78238
rect 196604 77694 199351 77696
rect 196604 77688 197186 77694
rect 199285 77691 199351 77694
rect 359273 76938 359339 76941
rect 356562 76936 359339 76938
rect 356562 76880 359278 76936
rect 359334 76880 359339 76936
rect 356562 76878 359339 76880
rect 199101 76394 199167 76397
rect 197126 76392 199167 76394
rect 197126 76388 199106 76392
rect 196604 76336 199106 76388
rect 199162 76336 199167 76392
rect 356562 76358 356622 76878
rect 359273 76875 359339 76878
rect 519077 76802 519143 76805
rect 516558 76800 519143 76802
rect 516558 76744 519082 76800
rect 519138 76744 519143 76800
rect 516558 76742 519143 76744
rect 516558 76358 516618 76742
rect 519077 76739 519143 76742
rect 196604 76334 199167 76336
rect 196604 76328 197186 76334
rect 199101 76331 199167 76334
rect 359181 75442 359247 75445
rect 519353 75442 519419 75445
rect 356562 75440 359247 75442
rect 356562 75384 359186 75440
rect 359242 75384 359247 75440
rect 356562 75382 359247 75384
rect 198733 74898 198799 74901
rect 197126 74896 198799 74898
rect 197126 74892 198738 74896
rect 196604 74840 198738 74892
rect 198794 74840 198799 74896
rect 356562 74862 356622 75382
rect 359181 75379 359247 75382
rect 516558 75440 519419 75442
rect 516558 75384 519358 75440
rect 519414 75384 519419 75440
rect 516558 75382 519419 75384
rect 516558 74862 516618 75382
rect 519353 75379 519419 75382
rect 196604 74838 198799 74840
rect 196604 74832 197186 74838
rect 198733 74835 198799 74838
rect 518985 74218 519051 74221
rect 516558 74216 519051 74218
rect 516558 74160 518990 74216
rect 519046 74160 519051 74216
rect 516558 74158 519051 74160
rect 358997 74082 359063 74085
rect 356562 74080 359063 74082
rect 356562 74024 359002 74080
rect 359058 74024 359063 74080
rect 356562 74022 359063 74024
rect 199193 73674 199259 73677
rect 197126 73672 199259 73674
rect 197126 73668 199198 73672
rect 196604 73616 199198 73668
rect 199254 73616 199259 73672
rect 356562 73638 356622 74022
rect 358997 74019 359063 74022
rect 516558 73638 516618 74158
rect 518985 74155 519051 74158
rect 196604 73614 199259 73616
rect 196604 73608 197186 73614
rect 199193 73611 199259 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 57462 70348 57468 70412
rect 57532 70410 57538 70412
rect 57532 70350 60062 70410
rect 57532 70348 57538 70350
rect 60002 69966 60062 70350
rect 216673 70002 216739 70005
rect 376937 70002 377003 70005
rect 216673 70000 219450 70002
rect 216673 69944 216678 70000
rect 216734 69996 219450 70000
rect 376937 70000 379530 70002
rect 216734 69944 220064 69996
rect 216673 69942 220064 69944
rect 216673 69939 216739 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 216673 68370 216739 68373
rect 217961 68370 218027 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68312 217966 68368
rect 218022 68364 219450 68368
rect 376937 68368 379530 68370
rect 218022 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 217961 68307 218027 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 44950 67764 44956 67828
rect 45020 67826 45026 67828
rect 60002 67826 60062 68062
rect 216070 68036 216076 68100
rect 216140 68098 216146 68100
rect 216140 68092 219450 68098
rect 216140 68038 220064 68092
rect 216140 68036 216146 68038
rect 219390 68032 220064 68038
rect 374678 68036 374684 68100
rect 374748 68098 374754 68100
rect 374748 68092 379530 68098
rect 374748 68038 380052 68092
rect 374748 68036 374754 68038
rect 379470 68032 380052 68038
rect 45020 67766 60062 67826
rect 45020 67764 45026 67766
rect 218697 60620 218763 60621
rect 219249 60620 219315 60621
rect 218646 60618 218652 60620
rect 218606 60558 218652 60618
rect 218716 60616 218763 60620
rect 219198 60618 219204 60620
rect 218758 60560 218763 60616
rect 218646 60556 218652 60558
rect 218716 60556 218763 60560
rect 219158 60558 219204 60618
rect 219268 60616 219315 60620
rect 219310 60560 219315 60616
rect 219198 60556 219204 60558
rect 219268 60556 219315 60560
rect 218697 60555 218763 60556
rect 219249 60555 219315 60556
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 94497 59804 94563 59805
rect 99465 59804 99531 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 94497 59800 94550 59804
rect 94614 59802 94620 59804
rect 99440 59802 99446 59804
rect 94497 59744 94502 59800
rect 83190 59740 83196 59742
rect 94497 59740 94550 59744
rect 94614 59742 94654 59802
rect 99374 59742 99446 59802
rect 99510 59800 99531 59804
rect 99526 59744 99531 59800
rect 94614 59740 94620 59742
rect 99440 59740 99446 59742
rect 99510 59740 99531 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 94497 59739 94563 59740
rect 99465 59739 99531 59740
rect 102777 59804 102843 59805
rect 105905 59804 105971 59805
rect 237097 59804 237163 59805
rect 255865 59804 255931 59805
rect 256969 59804 257035 59805
rect 262857 59804 262923 59805
rect 102777 59800 102846 59804
rect 102777 59744 102782 59800
rect 102838 59744 102846 59800
rect 102777 59740 102846 59744
rect 102910 59802 102916 59804
rect 102910 59742 102934 59802
rect 105905 59800 105974 59804
rect 105905 59744 105910 59800
rect 105966 59744 105974 59800
rect 102910 59740 102916 59742
rect 105905 59740 105974 59744
rect 106038 59802 106044 59804
rect 106038 59742 106062 59802
rect 237097 59800 237142 59804
rect 237206 59802 237212 59804
rect 237097 59744 237102 59800
rect 106038 59740 106044 59742
rect 237097 59740 237142 59744
rect 237206 59742 237254 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 255865 59744 255870 59800
rect 237206 59740 237212 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 256969 59800 256998 59804
rect 257062 59802 257068 59804
rect 262840 59802 262846 59804
rect 256969 59744 256974 59800
rect 255974 59740 255980 59742
rect 256969 59740 256998 59744
rect 257062 59742 257126 59802
rect 262766 59742 262846 59802
rect 262910 59800 262923 59804
rect 262918 59744 262923 59800
rect 257062 59740 257068 59742
rect 262840 59740 262846 59742
rect 262910 59740 262923 59744
rect 102777 59739 102843 59740
rect 105905 59739 105971 59740
rect 237097 59739 237163 59740
rect 255865 59739 255931 59740
rect 256969 59739 257035 59740
rect 262857 59739 262923 59740
rect 263869 59804 263935 59805
rect 396073 59804 396139 59805
rect 263869 59800 263934 59804
rect 263869 59744 263874 59800
rect 263930 59744 263934 59800
rect 263869 59740 263934 59744
rect 263998 59802 264004 59804
rect 396048 59802 396054 59804
rect 263998 59742 264026 59802
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 263998 59740 264004 59742
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 263869 59739 263935 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 416037 59804 416103 59805
rect 416957 59804 417023 59805
rect 422845 59804 422911 59805
rect 423949 59804 424015 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 416037 59800 416046 59804
rect 416110 59802 416116 59804
rect 416037 59744 416042 59800
rect 397206 59740 397212 59742
rect 416037 59740 416046 59744
rect 416110 59742 416194 59802
rect 416957 59800 416998 59804
rect 417062 59802 417068 59804
rect 422840 59802 422846 59804
rect 416957 59744 416962 59800
rect 416110 59740 416116 59742
rect 416957 59740 416998 59744
rect 417062 59742 417114 59802
rect 422754 59742 422846 59802
rect 417062 59740 417068 59742
rect 422840 59740 422846 59742
rect 422910 59740 422916 59804
rect 423928 59802 423934 59804
rect 423858 59742 423934 59802
rect 423998 59800 424015 59804
rect 424010 59744 424015 59800
rect 423928 59740 423934 59742
rect 423998 59740 424015 59744
rect 397085 59739 397151 59740
rect 416037 59739 416103 59740
rect 416957 59739 417023 59740
rect 422845 59739 422911 59740
rect 423949 59739 424015 59740
rect 107561 59668 107627 59669
rect 258073 59668 258139 59669
rect 260649 59668 260715 59669
rect 261753 59668 261819 59669
rect 308489 59668 308555 59669
rect 315849 59668 315915 59669
rect 403065 59668 403131 59669
rect 404169 59668 404235 59669
rect 105288 59666 105294 59668
rect 84150 59606 105294 59666
rect 57646 59468 57652 59532
rect 57716 59530 57722 59532
rect 84150 59530 84210 59606
rect 105288 59604 105294 59606
rect 105358 59604 105364 59668
rect 107561 59664 107606 59668
rect 107670 59666 107676 59668
rect 107561 59608 107566 59664
rect 107561 59604 107606 59608
rect 107670 59606 107718 59666
rect 258073 59664 258086 59668
rect 258150 59666 258156 59668
rect 258073 59608 258078 59664
rect 107670 59604 107676 59606
rect 258073 59604 258086 59608
rect 258150 59606 258230 59666
rect 260649 59664 260670 59668
rect 260734 59666 260740 59668
rect 260649 59608 260654 59664
rect 258150 59604 258156 59606
rect 260649 59604 260670 59608
rect 260734 59606 260806 59666
rect 260734 59604 260740 59606
rect 261752 59604 261758 59668
rect 261822 59666 261828 59668
rect 261822 59606 261910 59666
rect 308489 59664 308542 59668
rect 308606 59666 308612 59668
rect 308489 59608 308494 59664
rect 261822 59604 261828 59606
rect 308489 59604 308542 59608
rect 308606 59606 308646 59666
rect 315849 59664 315886 59668
rect 315950 59666 315956 59668
rect 315849 59608 315854 59664
rect 308606 59604 308612 59606
rect 315849 59604 315886 59608
rect 315950 59606 316006 59666
rect 403065 59664 403126 59668
rect 403065 59608 403070 59664
rect 315950 59604 315956 59606
rect 403065 59604 403126 59608
rect 403190 59666 403196 59668
rect 403190 59606 403222 59666
rect 404169 59664 404214 59668
rect 404278 59666 404284 59668
rect 412541 59666 412607 59669
rect 423489 59668 423555 59669
rect 413456 59666 413462 59668
rect 404169 59608 404174 59664
rect 403190 59604 403196 59606
rect 404169 59604 404214 59608
rect 404278 59606 404326 59666
rect 412541 59664 413462 59666
rect 412541 59608 412546 59664
rect 412602 59608 413462 59664
rect 412541 59606 413462 59608
rect 404278 59604 404284 59606
rect 107561 59603 107627 59604
rect 258073 59603 258139 59604
rect 260649 59603 260715 59604
rect 261753 59603 261819 59604
rect 308489 59603 308555 59604
rect 315849 59603 315915 59604
rect 403065 59603 403131 59604
rect 404169 59603 404235 59604
rect 412541 59603 412607 59606
rect 413456 59604 413462 59606
rect 413526 59604 413532 59668
rect 423489 59664 423526 59668
rect 423590 59666 423596 59668
rect 423489 59608 423494 59664
rect 423489 59604 423526 59608
rect 423590 59606 423646 59666
rect 423590 59604 423596 59606
rect 423489 59603 423555 59604
rect 57716 59470 84210 59530
rect 89989 59532 90055 59533
rect 95877 59532 95943 59533
rect 96981 59532 97047 59533
rect 100753 59532 100819 59533
rect 89989 59528 90036 59532
rect 90100 59530 90106 59532
rect 89989 59472 89994 59528
rect 57716 59468 57722 59470
rect 89989 59468 90036 59472
rect 90100 59470 90146 59530
rect 95877 59528 95924 59532
rect 95988 59530 95994 59532
rect 95877 59472 95882 59528
rect 90100 59468 90106 59470
rect 95877 59468 95924 59472
rect 95988 59470 96034 59530
rect 96981 59528 97028 59532
rect 97092 59530 97098 59532
rect 100702 59530 100708 59532
rect 96981 59472 96986 59528
rect 95988 59468 95994 59470
rect 96981 59468 97028 59472
rect 97092 59470 97138 59530
rect 100662 59470 100708 59530
rect 100772 59528 100819 59532
rect 100814 59472 100819 59528
rect 97092 59468 97098 59470
rect 100702 59468 100708 59470
rect 100772 59468 100819 59472
rect 89989 59467 90055 59468
rect 95877 59467 95943 59468
rect 96981 59467 97047 59468
rect 100753 59467 100819 59468
rect 101765 59532 101831 59533
rect 101765 59528 101812 59532
rect 101876 59530 101882 59532
rect 101765 59472 101770 59528
rect 101765 59468 101812 59472
rect 101876 59470 101922 59530
rect 583520 59516 584960 59756
rect 101876 59468 101882 59470
rect 101765 59467 101831 59468
rect 418153 59396 418219 59397
rect 48446 59332 48452 59396
rect 48516 59394 48522 59396
rect 113582 59394 113588 59396
rect 48516 59334 113588 59394
rect 48516 59332 48522 59334
rect 113582 59332 113588 59334
rect 113652 59332 113658 59396
rect 200614 59332 200620 59396
rect 200684 59394 200690 59396
rect 263542 59394 263548 59396
rect 200684 59334 263548 59394
rect 200684 59332 200690 59334
rect 263542 59332 263548 59334
rect 263612 59332 263618 59396
rect 418102 59394 418108 59396
rect 279006 59334 279434 59394
rect 418062 59334 418108 59394
rect 418172 59392 418219 59396
rect 418214 59336 418219 59392
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 52310 59196 52316 59260
rect 52380 59258 52386 59260
rect 143574 59258 143580 59260
rect 52380 59198 143580 59258
rect 52380 59196 52386 59198
rect 143574 59196 143580 59198
rect 143644 59196 143650 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 206686 59196 206692 59260
rect 206756 59258 206762 59260
rect 279006 59258 279066 59334
rect 279233 59260 279299 59261
rect 279182 59258 279188 59260
rect 206756 59198 279066 59258
rect 279142 59198 279188 59258
rect 279252 59256 279299 59260
rect 279294 59200 279299 59256
rect 206756 59196 206762 59198
rect 279182 59196 279188 59198
rect 279252 59196 279299 59200
rect 279374 59258 279434 59334
rect 418102 59332 418108 59334
rect 418172 59332 418219 59336
rect 418153 59331 418219 59332
rect 419349 59396 419415 59397
rect 420637 59396 420703 59397
rect 421741 59396 421807 59397
rect 425973 59396 426039 59397
rect 428181 59396 428247 59397
rect 453389 59396 453455 59397
rect 419349 59392 419396 59396
rect 419460 59394 419466 59396
rect 419349 59336 419354 59392
rect 419349 59332 419396 59336
rect 419460 59334 419506 59394
rect 420637 59392 420684 59396
rect 420748 59394 420754 59396
rect 420637 59336 420642 59392
rect 419460 59332 419466 59334
rect 420637 59332 420684 59336
rect 420748 59334 420794 59394
rect 421741 59392 421788 59396
rect 421852 59394 421858 59396
rect 421741 59336 421746 59392
rect 420748 59332 420754 59334
rect 421741 59332 421788 59336
rect 421852 59334 421898 59394
rect 425973 59392 426020 59396
rect 426084 59394 426090 59396
rect 425973 59336 425978 59392
rect 421852 59332 421858 59334
rect 425973 59332 426020 59336
rect 426084 59334 426130 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 426084 59332 426090 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 453389 59392 453436 59396
rect 453500 59394 453506 59396
rect 453389 59336 453394 59392
rect 428292 59332 428298 59334
rect 453389 59332 453436 59336
rect 453500 59334 453546 59394
rect 453500 59332 453506 59334
rect 419349 59331 419415 59332
rect 420637 59331 420703 59332
rect 421741 59331 421807 59332
rect 425973 59331 426039 59332
rect 428181 59331 428247 59332
rect 453389 59331 453455 59332
rect 290917 59260 290983 59261
rect 300853 59260 300919 59261
rect 320909 59260 320975 59261
rect 325877 59260 325943 59261
rect 285990 59258 285996 59260
rect 279374 59198 285996 59258
rect 285990 59196 285996 59198
rect 286060 59196 286066 59260
rect 290917 59256 290964 59260
rect 291028 59258 291034 59260
rect 290917 59200 290922 59256
rect 290917 59196 290964 59200
rect 291028 59198 291074 59258
rect 300853 59256 300900 59260
rect 300964 59258 300970 59260
rect 300853 59200 300858 59256
rect 291028 59196 291034 59198
rect 300853 59196 300900 59200
rect 300964 59198 301010 59258
rect 320909 59256 320956 59260
rect 321020 59258 321026 59260
rect 320909 59200 320914 59256
rect 300964 59196 300970 59198
rect 320909 59196 320956 59200
rect 321020 59198 321066 59258
rect 325877 59256 325924 59260
rect 325988 59258 325994 59260
rect 325877 59200 325882 59256
rect 321020 59196 321026 59198
rect 325877 59196 325924 59200
rect 325988 59198 326034 59258
rect 325988 59196 325994 59198
rect 360694 59196 360700 59260
rect 360764 59258 360770 59260
rect 483422 59258 483428 59260
rect 360764 59198 483428 59258
rect 360764 59196 360770 59198
rect 483422 59196 483428 59198
rect 483492 59196 483498 59260
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 279233 59195 279299 59196
rect 290917 59195 290983 59196
rect 300853 59195 300919 59196
rect 320909 59195 320975 59196
rect 325877 59195 325943 59196
rect 54886 59060 54892 59124
rect 54956 59122 54962 59124
rect 140814 59122 140820 59124
rect 54956 59062 140820 59122
rect 54956 59060 54962 59062
rect 140814 59060 140820 59062
rect 140884 59060 140890 59124
rect 209630 59060 209636 59124
rect 209700 59122 209706 59124
rect 280838 59122 280844 59124
rect 209700 59062 280844 59122
rect 209700 59060 209706 59062
rect 280838 59060 280844 59062
rect 280908 59060 280914 59124
rect 371918 59060 371924 59124
rect 371988 59122 371994 59124
rect 480846 59122 480852 59124
rect 371988 59062 480852 59122
rect 371988 59060 371994 59062
rect 480846 59060 480852 59062
rect 480916 59060 480922 59124
rect 138381 58988 138447 58989
rect 475837 58988 475903 58989
rect 52126 58924 52132 58988
rect 52196 58986 52202 58988
rect 135846 58986 135852 58988
rect 52196 58926 135852 58986
rect 52196 58924 52202 58926
rect 135846 58924 135852 58926
rect 135916 58924 135922 58988
rect 138381 58984 138428 58988
rect 138492 58986 138498 58988
rect 138381 58928 138386 58984
rect 138381 58924 138428 58928
rect 138492 58926 138538 58986
rect 138492 58924 138498 58926
rect 198038 58924 198044 58988
rect 198108 58986 198114 58988
rect 268326 58986 268332 58988
rect 198108 58926 268332 58986
rect 198108 58924 198114 58926
rect 268326 58924 268332 58926
rect 268396 58924 268402 58988
rect 366214 58924 366220 58988
rect 366284 58986 366290 58988
rect 468518 58986 468524 58988
rect 366284 58926 468524 58986
rect 366284 58924 366290 58926
rect 468518 58924 468524 58926
rect 468588 58924 468594 58988
rect 475837 58984 475884 58988
rect 475948 58986 475954 58988
rect 475837 58928 475842 58984
rect 475837 58924 475884 58928
rect 475948 58926 475994 58986
rect 475948 58924 475954 58926
rect 138381 58923 138447 58924
rect 475837 58923 475903 58924
rect 48630 58788 48636 58852
rect 48700 58850 48706 58852
rect 111006 58850 111012 58852
rect 48700 58790 111012 58850
rect 48700 58788 48706 58790
rect 111006 58788 111012 58790
rect 111076 58788 111082 58852
rect 206870 58788 206876 58852
rect 206940 58850 206946 58852
rect 276054 58850 276060 58852
rect 206940 58790 276060 58850
rect 206940 58788 206946 58790
rect 276054 58788 276060 58790
rect 276124 58788 276130 58852
rect 373758 58788 373764 58852
rect 373828 58850 373834 58852
rect 473486 58850 473492 58852
rect 373828 58790 473492 58850
rect 373828 58788 373834 58790
rect 473486 58788 473492 58790
rect 473556 58788 473562 58852
rect -960 58578 480 58668
rect 59302 58652 59308 58716
rect 59372 58714 59378 58716
rect 120942 58714 120948 58716
rect 59372 58654 120948 58714
rect 59372 58652 59378 58654
rect 120942 58652 120948 58654
rect 121012 58652 121018 58716
rect 197854 58652 197860 58716
rect 197924 58714 197930 58716
rect 253606 58714 253612 58716
rect 197924 58654 253612 58714
rect 197924 58652 197930 58654
rect 253606 58652 253612 58654
rect 253676 58652 253682 58716
rect 371734 58652 371740 58716
rect 371804 58714 371810 58716
rect 463550 58714 463556 58716
rect 371804 58654 463556 58714
rect 371804 58652 371810 58654
rect 463550 58652 463556 58654
rect 463620 58652 463626 58716
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 47894 58516 47900 58580
rect 47964 58578 47970 58580
rect 108246 58578 108252 58580
rect 47964 58518 108252 58578
rect 47964 58516 47970 58518
rect 108246 58516 108252 58518
rect 108316 58516 108322 58580
rect 202270 58516 202276 58580
rect 202340 58578 202346 58580
rect 250662 58578 250668 58580
rect 202340 58518 250668 58578
rect 202340 58516 202346 58518
rect 250662 58516 250668 58518
rect 250732 58516 250738 58580
rect 370446 58516 370452 58580
rect 370516 58578 370522 58580
rect 458398 58578 458404 58580
rect 370516 58518 458404 58578
rect 370516 58516 370522 58518
rect 458398 58516 458404 58518
rect 458468 58516 458474 58580
rect 59118 58380 59124 58444
rect 59188 58442 59194 58444
rect 101070 58442 101076 58444
rect 59188 58382 101076 58442
rect 59188 58380 59194 58382
rect 101070 58380 101076 58382
rect 101140 58380 101146 58444
rect 217542 58380 217548 58444
rect 217612 58442 217618 58444
rect 259494 58442 259500 58444
rect 217612 58382 259500 58442
rect 217612 58380 217618 58382
rect 259494 58380 259500 58382
rect 259564 58380 259570 58444
rect 376150 58380 376156 58444
rect 376220 58442 376226 58444
rect 410742 58442 410748 58444
rect 376220 58382 410748 58442
rect 376220 58380 376226 58382
rect 410742 58380 410748 58382
rect 410812 58380 410818 58444
rect 85430 58108 85436 58172
rect 85500 58108 85506 58172
rect 92422 58108 92428 58172
rect 92492 58108 92498 58172
rect 128302 58108 128308 58172
rect 128372 58108 128378 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 235942 58108 235948 58172
rect 236012 58108 236018 58172
rect 265198 58108 265204 58172
rect 265268 58108 265274 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 398230 58108 398236 58172
rect 398300 58108 398306 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 405406 58108 405412 58172
rect 405476 58108 405482 58172
rect 83958 57972 83964 58036
rect 84028 58034 84034 58036
rect 84193 58034 84259 58037
rect 84028 58032 84259 58034
rect 84028 57976 84198 58032
rect 84254 57976 84259 58032
rect 84028 57974 84259 57976
rect 84028 57972 84034 57974
rect 84193 57971 84259 57974
rect 85438 57901 85498 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78673 57898 78739 57901
rect 80421 57900 80487 57901
rect 79542 57898 79548 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 78673 57896 79548 57898
rect 78673 57840 78678 57896
rect 78734 57840 79548 57896
rect 78673 57838 79548 57840
rect 78324 57836 78330 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 78673 57835 78739 57838
rect 79542 57836 79548 57838
rect 79612 57836 79618 57900
rect 80421 57896 80468 57900
rect 80532 57898 80538 57900
rect 81433 57898 81499 57901
rect 81934 57898 81940 57900
rect 80421 57840 80426 57896
rect 80421 57836 80468 57840
rect 80532 57838 80578 57898
rect 81433 57896 81940 57898
rect 81433 57840 81438 57896
rect 81494 57840 81940 57896
rect 81433 57838 81940 57840
rect 80532 57836 80538 57838
rect 80421 57835 80487 57836
rect 81433 57835 81499 57838
rect 81934 57836 81940 57838
rect 82004 57836 82010 57900
rect 85389 57896 85498 57901
rect 85389 57840 85394 57896
rect 85450 57840 85498 57896
rect 85389 57838 85498 57840
rect 86493 57900 86559 57901
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 88333 57900 88399 57901
rect 88701 57900 88767 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 85389 57835 85455 57838
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88333 57896 88380 57900
rect 88444 57898 88450 57900
rect 88333 57840 88338 57896
rect 88333 57836 88380 57840
rect 88444 57838 88490 57898
rect 88701 57896 88748 57900
rect 88812 57898 88818 57900
rect 89713 57898 89779 57901
rect 90766 57898 90772 57900
rect 88701 57840 88706 57896
rect 88444 57836 88450 57838
rect 88701 57836 88748 57840
rect 88812 57838 88858 57898
rect 89713 57896 90772 57898
rect 89713 57840 89718 57896
rect 89774 57840 90772 57896
rect 89713 57838 90772 57840
rect 88812 57836 88818 57838
rect 88333 57835 88399 57836
rect 88701 57835 88767 57836
rect 89713 57835 89779 57838
rect 90766 57836 90772 57838
rect 90836 57836 90842 57900
rect 91093 57898 91159 57901
rect 91318 57898 91324 57900
rect 91093 57896 91324 57898
rect 91093 57840 91098 57896
rect 91154 57840 91324 57896
rect 91093 57838 91324 57840
rect 91093 57835 91159 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 91461 57898 91527 57901
rect 92430 57898 92490 58108
rect 93301 57900 93367 57901
rect 93669 57900 93735 57901
rect 98085 57900 98151 57901
rect 103789 57900 103855 57901
rect 108573 57900 108639 57901
rect 109493 57900 109559 57901
rect 112069 57900 112135 57901
rect 113173 57900 113239 57901
rect 93301 57898 93348 57900
rect 91461 57896 92490 57898
rect 91461 57840 91466 57896
rect 91522 57840 92490 57896
rect 91461 57838 92490 57840
rect 93256 57896 93348 57898
rect 93256 57840 93306 57896
rect 93256 57838 93348 57840
rect 91461 57835 91527 57838
rect 93301 57836 93348 57838
rect 93412 57836 93418 57900
rect 93669 57896 93716 57900
rect 93780 57898 93786 57900
rect 93669 57840 93674 57896
rect 93669 57836 93716 57840
rect 93780 57838 93826 57898
rect 98085 57896 98132 57900
rect 98196 57898 98202 57900
rect 98085 57840 98090 57896
rect 93780 57836 93786 57838
rect 98085 57836 98132 57840
rect 98196 57838 98242 57898
rect 103789 57896 103836 57900
rect 103900 57898 103906 57900
rect 103789 57840 103794 57896
rect 98196 57836 98202 57838
rect 103789 57836 103836 57840
rect 103900 57838 103946 57898
rect 108573 57896 108620 57900
rect 108684 57898 108690 57900
rect 108573 57840 108578 57896
rect 103900 57836 103906 57838
rect 108573 57836 108620 57840
rect 108684 57838 108730 57898
rect 109493 57896 109540 57900
rect 109604 57898 109610 57900
rect 109493 57840 109498 57896
rect 108684 57836 108690 57838
rect 109493 57836 109540 57840
rect 109604 57838 109650 57898
rect 112069 57896 112116 57900
rect 112180 57898 112186 57900
rect 112069 57840 112074 57896
rect 109604 57836 109610 57838
rect 112069 57836 112116 57840
rect 112180 57838 112226 57898
rect 113173 57896 113220 57900
rect 113284 57898 113290 57900
rect 114093 57898 114159 57901
rect 115933 57900 115999 57901
rect 114318 57898 114324 57900
rect 113173 57840 113178 57896
rect 112180 57836 112186 57838
rect 113173 57836 113220 57840
rect 113284 57838 113330 57898
rect 114093 57896 114324 57898
rect 114093 57840 114098 57896
rect 114154 57840 114324 57896
rect 114093 57838 114324 57840
rect 113284 57836 113290 57838
rect 93301 57835 93367 57836
rect 93669 57835 93735 57836
rect 98085 57835 98151 57836
rect 103789 57835 103855 57836
rect 108573 57835 108639 57836
rect 109493 57835 109559 57836
rect 112069 57835 112135 57836
rect 113173 57835 113239 57836
rect 114093 57835 114159 57838
rect 114318 57836 114324 57838
rect 114388 57836 114394 57900
rect 115933 57896 115980 57900
rect 116044 57898 116050 57900
rect 117865 57898 117931 57901
rect 119061 57900 119127 57901
rect 123477 57900 123543 57901
rect 117998 57898 118004 57900
rect 115933 57840 115938 57896
rect 115933 57836 115980 57840
rect 116044 57838 116090 57898
rect 117865 57896 118004 57898
rect 117865 57840 117870 57896
rect 117926 57840 118004 57896
rect 117865 57838 118004 57840
rect 116044 57836 116050 57838
rect 115933 57835 115999 57836
rect 117865 57835 117931 57838
rect 117998 57836 118004 57838
rect 118068 57836 118074 57900
rect 119061 57896 119108 57900
rect 119172 57898 119178 57900
rect 119061 57840 119066 57896
rect 119061 57836 119108 57840
rect 119172 57838 119218 57898
rect 123477 57896 123524 57900
rect 123588 57898 123594 57900
rect 123477 57840 123482 57896
rect 119172 57836 119178 57838
rect 123477 57836 123524 57840
rect 123588 57838 123634 57898
rect 123588 57836 123594 57838
rect 119061 57835 119127 57836
rect 123477 57835 123543 57836
rect 55070 57700 55076 57764
rect 55140 57762 55146 57764
rect 128310 57762 128370 58108
rect 153334 57901 153394 58108
rect 235950 57901 236010 58108
rect 130837 57900 130903 57901
rect 145557 57900 145623 57901
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 130837 57840 130842 57896
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 130948 57836 130954 57838
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 183461 57900 183527 57901
rect 183461 57896 183508 57900
rect 183572 57898 183578 57900
rect 183461 57840 183466 57896
rect 145668 57836 145674 57838
rect 130837 57835 130903 57836
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 183461 57836 183508 57840
rect 183572 57838 183618 57898
rect 235950 57896 236059 57901
rect 235950 57840 235998 57896
rect 236054 57840 236059 57896
rect 235950 57838 236059 57840
rect 183572 57836 183578 57838
rect 183461 57835 183527 57836
rect 235993 57835 236059 57838
rect 237373 57898 237439 57901
rect 238150 57898 238156 57900
rect 237373 57896 238156 57898
rect 237373 57840 237378 57896
rect 237434 57840 238156 57896
rect 237373 57838 238156 57840
rect 237373 57835 237439 57838
rect 238150 57836 238156 57838
rect 238220 57836 238226 57900
rect 239121 57898 239187 57901
rect 239254 57898 239260 57900
rect 239121 57896 239260 57898
rect 239121 57840 239126 57896
rect 239182 57840 239260 57896
rect 239121 57838 239260 57840
rect 239121 57835 239187 57838
rect 239254 57836 239260 57838
rect 239324 57836 239330 57900
rect 240133 57898 240199 57901
rect 241605 57900 241671 57901
rect 242893 57900 242959 57901
rect 240542 57898 240548 57900
rect 240133 57896 240548 57898
rect 240133 57840 240138 57896
rect 240194 57840 240548 57896
rect 240133 57838 240548 57840
rect 240133 57835 240199 57838
rect 240542 57836 240548 57838
rect 240612 57836 240618 57900
rect 241605 57896 241652 57900
rect 241716 57898 241722 57900
rect 241605 57840 241610 57896
rect 241605 57836 241652 57840
rect 241716 57838 241762 57898
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 242893 57840 242898 57896
rect 241716 57836 241722 57838
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 243004 57836 243010 57838
rect 244222 57836 244228 57900
rect 244292 57898 244298 57900
rect 244365 57898 244431 57901
rect 244292 57896 244431 57898
rect 244292 57840 244370 57896
rect 244426 57840 244431 57896
rect 244292 57838 244431 57840
rect 244292 57836 244298 57838
rect 241605 57835 241671 57836
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245285 57900 245351 57901
rect 245285 57896 245332 57900
rect 245396 57898 245402 57900
rect 245653 57898 245719 57901
rect 246430 57898 246436 57900
rect 245285 57840 245290 57896
rect 245285 57836 245332 57840
rect 245396 57838 245442 57898
rect 245653 57896 246436 57898
rect 245653 57840 245658 57896
rect 245714 57840 246436 57896
rect 245653 57838 246436 57840
rect 245396 57836 245402 57838
rect 245285 57835 245351 57836
rect 245653 57835 245719 57838
rect 246430 57836 246436 57838
rect 246500 57836 246506 57900
rect 247033 57898 247099 57901
rect 248597 57900 248663 57901
rect 247718 57898 247724 57900
rect 247033 57896 247724 57898
rect 247033 57840 247038 57896
rect 247094 57840 247724 57896
rect 247033 57838 247724 57840
rect 247033 57835 247099 57838
rect 247718 57836 247724 57838
rect 247788 57836 247794 57900
rect 248597 57896 248644 57900
rect 248708 57898 248714 57900
rect 249793 57898 249859 57901
rect 251173 57900 251239 57901
rect 250110 57898 250116 57900
rect 248597 57840 248602 57896
rect 248597 57836 248644 57840
rect 248708 57838 248754 57898
rect 249793 57896 250116 57898
rect 249793 57840 249798 57896
rect 249854 57840 250116 57896
rect 249793 57838 250116 57840
rect 248708 57836 248714 57838
rect 248597 57835 248663 57836
rect 249793 57835 249859 57838
rect 250110 57836 250116 57838
rect 250180 57836 250186 57900
rect 251173 57898 251220 57900
rect 251128 57896 251220 57898
rect 251128 57840 251178 57896
rect 251128 57838 251220 57840
rect 251173 57836 251220 57838
rect 251284 57836 251290 57900
rect 251357 57898 251423 57901
rect 253381 57900 253447 57901
rect 252318 57898 252324 57900
rect 251357 57896 252324 57898
rect 251357 57840 251362 57896
rect 251418 57840 252324 57896
rect 251357 57838 252324 57840
rect 251173 57835 251239 57836
rect 251357 57835 251423 57838
rect 252318 57836 252324 57838
rect 252388 57836 252394 57900
rect 253381 57896 253428 57900
rect 253492 57898 253498 57900
rect 253933 57898 253999 57901
rect 258349 57900 258415 57901
rect 254526 57898 254532 57900
rect 253381 57840 253386 57896
rect 253381 57836 253428 57840
rect 253492 57838 253538 57898
rect 253933 57896 254532 57898
rect 253933 57840 253938 57896
rect 253994 57840 254532 57896
rect 253933 57838 254532 57840
rect 253492 57836 253498 57838
rect 253381 57835 253447 57836
rect 253933 57835 253999 57838
rect 254526 57836 254532 57838
rect 254596 57836 254602 57900
rect 258349 57896 258396 57900
rect 258460 57898 258466 57900
rect 264973 57898 265039 57901
rect 265206 57898 265266 58108
rect 266353 57900 266419 57901
rect 266302 57898 266308 57900
rect 258349 57840 258354 57896
rect 258349 57836 258396 57840
rect 258460 57838 258506 57898
rect 264973 57896 265266 57898
rect 264973 57840 264978 57896
rect 265034 57840 265266 57896
rect 264973 57838 265266 57840
rect 266262 57838 266308 57898
rect 266372 57896 266419 57900
rect 266414 57840 266419 57896
rect 258460 57836 258466 57838
rect 258349 57835 258415 57836
rect 264973 57835 265039 57838
rect 266302 57836 266308 57838
rect 266372 57836 266419 57840
rect 266353 57835 266419 57836
rect 268469 57898 268535 57901
rect 271045 57900 271111 57901
rect 268694 57898 268700 57900
rect 268469 57896 268700 57898
rect 268469 57840 268474 57896
rect 268530 57840 268700 57896
rect 268469 57838 268700 57840
rect 268469 57835 268535 57838
rect 268694 57836 268700 57838
rect 268764 57836 268770 57900
rect 271045 57896 271092 57900
rect 271156 57898 271162 57900
rect 271873 57898 271939 57901
rect 272198 57898 272258 58108
rect 271045 57840 271050 57896
rect 271045 57836 271092 57840
rect 271156 57838 271202 57898
rect 271873 57896 272258 57898
rect 271873 57840 271878 57896
rect 271934 57840 272258 57896
rect 271873 57838 272258 57840
rect 273253 57900 273319 57901
rect 273253 57896 273300 57900
rect 273364 57898 273370 57900
rect 275093 57898 275159 57901
rect 275694 57898 275754 58108
rect 398238 57901 398298 58108
rect 273253 57840 273258 57896
rect 271156 57836 271162 57838
rect 271045 57835 271111 57836
rect 271873 57835 271939 57838
rect 273253 57836 273300 57840
rect 273364 57838 273410 57898
rect 275093 57896 275754 57898
rect 275093 57840 275098 57896
rect 275154 57840 275754 57896
rect 275093 57838 275754 57840
rect 283465 57898 283531 57901
rect 293309 57900 293375 57901
rect 295885 57900 295951 57901
rect 283782 57898 283788 57900
rect 283465 57896 283788 57898
rect 283465 57840 283470 57896
rect 283526 57840 283788 57896
rect 283465 57838 283788 57840
rect 273364 57836 273370 57838
rect 273253 57835 273319 57836
rect 275093 57835 275159 57838
rect 283465 57835 283531 57838
rect 283782 57836 283788 57838
rect 283852 57836 283858 57900
rect 293309 57896 293356 57900
rect 293420 57898 293426 57900
rect 293309 57840 293314 57896
rect 293309 57836 293356 57840
rect 293420 57838 293466 57898
rect 295885 57896 295932 57900
rect 295996 57898 296002 57900
rect 298093 57898 298159 57901
rect 303429 57900 303495 57901
rect 305821 57900 305887 57901
rect 310973 57900 311039 57901
rect 313365 57900 313431 57901
rect 318333 57900 318399 57901
rect 323301 57900 323367 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 298502 57898 298508 57900
rect 295885 57840 295890 57896
rect 293420 57836 293426 57838
rect 295885 57836 295932 57840
rect 295996 57838 296042 57898
rect 298093 57896 298508 57898
rect 298093 57840 298098 57896
rect 298154 57840 298508 57896
rect 298093 57838 298508 57840
rect 295996 57836 296002 57838
rect 293309 57835 293375 57836
rect 295885 57835 295951 57836
rect 298093 57835 298159 57838
rect 298502 57836 298508 57838
rect 298572 57836 298578 57900
rect 303429 57896 303476 57900
rect 303540 57898 303546 57900
rect 303429 57840 303434 57896
rect 303429 57836 303476 57840
rect 303540 57838 303586 57898
rect 305821 57896 305868 57900
rect 305932 57898 305938 57900
rect 305821 57840 305826 57896
rect 303540 57836 303546 57838
rect 305821 57836 305868 57840
rect 305932 57838 305978 57898
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 305932 57836 305938 57838
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 313365 57896 313412 57900
rect 313476 57898 313482 57900
rect 313365 57840 313370 57896
rect 311084 57836 311090 57838
rect 313365 57836 313412 57840
rect 313476 57838 313522 57898
rect 318333 57896 318380 57900
rect 318444 57898 318450 57900
rect 318333 57840 318338 57896
rect 313476 57836 313482 57838
rect 318333 57836 318380 57840
rect 318444 57838 318490 57898
rect 323301 57896 323348 57900
rect 323412 57898 323418 57900
rect 343173 57898 343220 57900
rect 323301 57840 323306 57896
rect 318444 57836 318450 57838
rect 323301 57836 323348 57840
rect 323412 57838 323458 57898
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 323412 57836 323418 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 303429 57835 303495 57836
rect 305821 57835 305887 57836
rect 310973 57835 311039 57836
rect 313365 57835 313431 57836
rect 318333 57835 318399 57836
rect 323301 57835 323367 57836
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 398189 57896 398298 57901
rect 398189 57840 398194 57896
rect 398250 57840 398298 57896
rect 398189 57838 398298 57840
rect 398833 57898 398899 57901
rect 400397 57900 400463 57901
rect 399518 57898 399524 57900
rect 398833 57896 399524 57898
rect 398833 57840 398838 57896
rect 398894 57840 399524 57896
rect 398833 57838 399524 57840
rect 398189 57835 398255 57838
rect 398833 57835 398899 57838
rect 399518 57836 399524 57838
rect 399588 57836 399594 57900
rect 400397 57896 400444 57900
rect 400508 57898 400514 57900
rect 401593 57898 401659 57901
rect 401734 57898 401794 58108
rect 400397 57840 400402 57896
rect 400397 57836 400444 57840
rect 400508 57838 400554 57898
rect 401593 57896 401794 57898
rect 401593 57840 401598 57896
rect 401654 57840 401794 57896
rect 401593 57838 401794 57840
rect 404353 57898 404419 57901
rect 405414 57898 405474 58108
rect 404353 57896 405474 57898
rect 404353 57840 404358 57896
rect 404414 57840 405474 57896
rect 404353 57838 405474 57840
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 400508 57836 400514 57838
rect 400397 57835 400463 57836
rect 401593 57835 401659 57838
rect 404353 57835 404419 57838
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407205 57898 407271 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407205 57896 407620 57898
rect 407205 57840 407210 57896
rect 407266 57840 407620 57896
rect 407205 57838 407620 57840
rect 407205 57835 407271 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 414565 57900 414631 57901
rect 415485 57900 415551 57901
rect 418429 57900 418495 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 414565 57896 414612 57900
rect 414676 57898 414682 57900
rect 414565 57840 414570 57896
rect 414565 57836 414612 57840
rect 414676 57838 414722 57898
rect 415485 57896 415532 57900
rect 415596 57898 415602 57900
rect 415485 57840 415490 57896
rect 414676 57836 414682 57838
rect 415485 57836 415532 57840
rect 415596 57838 415642 57898
rect 418429 57896 418476 57900
rect 418540 57898 418546 57900
rect 425053 57898 425119 57901
rect 426433 57900 426499 57901
rect 425278 57898 425284 57900
rect 418429 57840 418434 57896
rect 415596 57836 415602 57838
rect 418429 57836 418476 57840
rect 418540 57838 418586 57898
rect 425053 57896 425284 57898
rect 425053 57840 425058 57896
rect 425114 57840 425284 57896
rect 425053 57838 425284 57840
rect 418540 57836 418546 57838
rect 414565 57835 414631 57836
rect 415485 57835 415551 57836
rect 418429 57835 418495 57836
rect 425053 57835 425119 57838
rect 425278 57836 425284 57838
rect 425348 57836 425354 57900
rect 426382 57898 426388 57900
rect 426342 57838 426388 57898
rect 426452 57896 426499 57900
rect 427629 57900 427695 57901
rect 427629 57898 427676 57900
rect 426494 57840 426499 57896
rect 426382 57836 426388 57838
rect 426452 57836 426499 57840
rect 427584 57896 427676 57898
rect 427584 57840 427634 57896
rect 427584 57838 427676 57840
rect 426433 57835 426499 57836
rect 427629 57836 427676 57838
rect 427740 57836 427746 57900
rect 427813 57898 427879 57901
rect 428590 57898 428596 57900
rect 427813 57896 428596 57898
rect 427813 57840 427818 57896
rect 427874 57840 428596 57896
rect 427813 57838 428596 57840
rect 427629 57835 427695 57836
rect 427813 57835 427879 57838
rect 428590 57836 428596 57838
rect 428660 57836 428666 57900
rect 429193 57898 429259 57901
rect 431125 57900 431191 57901
rect 429694 57898 429700 57900
rect 429193 57896 429700 57898
rect 429193 57840 429198 57896
rect 429254 57840 429700 57896
rect 429193 57838 429700 57840
rect 429193 57835 429259 57838
rect 429694 57836 429700 57838
rect 429764 57836 429770 57900
rect 431125 57896 431172 57900
rect 431236 57898 431242 57900
rect 431953 57898 432019 57901
rect 433333 57900 433399 57901
rect 433517 57900 433583 57901
rect 435725 57900 435791 57901
rect 435909 57900 435975 57901
rect 438485 57900 438551 57901
rect 443453 57900 443519 57901
rect 445845 57900 445911 57901
rect 448237 57900 448303 57901
rect 465901 57900 465967 57901
rect 478413 57900 478479 57901
rect 485957 57900 486023 57901
rect 432270 57898 432276 57900
rect 431125 57840 431130 57896
rect 431125 57836 431172 57840
rect 431236 57838 431282 57898
rect 431953 57896 432276 57898
rect 431953 57840 431958 57896
rect 432014 57840 432276 57896
rect 431953 57838 432276 57840
rect 431236 57836 431242 57838
rect 431125 57835 431191 57836
rect 431953 57835 432019 57838
rect 432270 57836 432276 57838
rect 432340 57836 432346 57900
rect 433333 57898 433380 57900
rect 433288 57896 433380 57898
rect 433288 57840 433338 57896
rect 433288 57838 433380 57840
rect 433333 57836 433380 57838
rect 433444 57836 433450 57900
rect 433517 57896 433564 57900
rect 433628 57898 433634 57900
rect 435725 57898 435772 57900
rect 433517 57840 433522 57896
rect 433517 57836 433564 57840
rect 433628 57838 433674 57898
rect 435680 57896 435772 57898
rect 435680 57840 435730 57896
rect 435680 57838 435772 57840
rect 433628 57836 433634 57838
rect 435725 57836 435772 57838
rect 435836 57836 435842 57900
rect 435909 57896 435956 57900
rect 436020 57898 436026 57900
rect 435909 57840 435914 57896
rect 435909 57836 435956 57840
rect 436020 57838 436066 57898
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 438485 57840 438490 57896
rect 436020 57836 436026 57838
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 443453 57896 443500 57900
rect 443564 57898 443570 57900
rect 443453 57840 443458 57896
rect 438596 57836 438602 57838
rect 443453 57836 443500 57840
rect 443564 57838 443610 57898
rect 445845 57896 445892 57900
rect 445956 57898 445962 57900
rect 445845 57840 445850 57896
rect 443564 57836 443570 57838
rect 445845 57836 445892 57840
rect 445956 57838 446002 57898
rect 448237 57896 448284 57900
rect 448348 57898 448354 57900
rect 448237 57840 448242 57896
rect 445956 57836 445962 57838
rect 448237 57836 448284 57840
rect 448348 57838 448394 57898
rect 465901 57896 465948 57900
rect 466012 57898 466018 57900
rect 465901 57840 465906 57896
rect 448348 57836 448354 57838
rect 465901 57836 465948 57840
rect 466012 57838 466058 57898
rect 478413 57896 478460 57900
rect 478524 57898 478530 57900
rect 478413 57840 478418 57896
rect 466012 57836 466018 57838
rect 478413 57836 478460 57840
rect 478524 57838 478570 57898
rect 485957 57896 486004 57900
rect 486068 57898 486074 57900
rect 485957 57840 485962 57896
rect 478524 57836 478530 57838
rect 485957 57836 486004 57840
rect 486068 57838 486114 57898
rect 486068 57836 486074 57838
rect 503110 57836 503116 57900
rect 503180 57898 503186 57900
rect 503253 57898 503319 57901
rect 503529 57900 503595 57901
rect 503180 57896 503319 57898
rect 503180 57840 503258 57896
rect 503314 57840 503319 57896
rect 503180 57838 503319 57840
rect 503180 57836 503186 57838
rect 433333 57835 433399 57836
rect 433517 57835 433583 57836
rect 435725 57835 435791 57836
rect 435909 57835 435975 57836
rect 438485 57835 438551 57836
rect 443453 57835 443519 57836
rect 445845 57835 445911 57836
rect 448237 57835 448303 57836
rect 465901 57835 465967 57836
rect 478413 57835 478479 57836
rect 485957 57835 486023 57836
rect 503253 57835 503319 57838
rect 503478 57836 503484 57900
rect 503548 57898 503595 57900
rect 503548 57896 503640 57898
rect 503590 57840 503640 57896
rect 503548 57838 503640 57840
rect 503548 57836 503595 57838
rect 503529 57835 503595 57836
rect 183185 57764 183251 57765
rect 183134 57762 183140 57764
rect 55140 57702 128370 57762
rect 183094 57702 183140 57762
rect 183204 57760 183251 57764
rect 183246 57704 183251 57760
rect 55140 57700 55146 57702
rect 183134 57700 183140 57702
rect 183204 57700 183251 57704
rect 210734 57700 210740 57764
rect 210804 57762 210810 57764
rect 278446 57762 278452 57764
rect 210804 57702 278452 57762
rect 210804 57700 210810 57702
rect 278446 57700 278452 57702
rect 278516 57700 278522 57764
rect 378726 57700 378732 57764
rect 378796 57762 378802 57764
rect 470910 57762 470916 57764
rect 378796 57702 470916 57762
rect 378796 57700 378802 57702
rect 470910 57700 470916 57702
rect 470980 57700 470986 57764
rect 183185 57699 183251 57700
rect 60222 57564 60228 57628
rect 60292 57626 60298 57628
rect 125910 57626 125916 57628
rect 60292 57566 125916 57626
rect 60292 57564 60298 57566
rect 125910 57564 125916 57566
rect 125980 57564 125986 57628
rect 157333 57626 157399 57629
rect 158478 57626 158484 57628
rect 157333 57624 158484 57626
rect 157333 57568 157338 57624
rect 157394 57568 158484 57624
rect 157333 57566 158484 57568
rect 157333 57563 157399 57566
rect 158478 57564 158484 57566
rect 158548 57564 158554 57628
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 208894 57564 208900 57628
rect 208964 57626 208970 57628
rect 266445 57626 266511 57629
rect 267590 57626 267596 57628
rect 208964 57566 262908 57626
rect 208964 57564 208970 57566
rect 54702 57428 54708 57492
rect 54772 57490 54778 57492
rect 106273 57490 106339 57493
rect 106406 57490 106412 57492
rect 54772 57430 106106 57490
rect 54772 57428 54778 57430
rect 58566 57292 58572 57356
rect 58636 57354 58642 57356
rect 103830 57354 103836 57356
rect 58636 57294 103836 57354
rect 58636 57292 58642 57294
rect 103830 57292 103836 57294
rect 103900 57292 103906 57356
rect 106046 57354 106106 57430
rect 106273 57488 106412 57490
rect 106273 57432 106278 57488
rect 106334 57432 106412 57488
rect 106273 57430 106412 57432
rect 106273 57427 106339 57430
rect 106406 57428 106412 57430
rect 106476 57428 106482 57492
rect 110413 57490 110479 57493
rect 111190 57490 111196 57492
rect 110413 57488 111196 57490
rect 110413 57432 110418 57488
rect 110474 57432 111196 57488
rect 110413 57430 111196 57432
rect 110413 57427 110479 57430
rect 111190 57428 111196 57430
rect 111260 57428 111266 57492
rect 114553 57490 114619 57493
rect 115790 57490 115796 57492
rect 114553 57488 115796 57490
rect 114553 57432 114558 57488
rect 114614 57432 115796 57488
rect 114553 57430 115796 57432
rect 114553 57427 114619 57430
rect 115790 57428 115796 57430
rect 115860 57428 115866 57492
rect 116117 57490 116183 57493
rect 116894 57490 116900 57492
rect 116117 57488 116900 57490
rect 116117 57432 116122 57488
rect 116178 57432 116900 57488
rect 116117 57430 116900 57432
rect 116117 57427 116183 57430
rect 116894 57428 116900 57430
rect 116964 57428 116970 57492
rect 203190 57428 203196 57492
rect 203260 57490 203266 57492
rect 260966 57490 260972 57492
rect 203260 57430 260972 57490
rect 203260 57428 203266 57430
rect 260966 57428 260972 57430
rect 261036 57428 261042 57492
rect 262848 57490 262908 57566
rect 266445 57624 267596 57626
rect 266445 57568 266450 57624
rect 266506 57568 267596 57624
rect 266445 57566 267596 57568
rect 266445 57563 266511 57566
rect 267590 57564 267596 57566
rect 267660 57564 267666 57628
rect 269113 57626 269179 57629
rect 269798 57626 269804 57628
rect 269113 57624 269804 57626
rect 269113 57568 269118 57624
rect 269174 57568 269804 57624
rect 269113 57566 269804 57568
rect 269113 57563 269179 57566
rect 269798 57564 269804 57566
rect 269868 57564 269874 57628
rect 273345 57626 273411 57629
rect 274398 57626 274404 57628
rect 273345 57624 274404 57626
rect 273345 57568 273350 57624
rect 273406 57568 274404 57624
rect 273345 57566 274404 57568
rect 273345 57563 273411 57566
rect 274398 57564 274404 57566
rect 274468 57564 274474 57628
rect 277393 57626 277459 57629
rect 278078 57626 278084 57628
rect 277393 57624 278084 57626
rect 277393 57568 277398 57624
rect 277454 57568 278084 57624
rect 277393 57566 278084 57568
rect 277393 57563 277459 57566
rect 278078 57564 278084 57566
rect 278148 57564 278154 57628
rect 357934 57564 357940 57628
rect 358004 57626 358010 57628
rect 433241 57626 433307 57629
rect 358004 57624 433307 57626
rect 358004 57568 433246 57624
rect 433302 57568 433307 57624
rect 358004 57566 433307 57568
rect 358004 57564 358010 57566
rect 433241 57563 433307 57566
rect 433425 57626 433491 57629
rect 434662 57626 434668 57628
rect 433425 57624 434668 57626
rect 433425 57568 433430 57624
rect 433486 57568 434668 57624
rect 433425 57566 434668 57568
rect 433425 57563 433491 57566
rect 434662 57564 434668 57566
rect 434732 57564 434738 57628
rect 436093 57626 436159 57629
rect 436870 57626 436876 57628
rect 436093 57624 436876 57626
rect 436093 57568 436098 57624
rect 436154 57568 436876 57624
rect 436093 57566 436876 57568
rect 436093 57563 436159 57566
rect 436870 57564 436876 57566
rect 436940 57564 436946 57628
rect 438853 57626 438919 57629
rect 439078 57626 439084 57628
rect 438853 57624 439084 57626
rect 438853 57568 438858 57624
rect 438914 57568 439084 57624
rect 438853 57566 439084 57568
rect 438853 57563 438919 57566
rect 439078 57564 439084 57566
rect 439148 57564 439154 57628
rect 270902 57490 270908 57492
rect 262848 57430 270908 57490
rect 270902 57428 270908 57430
rect 270972 57428 270978 57492
rect 379094 57428 379100 57492
rect 379164 57490 379170 57492
rect 456374 57490 456380 57492
rect 379164 57430 456380 57490
rect 379164 57428 379170 57430
rect 456374 57428 456380 57430
rect 456444 57428 456450 57492
rect 118366 57354 118372 57356
rect 106046 57294 118372 57354
rect 118366 57292 118372 57294
rect 118436 57292 118442 57356
rect 205030 57292 205036 57356
rect 205100 57354 205106 57356
rect 255998 57354 256004 57356
rect 205100 57294 256004 57354
rect 205100 57292 205106 57294
rect 255998 57292 256004 57294
rect 256068 57292 256074 57356
rect 374494 57292 374500 57356
rect 374564 57354 374570 57356
rect 451038 57354 451044 57356
rect 374564 57294 451044 57354
rect 374564 57292 374570 57294
rect 451038 57292 451044 57294
rect 451108 57292 451114 57356
rect 58750 57156 58756 57220
rect 58820 57218 58826 57220
rect 98494 57218 98500 57220
rect 58820 57158 98500 57218
rect 58820 57156 58826 57158
rect 98494 57156 98500 57158
rect 98564 57156 98570 57220
rect 215886 57156 215892 57220
rect 215956 57218 215962 57220
rect 265934 57218 265940 57220
rect 215956 57158 265940 57218
rect 215956 57156 215962 57158
rect 265934 57156 265940 57158
rect 266004 57156 266010 57220
rect 379278 57156 379284 57220
rect 379348 57218 379354 57220
rect 430982 57218 430988 57220
rect 379348 57158 430988 57218
rect 379348 57156 379354 57158
rect 430982 57156 430988 57158
rect 431052 57156 431058 57220
rect 433241 57218 433307 57221
rect 440918 57218 440924 57220
rect 433241 57216 440924 57218
rect 433241 57160 433246 57216
rect 433302 57160 440924 57216
rect 433241 57158 440924 57160
rect 433241 57155 433307 57158
rect 440918 57156 440924 57158
rect 440988 57156 440994 57220
rect 58934 57020 58940 57084
rect 59004 57082 59010 57084
rect 96286 57082 96292 57084
rect 59004 57022 96292 57082
rect 59004 57020 59010 57022
rect 96286 57020 96292 57022
rect 96356 57020 96362 57084
rect 214414 57020 214420 57084
rect 214484 57082 214490 57084
rect 248270 57082 248276 57084
rect 214484 57022 248276 57082
rect 214484 57020 214490 57022
rect 248270 57020 248276 57022
rect 248340 57020 248346 57084
rect 378910 57020 378916 57084
rect 378980 57082 378986 57084
rect 413502 57082 413508 57084
rect 378980 57022 413508 57082
rect 378980 57020 378986 57022
rect 413502 57020 413508 57022
rect 413572 57020 413578 57084
rect 411253 56948 411319 56949
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 412541 56946 412607 56949
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 412541 56944 412650 56946
rect 412541 56888 412546 56944
rect 412602 56888 412650 56944
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 412541 56883 412650 56888
rect 412590 56813 412650 56883
rect 412590 56808 412699 56813
rect 412590 56752 412638 56808
rect 412694 56752 412699 56808
rect 412590 56750 412699 56752
rect 412633 56747 412699 56750
rect 55438 56612 55444 56676
rect 55508 56674 55514 56676
rect 133454 56674 133460 56676
rect 55508 56614 133460 56674
rect 55508 56612 55514 56614
rect 133454 56612 133460 56614
rect 133524 56612 133530 56676
rect 163262 56612 163268 56676
rect 163332 56612 163338 56676
rect 214598 56612 214604 56676
rect 214668 56674 214674 56676
rect 288198 56674 288204 56676
rect 214668 56614 288204 56674
rect 214668 56612 214674 56614
rect 288198 56612 288204 56614
rect 288268 56612 288274 56676
rect 367686 56612 367692 56676
rect 367756 56674 367762 56676
rect 460974 56674 460980 56676
rect 367756 56614 460980 56674
rect 367756 56612 367762 56614
rect 460974 56612 460980 56614
rect 461044 56612 461050 56676
rect 50654 56476 50660 56540
rect 50724 56538 50730 56540
rect 163270 56538 163330 56612
rect 50724 56478 163330 56538
rect 50724 56476 50730 56478
rect 219934 56476 219940 56540
rect 220004 56538 220010 56540
rect 421046 56538 421052 56540
rect 220004 56478 421052 56538
rect 220004 56476 220010 56478
rect 421046 56476 421052 56478
rect 421116 56476 421122 56540
rect 50470 56340 50476 56404
rect 50540 56402 50546 56404
rect 153285 56402 153351 56405
rect 50540 56400 153351 56402
rect 50540 56344 153290 56400
rect 153346 56344 153351 56400
rect 50540 56342 153351 56344
rect 50540 56340 50546 56342
rect 153285 56339 153351 56342
rect 201350 56340 201356 56404
rect 201420 56402 201426 56404
rect 273478 56402 273484 56404
rect 201420 56342 273484 56402
rect 201420 56340 201426 56342
rect 273478 56340 273484 56342
rect 273548 56340 273554 56404
rect 377254 56340 377260 56404
rect 377324 56402 377330 56404
rect 438342 56402 438348 56404
rect 377324 56342 438348 56402
rect 377324 56340 377330 56342
rect 438342 56340 438348 56342
rect 438412 56340 438418 56404
rect 55622 56204 55628 56268
rect 55692 56266 55698 56268
rect 155902 56266 155908 56268
rect 55692 56206 155908 56266
rect 55692 56204 55698 56206
rect 155902 56204 155908 56206
rect 155972 56204 155978 56268
rect 217358 56204 217364 56268
rect 217428 56266 217434 56268
rect 276974 56266 276980 56268
rect 217428 56206 276980 56266
rect 217428 56204 217434 56206
rect 276974 56204 276980 56206
rect 277044 56204 277050 56268
rect 57278 56068 57284 56132
rect 57348 56130 57354 56132
rect 119061 56130 119127 56133
rect 57348 56128 119127 56130
rect 57348 56072 119066 56128
rect 119122 56072 119127 56128
rect 57348 56070 119127 56072
rect 57348 56068 57354 56070
rect 119061 56067 119127 56070
rect 48078 55116 48084 55180
rect 48148 55178 48154 55180
rect 165613 55178 165679 55181
rect 48148 55176 165679 55178
rect 48148 55120 165618 55176
rect 165674 55120 165679 55176
rect 48148 55118 165679 55120
rect 48148 55116 48154 55118
rect 165613 55115 165679 55118
rect 214925 55178 214991 55181
rect 269113 55178 269179 55181
rect 214925 55176 269179 55178
rect 214925 55120 214930 55176
rect 214986 55120 269118 55176
rect 269174 55120 269179 55176
rect 214925 55118 269179 55120
rect 214925 55115 214991 55118
rect 269113 55115 269179 55118
rect 377806 55116 377812 55180
rect 377876 55178 377882 55180
rect 438853 55178 438919 55181
rect 377876 55176 438919 55178
rect 377876 55120 438858 55176
rect 438914 55120 438919 55176
rect 377876 55118 438919 55120
rect 377876 55116 377882 55118
rect 438853 55115 438919 55118
rect 50838 54980 50844 55044
rect 50908 55042 50914 55044
rect 157333 55042 157399 55045
rect 50908 55040 157399 55042
rect 50908 54984 157338 55040
rect 157394 54984 157399 55040
rect 50908 54982 157399 54984
rect 50908 54980 50914 54982
rect 157333 54979 157399 54982
rect 377622 54980 377628 55044
rect 377692 55042 377698 55044
rect 425053 55042 425119 55045
rect 377692 55040 425119 55042
rect 377692 54984 425058 55040
rect 425114 54984 425119 55040
rect 377692 54982 425119 54984
rect 377692 54980 377698 54982
rect 425053 54979 425119 54982
rect 53598 54844 53604 54908
rect 53668 54906 53674 54908
rect 160093 54906 160159 54909
rect 53668 54904 160159 54906
rect 53668 54848 160098 54904
rect 160154 54848 160159 54904
rect 53668 54846 160159 54848
rect 53668 54844 53674 54846
rect 160093 54843 160159 54846
rect 57830 54708 57836 54772
rect 57900 54770 57906 54772
rect 77845 54770 77911 54773
rect 57900 54768 77911 54770
rect 57900 54712 77850 54768
rect 77906 54712 77911 54768
rect 57900 54710 77911 54712
rect 57900 54708 57906 54710
rect 77845 54707 77911 54710
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 140037 4042 140103 4045
rect 210366 4042 210372 4044
rect 140037 4040 210372 4042
rect 140037 3984 140042 4040
rect 140098 3984 210372 4040
rect 140037 3982 210372 3984
rect 140037 3979 140103 3982
rect 210366 3980 210372 3982
rect 210436 3980 210442 4044
rect 129365 3906 129431 3909
rect 202086 3906 202092 3908
rect 129365 3904 202092 3906
rect 129365 3848 129370 3904
rect 129426 3848 202092 3904
rect 129365 3846 202092 3848
rect 129365 3843 129431 3846
rect 202086 3844 202092 3846
rect 202156 3844 202162 3908
rect 147121 3770 147187 3773
rect 364926 3770 364932 3772
rect 147121 3768 364932 3770
rect 147121 3712 147126 3768
rect 147182 3712 364932 3768
rect 147121 3710 364932 3712
rect 147121 3707 147187 3710
rect 364926 3708 364932 3710
rect 364996 3708 365002 3772
rect 143533 3634 143599 3637
rect 363454 3634 363460 3636
rect 143533 3632 363460 3634
rect 143533 3576 143538 3632
rect 143594 3576 363460 3632
rect 143533 3574 363460 3576
rect 143533 3571 143599 3574
rect 363454 3572 363460 3574
rect 363524 3572 363530 3636
rect 150617 3498 150683 3501
rect 375966 3498 375972 3500
rect 150617 3496 375972 3498
rect 150617 3440 150622 3496
rect 150678 3440 375972 3496
rect 150617 3438 375972 3440
rect 150617 3435 150683 3438
rect 375966 3436 375972 3438
rect 376036 3436 376042 3500
rect 132953 3362 133019 3365
rect 365110 3362 365116 3364
rect 132953 3360 365116 3362
rect 132953 3304 132958 3360
rect 133014 3304 365116 3360
rect 132953 3302 365116 3304
rect 132953 3299 133019 3302
rect 365110 3300 365116 3302
rect 365180 3300 365186 3364
rect 136449 3226 136515 3229
rect 204846 3226 204852 3228
rect 136449 3224 204852 3226
rect 136449 3168 136454 3224
rect 136510 3168 204852 3224
rect 136449 3166 204852 3168
rect 136449 3163 136515 3166
rect 204846 3164 204852 3166
rect 204916 3164 204922 3228
rect 367093 2954 367159 2957
rect 368238 2954 368244 2956
rect 367093 2952 368244 2954
rect 367093 2896 367098 2952
rect 367154 2896 368244 2952
rect 367093 2894 368244 2896
rect 367093 2891 367159 2894
rect 368238 2892 368244 2894
rect 368308 2892 368314 2956
<< via3 >>
rect 53052 639236 53116 639300
rect 51580 639100 51644 639164
rect 54340 638964 54404 639028
rect 476068 627812 476132 627876
rect 488580 627812 488644 627876
rect 506612 627812 506676 627876
rect 430620 615028 430684 615092
rect 430804 600748 430868 600812
rect 430804 527036 430868 527100
rect 430620 526900 430684 526964
rect 368244 518060 368308 518124
rect 506612 518060 506676 518124
rect 360884 489092 360948 489156
rect 364932 487732 364996 487796
rect 363460 486372 363524 486436
rect 488580 486372 488644 486436
rect 199332 485692 199396 485756
rect 366220 485692 366284 485756
rect 55076 485556 55140 485620
rect 198228 485556 198292 485620
rect 206876 485556 206940 485620
rect 209636 485556 209700 485620
rect 371924 485556 371988 485620
rect 54892 485420 54956 485484
rect 198044 485420 198108 485484
rect 371740 485420 371804 485484
rect 44956 485284 45020 485348
rect 197860 485284 197924 485348
rect 199148 485284 199212 485348
rect 370452 485284 370516 485348
rect 57836 485148 57900 485212
rect 200620 485148 200684 485212
rect 206324 485148 206388 485212
rect 219204 485148 219268 485212
rect 373764 485148 373828 485212
rect 375972 485148 376036 485212
rect 202276 485012 202340 485076
rect 217548 485012 217612 485076
rect 376156 485012 376220 485076
rect 59124 484876 59188 484940
rect 196572 484876 196636 484940
rect 198412 484876 198476 484940
rect 202460 484876 202524 484940
rect 211660 484876 211724 484940
rect 360700 484876 360764 484940
rect 59308 484740 59372 484804
rect 200988 484740 201052 484804
rect 211844 484740 211908 484804
rect 201356 484468 201420 484532
rect 206692 484468 206756 484532
rect 216996 484468 217060 484532
rect 219940 484468 220004 484532
rect 216260 483924 216324 483988
rect 213868 483788 213932 483852
rect 214420 483652 214484 483716
rect 57100 482700 57164 482764
rect 359780 482564 359844 482628
rect 212580 482428 212644 482492
rect 375420 482428 375484 482492
rect 46612 482292 46676 482356
rect 215892 482292 215956 482356
rect 374684 482292 374748 482356
rect 377260 481068 377324 481132
rect 217180 480932 217244 480996
rect 374868 480932 374932 480996
rect 203196 480796 203260 480860
rect 378732 480796 378796 480860
rect 57468 479708 57532 479772
rect 213132 479708 213196 479772
rect 359412 479708 359476 479772
rect 215340 479572 215404 479636
rect 374500 479572 374564 479636
rect 208900 479436 208964 479500
rect 210372 479436 210436 479500
rect 377444 478484 377508 478548
rect 205036 478348 205100 478412
rect 357572 478348 357636 478412
rect 214604 478212 214668 478276
rect 378916 478212 378980 478276
rect 204852 478076 204916 478140
rect 46796 476852 46860 476916
rect 213316 476852 213380 476916
rect 357940 476852 358004 476916
rect 44772 476716 44836 476780
rect 209820 476716 209884 476780
rect 379100 476716 379164 476780
rect 376892 475900 376956 475964
rect 367692 475764 367756 475828
rect 207980 475628 208044 475692
rect 379468 475628 379532 475692
rect 218652 475492 218716 475556
rect 379284 475492 379348 475556
rect 202092 475356 202156 475420
rect 218836 474268 218900 474332
rect 196756 474132 196820 474196
rect 216076 473996 216140 474060
rect 203012 472636 203076 472700
rect 204300 472500 204364 472564
rect 365116 472500 365180 472564
rect 476068 472500 476132 472564
rect 199516 471820 199580 471884
rect 217364 471684 217428 471748
rect 377628 471140 377692 471204
rect 206140 469916 206204 469980
rect 58940 469780 59004 469844
rect 200804 469780 200868 469844
rect 47900 469100 47964 469164
rect 48636 468964 48700 469028
rect 55628 468828 55692 468892
rect 53604 468692 53668 468756
rect 50476 468556 50540 468620
rect 50844 468420 50908 468484
rect 213500 468420 213564 468484
rect 359596 468420 359660 468484
rect 58756 468284 58820 468348
rect 48084 467876 48148 467940
rect 50660 467936 50724 467940
rect 50660 467880 50710 467936
rect 50710 467880 50724 467936
rect 50660 467876 50724 467880
rect 208348 467196 208412 467260
rect 60228 467060 60292 467124
rect 210004 467060 210068 467124
rect 179644 466924 179708 466988
rect 178356 466516 178420 466580
rect 190868 466576 190932 466580
rect 190868 466520 190918 466576
rect 190918 466520 190932 466576
rect 190868 466516 190932 466520
rect 338436 466576 338500 466580
rect 338436 466520 338486 466576
rect 338486 466520 338500 466576
rect 338436 466516 338500 466520
rect 339724 466576 339788 466580
rect 339724 466520 339774 466576
rect 339774 466520 339788 466576
rect 339724 466516 339788 466520
rect 350948 466576 351012 466580
rect 350948 466520 350998 466576
rect 350998 466520 351012 466576
rect 350948 466516 351012 466520
rect 498516 466516 498580 466580
rect 499804 466576 499868 466580
rect 499804 466520 499818 466576
rect 499818 466520 499868 466576
rect 499804 466516 499868 466520
rect 510844 466576 510908 466580
rect 510844 466520 510894 466576
rect 510894 466520 510908 466576
rect 510844 466516 510908 466520
rect 54708 466380 54772 466444
rect 57652 466244 57716 466308
rect 48452 466108 48516 466172
rect 53236 465972 53300 466036
rect 55444 466108 55508 466172
rect 198780 466108 198844 466172
rect 52132 465836 52196 465900
rect 205220 465836 205284 465900
rect 52316 465700 52380 465764
rect 359964 465700 360028 465764
rect 58572 465564 58636 465628
rect 51764 465156 51828 465220
rect 208164 464340 208228 464404
rect 357572 417420 357636 417484
rect 204300 413884 204364 413948
rect 208348 390628 208412 390692
rect 57652 388588 57716 388652
rect 57652 388452 57716 388516
rect 198412 380972 198476 381036
rect 210740 380972 210804 381036
rect 376892 381032 376956 381036
rect 376892 380976 376942 381032
rect 376942 380976 376956 381032
rect 376892 380972 376956 380976
rect 236054 380836 236118 380900
rect 237142 380896 237206 380900
rect 237142 380840 237158 380896
rect 237158 380840 237206 380896
rect 237142 380836 237206 380840
rect 243126 380896 243190 380900
rect 243126 380840 243138 380896
rect 243138 380840 243190 380896
rect 243126 380836 243190 380840
rect 245438 380836 245502 380900
rect 247614 380896 247678 380900
rect 247614 380840 247646 380896
rect 247646 380840 247678 380896
rect 247614 380836 247678 380840
rect 254550 380836 254614 380900
rect 255910 380896 255974 380900
rect 255910 380840 255926 380896
rect 255926 380840 255974 380896
rect 255910 380836 255974 380840
rect 256998 380896 257062 380900
rect 256998 380840 257030 380896
rect 257030 380840 257062 380896
rect 256998 380836 257062 380840
rect 76054 380700 76118 380764
rect 263934 380700 263998 380764
rect 83126 380564 83190 380628
rect 258086 380564 258150 380628
rect 259446 380624 259510 380628
rect 259446 380568 259458 380624
rect 259458 380568 259510 380624
rect 259446 380564 259510 380568
rect 260670 380564 260734 380628
rect 265294 380624 265358 380628
rect 265294 380568 265310 380624
rect 265310 380568 265358 380624
rect 265294 380564 265358 380568
rect 84516 380428 84580 380492
rect 216628 380428 216692 380492
rect 216996 380428 217060 380492
rect 105860 380352 105924 380356
rect 105860 380296 105874 380352
rect 105874 380296 105924 380352
rect 105860 380292 105924 380296
rect 111012 380352 111076 380356
rect 111012 380296 111026 380352
rect 111026 380296 111076 380352
rect 111012 380292 111076 380296
rect 113588 380352 113652 380356
rect 113588 380296 113602 380352
rect 113602 380296 113652 380352
rect 113588 380292 113652 380296
rect 115980 380352 116044 380356
rect 115980 380296 115994 380352
rect 115994 380296 116044 380352
rect 115980 380292 116044 380296
rect 118372 380352 118436 380356
rect 118372 380296 118386 380352
rect 118386 380296 118436 380352
rect 118372 380292 118436 380296
rect 120948 380352 121012 380356
rect 120948 380296 120962 380352
rect 120962 380296 121012 380352
rect 120948 380292 121012 380296
rect 123524 380352 123588 380356
rect 123524 380296 123574 380352
rect 123574 380296 123588 380352
rect 123524 380292 123588 380296
rect 128308 380352 128372 380356
rect 128308 380296 128358 380352
rect 128358 380296 128372 380352
rect 128308 380292 128372 380296
rect 133460 380352 133524 380356
rect 133460 380296 133510 380352
rect 133510 380296 133524 380352
rect 133460 380292 133524 380296
rect 135852 380352 135916 380356
rect 135852 380296 135902 380352
rect 135902 380296 135916 380352
rect 135852 380292 135916 380296
rect 138428 380352 138492 380356
rect 138428 380296 138478 380352
rect 138478 380296 138492 380352
rect 138428 380292 138492 380296
rect 148548 380352 148612 380356
rect 148548 380296 148598 380352
rect 148598 380296 148612 380352
rect 148548 380292 148612 380296
rect 155908 380352 155972 380356
rect 155908 380296 155958 380352
rect 155958 380296 155972 380352
rect 155908 380292 155972 380296
rect 158484 380352 158548 380356
rect 158484 380296 158534 380352
rect 158534 380296 158548 380352
rect 158484 380292 158548 380296
rect 160876 380352 160940 380356
rect 160876 380296 160926 380352
rect 160926 380296 160940 380352
rect 160876 380292 160940 380296
rect 163452 380352 163516 380356
rect 163452 380296 163502 380352
rect 163502 380296 163516 380352
rect 163452 380292 163516 380296
rect 166028 380352 166092 380356
rect 166028 380296 166078 380352
rect 166078 380296 166092 380352
rect 166028 380292 166092 380296
rect 244228 380352 244292 380356
rect 244228 380296 244278 380352
rect 244278 380296 244292 380352
rect 244228 380292 244292 380296
rect 119108 380156 119172 380220
rect 51764 379476 51828 379540
rect 200988 379476 201052 379540
rect 202460 379476 202524 379540
rect 206324 379476 206388 379540
rect 78260 379340 78324 379404
rect 80468 379340 80532 379404
rect 85436 379400 85500 379404
rect 85436 379344 85486 379400
rect 85486 379344 85500 379400
rect 85436 379340 85500 379344
rect 86540 379400 86604 379404
rect 86540 379344 86590 379400
rect 86590 379344 86604 379400
rect 86540 379340 86604 379344
rect 87644 379400 87708 379404
rect 87644 379344 87694 379400
rect 87694 379344 87708 379400
rect 87644 379340 87708 379344
rect 88380 379400 88444 379404
rect 88380 379344 88394 379400
rect 88394 379344 88444 379400
rect 88380 379340 88444 379344
rect 88748 379400 88812 379404
rect 88748 379344 88798 379400
rect 88798 379344 88812 379400
rect 88748 379340 88812 379344
rect 90772 379340 90836 379404
rect 91324 379400 91388 379404
rect 91324 379344 91374 379400
rect 91374 379344 91388 379400
rect 91324 379340 91388 379344
rect 92428 379400 92492 379404
rect 92428 379344 92442 379400
rect 92442 379344 92492 379400
rect 92428 379340 92492 379344
rect 93348 379340 93412 379404
rect 96108 379400 96172 379404
rect 96108 379344 96122 379400
rect 96122 379344 96172 379400
rect 96108 379340 96172 379344
rect 98500 379340 98564 379404
rect 101076 379400 101140 379404
rect 101076 379344 101090 379400
rect 101090 379344 101140 379400
rect 101076 379340 101140 379344
rect 103284 379340 103348 379404
rect 105308 379400 105372 379404
rect 105308 379344 105358 379400
rect 105358 379344 105372 379400
rect 105308 379340 105372 379344
rect 108252 379400 108316 379404
rect 108252 379344 108266 379400
rect 108266 379344 108316 379400
rect 108252 379340 108316 379344
rect 108804 379400 108868 379404
rect 108804 379344 108854 379400
rect 108854 379344 108868 379400
rect 108804 379340 108868 379344
rect 111196 379400 111260 379404
rect 111196 379344 111246 379400
rect 111246 379344 111260 379400
rect 111196 379340 111260 379344
rect 112300 379400 112364 379404
rect 112300 379344 112350 379400
rect 112350 379344 112364 379400
rect 112300 379340 112364 379344
rect 113404 379400 113468 379404
rect 113404 379344 113454 379400
rect 113454 379344 113468 379400
rect 113404 379340 113468 379344
rect 114508 379400 114572 379404
rect 114508 379344 114522 379400
rect 114522 379344 114572 379400
rect 114508 379340 114572 379344
rect 115796 379400 115860 379404
rect 115796 379344 115846 379400
rect 115846 379344 115860 379400
rect 115796 379340 115860 379344
rect 141004 379400 141068 379404
rect 141004 379344 141054 379400
rect 141054 379344 141068 379400
rect 141004 379340 141068 379344
rect 143580 379400 143644 379404
rect 143580 379344 143630 379400
rect 143630 379344 143644 379400
rect 143580 379340 143644 379344
rect 145972 379400 146036 379404
rect 145972 379344 146022 379400
rect 146022 379344 146036 379400
rect 145972 379340 146036 379344
rect 150940 379400 151004 379404
rect 150940 379344 150990 379400
rect 150990 379344 151004 379400
rect 150940 379340 151004 379344
rect 153516 379400 153580 379404
rect 153516 379344 153566 379400
rect 153566 379344 153580 379400
rect 153516 379340 153580 379344
rect 199148 379340 199212 379404
rect 79548 379204 79612 379268
rect 90036 379204 90100 379268
rect 93716 379204 93780 379268
rect 95924 379264 95988 379268
rect 95924 379208 95974 379264
rect 95974 379208 95988 379264
rect 95924 379204 95988 379208
rect 98132 379204 98196 379268
rect 99420 379264 99484 379268
rect 99420 379208 99470 379264
rect 99470 379208 99484 379264
rect 99420 379204 99484 379208
rect 102916 379264 102980 379268
rect 102916 379208 102966 379264
rect 102966 379208 102980 379264
rect 102916 379204 102980 379208
rect 109724 379204 109788 379268
rect 209820 379204 209884 379268
rect 269782 380836 269846 380900
rect 276038 380896 276102 380900
rect 276038 380840 276074 380896
rect 276074 380840 276102 380896
rect 276038 380836 276102 380840
rect 485950 380836 486014 380900
rect 421078 380760 421142 380764
rect 421078 380704 421102 380760
rect 421102 380704 421142 380760
rect 421078 380700 421142 380704
rect 421758 380760 421822 380764
rect 421758 380704 421802 380760
rect 421802 380704 421822 380760
rect 421758 380700 421822 380704
rect 425974 380760 426038 380764
rect 425974 380704 425978 380760
rect 425978 380704 426034 380760
rect 426034 380704 426038 380760
rect 425974 380700 426038 380704
rect 433590 380760 433654 380764
rect 433590 380704 433614 380760
rect 433614 380704 433654 380760
rect 433590 380700 433654 380704
rect 434406 380700 434470 380764
rect 436038 380760 436102 380764
rect 436038 380704 436062 380760
rect 436062 380704 436102 380760
rect 436038 380700 436102 380704
rect 438486 380760 438550 380764
rect 438486 380704 438490 380760
rect 438490 380704 438546 380760
rect 438546 380704 438550 380760
rect 438486 380700 438550 380704
rect 440934 380760 440998 380764
rect 440934 380704 440938 380760
rect 440938 380704 440998 380760
rect 440934 380700 440998 380704
rect 443518 380700 443582 380764
rect 271006 380624 271070 380628
rect 271006 380568 271014 380624
rect 271014 380568 271070 380624
rect 271006 380564 271070 380568
rect 408702 380624 408766 380628
rect 408702 380568 408738 380624
rect 408738 380568 408766 380624
rect 408702 380564 408766 380568
rect 413462 380624 413526 380628
rect 413462 380568 413466 380624
rect 413466 380568 413522 380624
rect 413522 380568 413526 380624
rect 413462 380564 413526 380568
rect 422846 380624 422910 380628
rect 422846 380568 422850 380624
rect 422850 380568 422906 380624
rect 422906 380568 422910 380624
rect 422846 380564 422910 380568
rect 425294 380624 425358 380628
rect 425294 380568 425298 380624
rect 425298 380568 425358 380624
rect 425294 380564 425358 380568
rect 436990 380564 437054 380628
rect 465958 380624 466022 380628
rect 465958 380568 465962 380624
rect 465962 380568 466022 380624
rect 465958 380564 466022 380568
rect 376892 379476 376956 379540
rect 268700 379400 268764 379404
rect 268700 379344 268714 379400
rect 268714 379344 268764 379400
rect 268700 379340 268764 379344
rect 271092 379400 271156 379404
rect 271092 379344 271106 379400
rect 271106 379344 271156 379400
rect 271092 379340 271156 379344
rect 272196 379340 272260 379404
rect 273300 379400 273364 379404
rect 273300 379344 273314 379400
rect 273314 379344 273364 379400
rect 273300 379340 273364 379344
rect 274404 379400 274468 379404
rect 274404 379344 274418 379400
rect 274418 379344 274468 379400
rect 274404 379340 274468 379344
rect 275692 379400 275756 379404
rect 275692 379344 275706 379400
rect 275706 379344 275756 379400
rect 275692 379340 275756 379344
rect 285996 379400 286060 379404
rect 285996 379344 286010 379400
rect 286010 379344 286060 379400
rect 285996 379340 286060 379344
rect 288204 379340 288268 379404
rect 290964 379400 291028 379404
rect 290964 379344 290978 379400
rect 290978 379344 291028 379400
rect 290964 379340 291028 379344
rect 293356 379400 293420 379404
rect 293356 379344 293370 379400
rect 293370 379344 293420 379400
rect 293356 379340 293420 379344
rect 295932 379400 295996 379404
rect 295932 379344 295946 379400
rect 295946 379344 295996 379400
rect 295932 379340 295996 379344
rect 298508 379340 298572 379404
rect 300900 379400 300964 379404
rect 300900 379344 300914 379400
rect 300914 379344 300964 379400
rect 300900 379340 300964 379344
rect 303476 379340 303540 379404
rect 305868 379340 305932 379404
rect 308444 379400 308508 379404
rect 308444 379344 308458 379400
rect 308458 379344 308508 379400
rect 308444 379340 308508 379344
rect 311020 379400 311084 379404
rect 311020 379344 311034 379400
rect 311034 379344 311084 379400
rect 311020 379340 311084 379344
rect 313412 379400 313476 379404
rect 313412 379344 313426 379400
rect 313426 379344 313476 379400
rect 313412 379340 313476 379344
rect 315804 379400 315868 379404
rect 315804 379344 315818 379400
rect 315818 379344 315868 379400
rect 315804 379340 315868 379344
rect 318380 379400 318444 379404
rect 318380 379344 318394 379400
rect 318394 379344 318444 379400
rect 318380 379340 318444 379344
rect 323348 379400 323412 379404
rect 323348 379344 323362 379400
rect 323362 379344 323412 379400
rect 323348 379340 323412 379344
rect 377444 379340 377508 379404
rect 397132 379340 397196 379404
rect 246436 379204 246500 379268
rect 248644 379264 248708 379268
rect 248644 379208 248658 379264
rect 248658 379208 248708 379264
rect 248644 379204 248708 379208
rect 250116 379264 250180 379268
rect 250116 379208 250130 379264
rect 250130 379208 250180 379264
rect 250116 379204 250180 379208
rect 251220 379264 251284 379268
rect 251220 379208 251234 379264
rect 251234 379208 251284 379264
rect 251220 379204 251284 379208
rect 252324 379264 252388 379268
rect 252324 379208 252338 379264
rect 252338 379208 252388 379264
rect 252324 379204 252388 379208
rect 253428 379264 253492 379268
rect 253428 379208 253442 379264
rect 253442 379208 253492 379264
rect 253428 379204 253492 379208
rect 261708 379264 261772 379268
rect 261708 379208 261722 379264
rect 261722 379208 261772 379264
rect 261708 379204 261772 379208
rect 273484 379264 273548 379268
rect 273484 379208 273498 379264
rect 273498 379208 273548 379264
rect 273484 379204 273548 379208
rect 276980 379264 277044 379268
rect 276980 379208 277030 379264
rect 277030 379208 277044 379264
rect 276980 379204 277044 379208
rect 278452 379204 278516 379268
rect 279188 379264 279252 379268
rect 279188 379208 279202 379264
rect 279202 379208 279252 379264
rect 279188 379204 279252 379208
rect 280844 379264 280908 379268
rect 280844 379208 280858 379264
rect 280858 379208 280908 379264
rect 280844 379204 280908 379208
rect 283420 379204 283484 379268
rect 325924 379264 325988 379268
rect 400444 379340 400508 379404
rect 406516 379340 406580 379404
rect 407620 379400 407684 379404
rect 407620 379344 407634 379400
rect 407634 379344 407684 379400
rect 407620 379340 407684 379344
rect 408356 379400 408420 379404
rect 408356 379344 408370 379400
rect 408370 379344 408420 379400
rect 408356 379340 408420 379344
rect 410748 379340 410812 379404
rect 411300 379400 411364 379404
rect 411300 379344 411314 379400
rect 411314 379344 411364 379400
rect 411300 379340 411364 379344
rect 412404 379400 412468 379404
rect 412404 379344 412418 379400
rect 412418 379344 412468 379400
rect 412404 379340 412468 379344
rect 413508 379340 413572 379404
rect 423444 379400 423508 379404
rect 423444 379344 423458 379400
rect 423458 379344 423508 379400
rect 423444 379340 423508 379344
rect 427492 379400 427556 379404
rect 427492 379344 427506 379400
rect 427506 379344 427556 379400
rect 427492 379340 427556 379344
rect 439084 379400 439148 379404
rect 439084 379344 439098 379400
rect 439098 379344 439148 379400
rect 439084 379340 439148 379344
rect 445892 379400 445956 379404
rect 445892 379344 445906 379400
rect 445906 379344 445956 379400
rect 445892 379340 445956 379344
rect 448284 379340 448348 379404
rect 451044 379400 451108 379404
rect 451044 379344 451058 379400
rect 451058 379344 451108 379400
rect 451044 379340 451108 379344
rect 453436 379340 453500 379404
rect 455828 379340 455892 379404
rect 458404 379400 458468 379404
rect 458404 379344 458418 379400
rect 458418 379344 458468 379400
rect 458404 379340 458468 379344
rect 325924 379208 325938 379264
rect 325938 379208 325988 379264
rect 325924 379204 325988 379208
rect 401732 379204 401796 379268
rect 403020 379264 403084 379268
rect 403020 379208 403034 379264
rect 403034 379208 403084 379264
rect 403020 379204 403084 379208
rect 405412 379264 405476 379268
rect 405412 379208 405426 379264
rect 405426 379208 405476 379264
rect 405412 379204 405476 379208
rect 410012 379264 410076 379268
rect 410012 379208 410026 379264
rect 410026 379208 410076 379264
rect 410012 379204 410076 379208
rect 414612 379264 414676 379268
rect 414612 379208 414626 379264
rect 414626 379208 414676 379264
rect 414612 379204 414676 379208
rect 240548 379068 240612 379132
rect 241468 379068 241532 379132
rect 415900 379204 415964 379268
rect 416084 379264 416148 379268
rect 416084 379208 416098 379264
rect 416098 379208 416148 379264
rect 416084 379204 416148 379208
rect 419396 379204 419460 379268
rect 437980 379204 438044 379268
rect 463556 379264 463620 379268
rect 463556 379208 463570 379264
rect 463570 379208 463620 379264
rect 463556 379204 463620 379208
rect 473492 379264 473556 379268
rect 473492 379208 473506 379264
rect 473506 379208 473556 379264
rect 473492 379204 473556 379208
rect 475884 379204 475948 379268
rect 480852 379264 480916 379268
rect 480852 379208 480866 379264
rect 480866 379208 480916 379264
rect 480852 379204 480916 379208
rect 503116 379264 503180 379268
rect 503116 379208 503130 379264
rect 503130 379208 503180 379264
rect 503116 379204 503180 379208
rect 503484 379264 503548 379268
rect 503484 379208 503534 379264
rect 503534 379208 503548 379264
rect 503484 379204 503548 379208
rect 57100 378932 57164 378996
rect 77156 378992 77220 378996
rect 77156 378936 77206 378992
rect 77206 378936 77220 378992
rect 77156 378932 77220 378936
rect 78260 378932 78324 378996
rect 238156 378932 238220 378996
rect 397500 378932 397564 378996
rect 53236 378796 53300 378860
rect 81940 378796 82004 378860
rect 241468 378796 241532 378860
rect 433380 379068 433444 379132
rect 418476 378796 418540 378860
rect 468524 378796 468588 378860
rect 470916 378856 470980 378860
rect 470916 378800 470930 378856
rect 470930 378800 470980 378856
rect 470916 378796 470980 378800
rect 478460 378796 478524 378860
rect 483428 378856 483492 378860
rect 483428 378800 483442 378856
rect 483442 378800 483492 378856
rect 483428 378796 483492 378800
rect 239260 378660 239324 378724
rect 94636 378584 94700 378588
rect 94636 378528 94686 378584
rect 94686 378528 94700 378584
rect 94636 378524 94700 378528
rect 97028 378524 97092 378588
rect 117084 378524 117148 378588
rect 210004 378524 210068 378588
rect 278084 378524 278148 378588
rect 320956 378584 321020 378588
rect 320956 378528 320970 378584
rect 320970 378528 321020 378584
rect 320956 378524 321020 378528
rect 100708 378448 100772 378452
rect 100708 378392 100758 378448
rect 100758 378392 100772 378448
rect 100708 378388 100772 378392
rect 104020 378448 104084 378452
rect 104020 378392 104070 378448
rect 104070 378392 104084 378448
rect 104020 378388 104084 378392
rect 125916 378448 125980 378452
rect 125916 378392 125966 378448
rect 125966 378392 125980 378448
rect 125916 378388 125980 378392
rect 131068 378448 131132 378452
rect 131068 378392 131082 378448
rect 131082 378392 131132 378448
rect 131068 378388 131132 378392
rect 183140 378388 183204 378452
rect 248276 378448 248340 378452
rect 248276 378392 248290 378448
rect 248290 378392 248340 378448
rect 248276 378388 248340 378392
rect 250668 378448 250732 378452
rect 250668 378392 250682 378448
rect 250682 378392 250732 378448
rect 250668 378388 250732 378392
rect 253612 378448 253676 378452
rect 253612 378392 253626 378448
rect 253626 378392 253676 378448
rect 253612 378388 253676 378392
rect 256004 378448 256068 378452
rect 256004 378392 256018 378448
rect 256018 378392 256068 378448
rect 256004 378388 256068 378392
rect 258396 378448 258460 378452
rect 258396 378392 258410 378448
rect 258410 378392 258460 378448
rect 258396 378388 258460 378392
rect 260972 378448 261036 378452
rect 260972 378392 260986 378448
rect 260986 378392 261036 378448
rect 260972 378388 261036 378392
rect 263548 378448 263612 378452
rect 263548 378392 263598 378448
rect 263598 378392 263612 378448
rect 263548 378388 263612 378392
rect 265940 378388 266004 378452
rect 268332 378388 268396 378452
rect 343220 378448 343284 378452
rect 377628 378660 377692 378724
rect 435772 378660 435836 378724
rect 396028 378584 396092 378588
rect 396028 378528 396078 378584
rect 396078 378528 396092 378584
rect 396028 378524 396092 378528
rect 404124 378524 404188 378588
rect 428228 378584 428292 378588
rect 428228 378528 428242 378584
rect 428242 378528 428292 378584
rect 428228 378524 428292 378528
rect 430988 378524 431052 378588
rect 343220 378392 343234 378448
rect 343234 378392 343284 378448
rect 343220 378388 343284 378392
rect 399524 378388 399588 378452
rect 101812 378252 101876 378316
rect 118188 378252 118252 378316
rect 241836 378252 241900 378316
rect 262812 378312 262876 378316
rect 262812 378256 262826 378312
rect 262826 378256 262876 378312
rect 262812 378252 262876 378256
rect 266308 378312 266372 378316
rect 266308 378256 266358 378312
rect 266358 378256 266372 378312
rect 266308 378252 266372 378256
rect 267596 378312 267660 378316
rect 267596 378256 267610 378312
rect 267610 378256 267660 378312
rect 267596 378252 267660 378256
rect 343404 378252 343468 378316
rect 428596 378252 428660 378316
rect 106412 378176 106476 378180
rect 106412 378120 106462 378176
rect 106462 378120 106476 378176
rect 106412 378116 106476 378120
rect 107516 378176 107580 378180
rect 107516 378120 107566 378176
rect 107566 378120 107580 378176
rect 107516 378116 107580 378120
rect 183508 378116 183572 378180
rect 377996 378116 378060 378180
rect 417004 378176 417068 378180
rect 417004 378120 417018 378176
rect 417018 378120 417068 378176
rect 417004 378116 417068 378120
rect 418108 378176 418172 378180
rect 418108 378120 418158 378176
rect 418158 378120 418172 378176
rect 418108 378116 418172 378120
rect 420684 378116 420748 378180
rect 423996 378176 424060 378180
rect 423996 378120 424010 378176
rect 424010 378120 424060 378176
rect 423996 378116 424060 378120
rect 426388 378176 426452 378180
rect 426388 378120 426438 378176
rect 426438 378120 426452 378176
rect 426388 378116 426452 378120
rect 429700 378116 429764 378180
rect 431172 378176 431236 378180
rect 431172 378120 431186 378176
rect 431186 378120 431236 378176
rect 431172 378116 431236 378120
rect 432276 378176 432340 378180
rect 432276 378120 432290 378176
rect 432290 378120 432340 378176
rect 432276 378116 432340 378120
rect 460980 378116 461044 378180
rect 359780 377980 359844 378044
rect 211844 377844 211908 377908
rect 212580 377844 212644 377908
rect 215340 377844 215404 377908
rect 211660 376620 211724 376684
rect 213868 376620 213932 376684
rect 216628 376620 216692 376684
rect 377260 376620 377324 376684
rect 217548 375260 217612 375324
rect 217548 375048 217612 375052
rect 217548 374992 217562 375048
rect 217562 374992 217612 375048
rect 217548 374988 217612 374992
rect 359964 374580 360028 374644
rect 178540 358864 178604 358868
rect 178540 358808 178590 358864
rect 178590 358808 178604 358864
rect 178540 358804 178604 358808
rect 179644 358864 179708 358868
rect 179644 358808 179694 358864
rect 179694 358808 179708 358864
rect 179644 358804 179708 358808
rect 190868 358864 190932 358868
rect 190868 358808 190918 358864
rect 190918 358808 190932 358864
rect 190868 358804 190932 358808
rect 338436 358864 338500 358868
rect 338436 358808 338486 358864
rect 338486 358808 338500 358864
rect 338436 358804 338500 358808
rect 339724 358804 339788 358868
rect 350948 358804 351012 358868
rect 498516 358804 498580 358868
rect 499804 358804 499868 358868
rect 510844 358864 510908 358868
rect 510844 358808 510894 358864
rect 510894 358808 510908 358864
rect 510844 358804 510908 358808
rect 54340 304948 54404 305012
rect 376892 274620 376956 274684
rect 95910 273804 95974 273868
rect 266382 273728 266446 273732
rect 266382 273672 266414 273728
rect 266414 273672 266446 273728
rect 266382 273668 266446 273672
rect 278078 273728 278142 273732
rect 278078 273672 278098 273728
rect 278098 273672 278142 273728
rect 278078 273668 278142 273672
rect 111006 273592 111070 273596
rect 111006 273536 111026 273592
rect 111026 273536 111070 273592
rect 111006 273532 111070 273536
rect 133446 273592 133510 273596
rect 133446 273536 133474 273592
rect 133474 273536 133510 273592
rect 133446 273532 133510 273536
rect 135894 273592 135958 273596
rect 135894 273536 135902 273592
rect 135902 273536 135958 273592
rect 135894 273532 135958 273536
rect 138478 273592 138542 273596
rect 138478 273536 138534 273592
rect 138534 273536 138542 273592
rect 138478 273532 138542 273536
rect 140926 273532 140990 273596
rect 250742 273592 250806 273596
rect 250742 273536 250774 273592
rect 250774 273536 250806 273592
rect 250742 273532 250806 273536
rect 273318 273592 273382 273596
rect 273318 273536 273350 273592
rect 273350 273536 273382 273592
rect 273318 273532 273382 273536
rect 275766 273592 275830 273596
rect 275766 273536 275798 273592
rect 275798 273536 275830 273592
rect 275766 273532 275830 273536
rect 283518 273592 283582 273596
rect 283518 273536 283526 273592
rect 283526 273536 283582 273592
rect 283518 273532 283582 273536
rect 421078 273592 421142 273596
rect 421078 273536 421102 273592
rect 421102 273536 421142 273592
rect 421078 273532 421142 273536
rect 450998 273592 451062 273596
rect 450998 273536 451002 273592
rect 451002 273536 451058 273592
rect 451058 273536 451062 273592
rect 450998 273532 451062 273536
rect 376892 273396 376956 273460
rect 422892 273396 422956 273460
rect 218836 273260 218900 273324
rect 285996 273320 286060 273324
rect 285996 273264 286010 273320
rect 286010 273264 286060 273320
rect 285996 273260 286060 273264
rect 359412 273260 359476 273324
rect 430988 273396 431052 273460
rect 423444 273320 423508 273324
rect 423444 273264 423458 273320
rect 423458 273264 423508 273320
rect 423444 273260 423508 273264
rect 423812 273320 423876 273324
rect 423812 273264 423826 273320
rect 423826 273264 423876 273320
rect 423812 273260 423876 273264
rect 426388 273320 426452 273324
rect 426388 273264 426438 273320
rect 426438 273264 426452 273320
rect 426388 273260 426452 273264
rect 100708 273184 100772 273188
rect 100708 273128 100758 273184
rect 100758 273128 100772 273184
rect 100708 273124 100772 273128
rect 199332 273124 199396 273188
rect 318380 273124 318444 273188
rect 359596 273124 359660 273188
rect 486004 273124 486068 273188
rect 102732 272988 102796 273052
rect 196572 272988 196636 273052
rect 311020 272988 311084 273052
rect 483244 272988 483308 273052
rect 76052 272912 76116 272916
rect 76052 272856 76066 272912
rect 76066 272856 76116 272912
rect 76052 272852 76116 272856
rect 90772 272912 90836 272916
rect 90772 272856 90786 272912
rect 90786 272856 90836 272912
rect 90772 272852 90836 272856
rect 93716 272912 93780 272916
rect 93716 272856 93730 272912
rect 93730 272856 93780 272912
rect 93716 272852 93780 272856
rect 95924 272912 95988 272916
rect 95924 272856 95938 272912
rect 95938 272856 95988 272912
rect 95924 272852 95988 272856
rect 98500 272912 98564 272916
rect 98500 272856 98514 272912
rect 98514 272856 98564 272912
rect 98500 272852 98564 272856
rect 99420 272912 99484 272916
rect 99420 272856 99434 272912
rect 99434 272856 99484 272912
rect 99420 272852 99484 272856
rect 199516 272852 199580 272916
rect 288204 272912 288268 272916
rect 288204 272856 288218 272912
rect 288218 272856 288268 272912
rect 288204 272852 288268 272856
rect 290964 272912 291028 272916
rect 290964 272856 290978 272912
rect 290978 272856 291028 272912
rect 290964 272852 291028 272856
rect 293356 272912 293420 272916
rect 293356 272856 293370 272912
rect 293370 272856 293420 272912
rect 293356 272852 293420 272856
rect 300900 272912 300964 272916
rect 300900 272856 300914 272912
rect 300914 272856 300964 272912
rect 300900 272852 300964 272856
rect 480852 272852 480916 272916
rect 103836 272716 103900 272780
rect 217364 272716 217428 272780
rect 298508 272776 298572 272780
rect 298508 272720 298522 272776
rect 298522 272720 298572 272776
rect 118004 272580 118068 272644
rect 143580 272640 143644 272644
rect 143580 272584 143594 272640
rect 143594 272584 143644 272640
rect 143580 272580 143644 272584
rect 295932 272580 295996 272644
rect 298508 272716 298572 272720
rect 426020 272776 426084 272780
rect 426020 272720 426034 272776
rect 426034 272720 426084 272776
rect 426020 272716 426084 272720
rect 428228 272776 428292 272780
rect 428228 272720 428242 272776
rect 428242 272720 428292 272776
rect 428228 272716 428292 272720
rect 431172 272776 431236 272780
rect 431172 272720 431186 272776
rect 431186 272720 431236 272776
rect 431172 272716 431236 272720
rect 468524 272776 468588 272780
rect 468524 272720 468538 272776
rect 468538 272720 468588 272776
rect 468524 272716 468588 272720
rect 470916 272776 470980 272780
rect 470916 272720 470930 272776
rect 470930 272720 470980 272776
rect 470916 272716 470980 272720
rect 473492 272776 473556 272780
rect 473492 272720 473506 272776
rect 473506 272720 473556 272776
rect 473492 272716 473556 272720
rect 303476 272580 303540 272644
rect 305868 272640 305932 272644
rect 305868 272584 305882 272640
rect 305882 272584 305932 272640
rect 305868 272580 305932 272584
rect 320956 272640 321020 272644
rect 320956 272584 320970 272640
rect 320970 272584 321020 272640
rect 320956 272580 321020 272584
rect 475884 272640 475948 272644
rect 475884 272584 475898 272640
rect 475898 272584 475948 272640
rect 475884 272580 475948 272584
rect 478460 272640 478524 272644
rect 478460 272584 478474 272640
rect 478474 272584 478524 272640
rect 478460 272580 478524 272584
rect 119108 272444 119172 272508
rect 97028 272368 97092 272372
rect 97028 272312 97042 272368
rect 97042 272312 97092 272368
rect 97028 272308 97092 272312
rect 113588 272232 113652 272236
rect 113588 272176 113602 272232
rect 113602 272176 113652 272232
rect 113588 272172 113652 272176
rect 235948 272232 236012 272236
rect 235948 272176 235998 272232
rect 235998 272176 236012 272232
rect 235948 272172 236012 272176
rect 265204 272232 265268 272236
rect 265204 272176 265218 272232
rect 265218 272176 265268 272232
rect 265204 272172 265268 272176
rect 401732 272232 401796 272236
rect 401732 272176 401746 272232
rect 401746 272176 401796 272232
rect 401732 272172 401796 272176
rect 416084 272232 416148 272236
rect 416084 272176 416098 272232
rect 416098 272176 416148 272232
rect 416084 272172 416148 272176
rect 437980 272232 438044 272236
rect 437980 272176 437994 272232
rect 437994 272176 438044 272232
rect 437980 272172 438044 272176
rect 455828 272232 455892 272236
rect 455828 272176 455842 272232
rect 455842 272176 455892 272232
rect 455828 272172 455892 272176
rect 77156 271764 77220 271828
rect 83044 271764 83108 271828
rect 83964 271764 84028 271828
rect 87644 271764 87708 271828
rect 94452 271764 94516 271828
rect 98132 271764 98196 271828
rect 101812 271764 101876 271828
rect 114508 271824 114572 271828
rect 114508 271768 114522 271824
rect 114522 271768 114572 271824
rect 114508 271764 114572 271768
rect 123524 271764 123588 271828
rect 128676 271764 128740 271828
rect 130884 271764 130948 271828
rect 150940 271764 151004 271828
rect 154068 271764 154132 271828
rect 155908 271764 155972 271828
rect 196756 271764 196820 271828
rect 268700 271764 268764 271828
rect 270908 271764 270972 271828
rect 276244 271764 276308 271828
rect 280844 271764 280908 271828
rect 308628 271764 308692 271828
rect 313412 271764 313476 271828
rect 343404 271764 343468 271828
rect 403020 271824 403084 271828
rect 403020 271768 403034 271824
rect 403034 271768 403084 271824
rect 403020 271764 403084 271768
rect 418476 271764 418540 271828
rect 433564 271764 433628 271828
rect 435956 271764 436020 271828
rect 438532 271764 438596 271828
rect 445892 271764 445956 271828
rect 448284 271764 448348 271828
rect 453436 271764 453500 271828
rect 458404 271764 458468 271828
rect 81940 271628 82004 271692
rect 84700 271688 84764 271692
rect 84700 271632 84714 271688
rect 84714 271632 84764 271688
rect 84700 271628 84764 271632
rect 103836 271628 103900 271692
rect 120764 271628 120828 271692
rect 125916 271628 125980 271692
rect 158484 271628 158548 271692
rect 160876 271628 160940 271692
rect 163452 271628 163516 271692
rect 166028 271628 166092 271692
rect 198780 271628 198844 271692
rect 315068 271628 315132 271692
rect 465948 271628 466012 271692
rect 503116 271628 503180 271692
rect 80468 271492 80532 271556
rect 115980 271552 116044 271556
rect 115980 271496 115994 271552
rect 115994 271496 116044 271552
rect 115980 271492 116044 271496
rect 118372 271492 118436 271556
rect 217180 271492 217244 271556
rect 101076 271356 101140 271420
rect 105860 271356 105924 271420
rect 183140 271356 183204 271420
rect 237052 271356 237116 271420
rect 258396 271492 258460 271556
rect 263548 271552 263612 271556
rect 263548 271496 263598 271552
rect 263598 271496 263612 271552
rect 263548 271492 263612 271496
rect 265940 271492 266004 271556
rect 268332 271492 268396 271556
rect 272564 271492 272628 271556
rect 276980 271492 277044 271556
rect 343220 271492 343284 271556
rect 460980 271492 461044 271556
rect 273484 271356 273548 271420
rect 278452 271356 278516 271420
rect 377812 271356 377876 271420
rect 253612 271220 253676 271284
rect 260972 271220 261036 271284
rect 78260 271084 78324 271148
rect 88380 271144 88444 271148
rect 88380 271088 88394 271144
rect 88394 271088 88444 271144
rect 88380 271084 88444 271088
rect 183508 271144 183572 271148
rect 183508 271088 183522 271144
rect 183522 271088 183572 271144
rect 183508 271084 183572 271088
rect 248276 271084 248340 271148
rect 256188 271084 256252 271148
rect 79548 270948 79612 271012
rect 88748 270948 88812 271012
rect 90036 270948 90100 271012
rect 107516 270948 107580 271012
rect 108620 270948 108684 271012
rect 112116 270948 112180 271012
rect 325556 270948 325620 271012
rect 396028 271220 396092 271284
rect 415532 271356 415596 271420
rect 440924 271356 440988 271420
rect 413692 271220 413756 271284
rect 439268 271220 439332 271284
rect 443500 271220 443564 271284
rect 503484 271220 503548 271284
rect 410748 271084 410812 271148
rect 414428 271084 414492 271148
rect 417004 271084 417068 271148
rect 434668 271084 434732 271148
rect 405044 270948 405108 271012
rect 408172 270948 408236 271012
rect 412404 270948 412468 271012
rect 428596 270948 428660 271012
rect 429700 270948 429764 271012
rect 433380 270948 433444 271012
rect 435772 270948 435836 271012
rect 86540 270812 86604 270876
rect 93348 270812 93412 270876
rect 105308 270812 105372 270876
rect 106412 270812 106476 270876
rect 254532 270812 254596 270876
rect 279004 270812 279068 270876
rect 462636 270812 462700 270876
rect 111196 270676 111260 270740
rect 244228 270676 244292 270740
rect 252324 270676 252388 270740
rect 255820 270676 255884 270740
rect 260604 270676 260668 270740
rect 413324 270676 413388 270740
rect 419212 270676 419276 270740
rect 427676 270676 427740 270740
rect 91324 270540 91388 270604
rect 108252 270540 108316 270604
rect 109540 270540 109604 270604
rect 113220 270600 113284 270604
rect 113220 270544 113234 270600
rect 113234 270544 113284 270600
rect 113220 270540 113284 270544
rect 115796 270600 115860 270604
rect 115796 270544 115846 270600
rect 115846 270544 115860 270600
rect 115796 270540 115860 270544
rect 117084 270540 117148 270604
rect 145604 270540 145668 270604
rect 148548 270540 148612 270604
rect 239260 270540 239324 270604
rect 242940 270600 243004 270604
rect 242940 270544 242954 270600
rect 242954 270544 243004 270600
rect 242940 270540 243004 270544
rect 245332 270540 245396 270604
rect 246436 270540 246500 270604
rect 247724 270540 247788 270604
rect 248644 270540 248708 270604
rect 250116 270540 250180 270604
rect 251220 270600 251284 270604
rect 251220 270544 251234 270600
rect 251234 270544 251284 270600
rect 251220 270540 251284 270544
rect 253428 270540 253492 270604
rect 256924 270540 256988 270604
rect 258396 270540 258460 270604
rect 259500 270600 259564 270604
rect 259500 270544 259514 270600
rect 259514 270544 259564 270600
rect 259500 270540 259564 270544
rect 262076 270540 262140 270604
rect 262812 270540 262876 270604
rect 263916 270540 263980 270604
rect 267596 270540 267660 270604
rect 269804 270540 269868 270604
rect 271276 270540 271340 270604
rect 274404 270540 274468 270604
rect 397132 270540 397196 270604
rect 397500 270600 397564 270604
rect 397500 270544 397514 270600
rect 397514 270544 397564 270600
rect 397500 270540 397564 270544
rect 399524 270540 399588 270604
rect 400444 270540 400508 270604
rect 404124 270540 404188 270604
rect 406516 270540 406580 270604
rect 407620 270540 407684 270604
rect 408724 270540 408788 270604
rect 410012 270540 410076 270604
rect 411300 270600 411364 270604
rect 411300 270544 411350 270600
rect 411350 270544 411364 270600
rect 411300 270540 411364 270544
rect 418108 270600 418172 270604
rect 418108 270544 418158 270600
rect 418158 270544 418172 270600
rect 418108 270540 418172 270544
rect 420684 270540 420748 270604
rect 421788 270540 421852 270604
rect 436876 270540 436940 270604
rect 57468 270268 57532 270332
rect 91508 270404 91572 270468
rect 323348 270404 323412 270468
rect 241652 270268 241716 270332
rect 240548 270132 240612 270196
rect 432276 270404 432340 270468
rect 425284 270268 425348 270332
rect 238156 269724 238220 269788
rect 375420 269044 375484 269108
rect 44772 268364 44836 268428
rect 217548 268364 217612 268428
rect 46612 267684 46676 267748
rect 53052 253948 53116 254012
rect 190868 253676 190932 253740
rect 339724 253404 339788 253468
rect 499804 253268 499868 253332
rect 178540 253132 178604 253196
rect 179644 253132 179708 253196
rect 350948 253132 351012 253196
rect 338436 252996 338500 253060
rect 498516 252724 498580 252788
rect 510844 252648 510908 252652
rect 510844 252592 510894 252648
rect 510894 252592 510908 252648
rect 510844 252588 510908 252592
rect 57468 252452 57532 252516
rect 57284 252316 57348 252380
rect 217548 251772 217612 251836
rect 377996 251772 378060 251836
rect 46796 251092 46860 251156
rect 51580 201452 51644 201516
rect 57652 175068 57716 175132
rect 57836 166908 57900 166972
rect 198228 166908 198292 166972
rect 101078 166832 101142 166836
rect 101078 166776 101090 166832
rect 101090 166776 101142 166832
rect 101078 166772 101142 166776
rect 103526 166832 103590 166836
rect 103526 166776 103574 166832
rect 103574 166776 103590 166832
rect 103526 166772 103590 166776
rect 108286 166832 108350 166836
rect 108286 166776 108302 166832
rect 108302 166776 108350 166832
rect 108286 166772 108350 166776
rect 138478 166832 138542 166836
rect 138478 166776 138534 166832
rect 138534 166776 138542 166832
rect 138478 166772 138542 166776
rect 140926 166772 140990 166836
rect 143510 166772 143574 166836
rect 145958 166832 146022 166836
rect 145958 166776 145986 166832
rect 145986 166776 146022 166832
rect 145958 166772 146022 166776
rect 213500 166772 213564 166836
rect 303510 166772 303574 166836
rect 313438 166772 313502 166836
rect 418476 166832 418540 166836
rect 418476 166776 418490 166832
rect 418490 166776 418540 166832
rect 418476 166772 418540 166776
rect 421052 166832 421116 166836
rect 421052 166776 421066 166832
rect 421066 166776 421116 166832
rect 421052 166772 421116 166776
rect 423444 166832 423508 166836
rect 423444 166776 423458 166832
rect 423458 166776 423508 166832
rect 423444 166772 423508 166776
rect 445892 166832 445956 166836
rect 445892 166776 445906 166832
rect 445906 166776 445956 166832
rect 445892 166772 445956 166776
rect 470990 166832 471054 166836
rect 470990 166776 471022 166832
rect 471022 166776 471054 166832
rect 470990 166772 471054 166776
rect 473438 166832 473502 166836
rect 473438 166776 473450 166832
rect 473450 166776 473502 166832
rect 473438 166772 473502 166776
rect 475886 166832 475950 166836
rect 475886 166776 475898 166832
rect 475898 166776 475950 166832
rect 475886 166772 475950 166776
rect 478470 166832 478534 166836
rect 478470 166776 478474 166832
rect 478474 166776 478534 166832
rect 478470 166772 478534 166776
rect 480918 166832 480982 166836
rect 480918 166776 480958 166832
rect 480958 166776 480982 166832
rect 480918 166772 480982 166776
rect 148548 166696 148612 166700
rect 148548 166640 148562 166696
rect 148562 166640 148612 166696
rect 148548 166636 148612 166640
rect 163366 166696 163430 166700
rect 163366 166640 163374 166696
rect 163374 166640 163430 166696
rect 163366 166636 163430 166640
rect 165950 166636 166014 166700
rect 205220 166636 205284 166700
rect 107606 166560 107670 166564
rect 107606 166504 107658 166560
rect 107658 166504 107670 166560
rect 107606 166500 107670 166504
rect 150940 166560 151004 166564
rect 150940 166504 150954 166560
rect 150954 166504 151004 166560
rect 150940 166500 151004 166504
rect 153332 166560 153396 166564
rect 153332 166504 153346 166560
rect 153346 166504 153396 166560
rect 153332 166500 153396 166504
rect 183222 166560 183286 166564
rect 183222 166504 183282 166560
rect 183282 166504 183286 166560
rect 183222 166500 183286 166504
rect 260972 166560 261036 166564
rect 260972 166504 260986 166560
rect 260986 166504 261036 166560
rect 260972 166500 261036 166504
rect 265940 166560 266004 166564
rect 265940 166504 265954 166560
rect 265954 166504 266004 166560
rect 265940 166500 266004 166504
rect 270908 166560 270972 166564
rect 270908 166504 270922 166560
rect 270922 166504 270972 166560
rect 270908 166500 270972 166504
rect 285966 166696 286030 166700
rect 285966 166640 286010 166696
rect 286010 166640 286030 166696
rect 285966 166636 286030 166640
rect 290998 166696 291062 166700
rect 290998 166640 291014 166696
rect 291014 166640 291062 166696
rect 290998 166636 291062 166640
rect 293446 166696 293510 166700
rect 293446 166640 293462 166696
rect 293462 166640 293510 166696
rect 293446 166636 293510 166640
rect 295894 166696 295958 166700
rect 295894 166640 295946 166696
rect 295946 166640 295958 166696
rect 295894 166636 295958 166640
rect 298478 166696 298542 166700
rect 298478 166640 298522 166696
rect 298522 166640 298542 166696
rect 298478 166636 298542 166640
rect 305958 166696 306022 166700
rect 305958 166640 305974 166696
rect 305974 166640 306022 166696
rect 305958 166636 306022 166640
rect 483366 166696 483430 166700
rect 483366 166640 483386 166696
rect 483386 166640 483430 166696
rect 483366 166636 483430 166640
rect 485950 166696 486014 166700
rect 485950 166640 485962 166696
rect 485962 166640 486014 166696
rect 485950 166636 486014 166640
rect 288278 166500 288342 166564
rect 503222 166560 503286 166564
rect 503222 166504 503258 166560
rect 503258 166504 503286 166560
rect 503222 166500 503286 166504
rect 96108 166288 96172 166292
rect 96108 166232 96122 166288
rect 96122 166232 96172 166288
rect 96108 166228 96172 166232
rect 98500 166288 98564 166292
rect 98500 166232 98514 166288
rect 98514 166232 98564 166288
rect 98500 166228 98564 166232
rect 428228 166288 428292 166292
rect 428228 166232 428242 166288
rect 428242 166232 428292 166288
rect 428228 166228 428292 166232
rect 430988 166288 431052 166292
rect 430988 166232 431002 166288
rect 431002 166232 431052 166288
rect 430988 166228 431052 166232
rect 81756 165548 81820 165612
rect 85436 165548 85500 165612
rect 92428 165548 92492 165612
rect 95740 165548 95804 165612
rect 99420 165608 99484 165612
rect 99420 165552 99434 165608
rect 99434 165552 99484 165608
rect 99420 165548 99484 165552
rect 100708 165548 100772 165612
rect 105308 165548 105372 165612
rect 105860 165548 105924 165612
rect 106412 165608 106476 165612
rect 106412 165552 106426 165608
rect 106426 165552 106476 165608
rect 106412 165548 106476 165552
rect 108620 165548 108684 165612
rect 109724 165608 109788 165612
rect 109724 165552 109738 165608
rect 109738 165552 109788 165608
rect 109724 165548 109788 165552
rect 111012 165608 111076 165612
rect 111012 165552 111026 165608
rect 111026 165552 111076 165608
rect 111012 165548 111076 165552
rect 112116 165548 112180 165612
rect 113588 165608 113652 165612
rect 113588 165552 113602 165608
rect 113602 165552 113652 165608
rect 113588 165548 113652 165552
rect 115980 165608 116044 165612
rect 115980 165552 115994 165608
rect 115994 165552 116044 165608
rect 115980 165548 116044 165552
rect 118004 165548 118068 165612
rect 118372 165608 118436 165612
rect 118372 165552 118386 165608
rect 118386 165552 118436 165608
rect 118372 165548 118436 165552
rect 119108 165608 119172 165612
rect 119108 165552 119122 165608
rect 119122 165552 119172 165608
rect 119108 165548 119172 165552
rect 120948 165608 121012 165612
rect 120948 165552 120962 165608
rect 120962 165552 121012 165608
rect 120948 165548 121012 165552
rect 123524 165608 123588 165612
rect 123524 165552 123538 165608
rect 123538 165552 123588 165608
rect 123524 165548 123588 165552
rect 125916 165608 125980 165612
rect 125916 165552 125930 165608
rect 125930 165552 125980 165608
rect 125916 165548 125980 165552
rect 128492 165548 128556 165612
rect 130884 165548 130948 165612
rect 133460 165548 133524 165612
rect 183324 165608 183388 165612
rect 183324 165552 183374 165608
rect 183374 165552 183388 165608
rect 183324 165548 183388 165552
rect 235948 165608 236012 165612
rect 235948 165552 235998 165608
rect 235998 165552 236012 165608
rect 235948 165548 236012 165552
rect 239628 165548 239692 165612
rect 243124 165548 243188 165612
rect 247540 165548 247604 165612
rect 248276 165548 248340 165612
rect 250668 165548 250732 165612
rect 253612 165548 253676 165612
rect 258396 165548 258460 165612
rect 261708 165548 261772 165612
rect 265204 165548 265268 165612
rect 266492 165548 266556 165612
rect 268332 165548 268396 165612
rect 280844 165548 280908 165612
rect 283420 165608 283484 165612
rect 283420 165552 283434 165608
rect 283434 165552 283484 165608
rect 283420 165548 283484 165552
rect 300900 165608 300964 165612
rect 300900 165552 300914 165608
rect 300914 165552 300964 165608
rect 300900 165548 300964 165552
rect 308444 165608 308508 165612
rect 308444 165552 308458 165608
rect 308458 165552 308508 165608
rect 308444 165548 308508 165552
rect 323348 165548 323412 165612
rect 325924 165608 325988 165612
rect 325924 165552 325938 165608
rect 325938 165552 325988 165608
rect 325924 165548 325988 165552
rect 343220 165608 343284 165612
rect 343220 165552 343270 165608
rect 343270 165552 343284 165608
rect 343220 165548 343284 165552
rect 343404 165608 343468 165612
rect 343404 165552 343454 165608
rect 343454 165552 343468 165608
rect 343404 165548 343468 165552
rect 398236 165548 398300 165612
rect 401732 165548 401796 165612
rect 405412 165548 405476 165612
rect 408172 165548 408236 165612
rect 410748 165548 410812 165612
rect 415900 165548 415964 165612
rect 416084 165608 416148 165612
rect 416084 165552 416098 165608
rect 416098 165552 416148 165608
rect 416084 165548 416148 165552
rect 419396 165548 419460 165612
rect 423812 165548 423876 165612
rect 426388 165548 426452 165612
rect 433380 165608 433444 165612
rect 433380 165552 433394 165608
rect 433394 165552 433444 165608
rect 433380 165548 433444 165552
rect 434300 165548 434364 165612
rect 435956 165548 436020 165612
rect 437796 165608 437860 165612
rect 437796 165552 437810 165608
rect 437810 165552 437860 165608
rect 437796 165548 437860 165552
rect 438532 165548 438596 165612
rect 443500 165548 443564 165612
rect 448284 165548 448348 165612
rect 451044 165548 451108 165612
rect 453436 165548 453500 165612
rect 455828 165548 455892 165612
rect 458404 165608 458468 165612
rect 458404 165552 458418 165608
rect 458418 165552 458468 165608
rect 458404 165548 458468 165552
rect 503300 165608 503364 165612
rect 503300 165552 503350 165608
rect 503350 165552 503364 165608
rect 503300 165548 503364 165552
rect 155908 165412 155972 165476
rect 213132 165412 213196 165476
rect 320956 165412 321020 165476
rect 468524 165412 468588 165476
rect 158484 165276 158548 165340
rect 206140 165276 206204 165340
rect 311020 165276 311084 165340
rect 465948 165276 466012 165340
rect 135852 165140 135916 165204
rect 213316 165140 213380 165204
rect 90772 165004 90836 165068
rect 113220 165064 113284 165068
rect 113220 165008 113234 165064
rect 113234 165008 113284 165064
rect 113220 165004 113284 165008
rect 216260 165004 216324 165068
rect 272196 165140 272260 165204
rect 275876 165200 275940 165204
rect 275876 165144 275926 165200
rect 275926 165144 275940 165200
rect 275876 165140 275940 165144
rect 276060 165140 276124 165204
rect 79548 164868 79612 164932
rect 88380 164928 88444 164932
rect 88380 164872 88394 164928
rect 88394 164872 88444 164928
rect 88380 164868 88444 164872
rect 93716 164868 93780 164932
rect 114508 164928 114572 164932
rect 114508 164872 114522 164928
rect 114522 164872 114572 164928
rect 114508 164868 114572 164872
rect 207980 164868 208044 164932
rect 263732 164868 263796 164932
rect 273484 165004 273548 165068
rect 278452 165140 278516 165204
rect 279188 165140 279252 165204
rect 374868 165140 374932 165204
rect 463556 165140 463620 165204
rect 379468 165004 379532 165068
rect 426020 165004 426084 165068
rect 433564 165004 433628 165068
rect 440924 164868 440988 164932
rect 160876 164732 160940 164796
rect 200804 164732 200868 164796
rect 256188 164732 256252 164796
rect 413692 164732 413756 164796
rect 421788 164732 421852 164796
rect 111196 164656 111260 164660
rect 111196 164600 111210 164656
rect 111210 164600 111260 164656
rect 111196 164596 111260 164600
rect 460980 164596 461044 164660
rect 115796 164460 115860 164524
rect 117084 164460 117148 164524
rect 244412 164460 244476 164524
rect 252324 164460 252388 164524
rect 260604 164460 260668 164524
rect 267596 164460 267660 164524
rect 273300 164460 273364 164524
rect 436876 164460 436940 164524
rect 77156 164324 77220 164388
rect 203012 164324 203076 164388
rect 315068 164324 315132 164388
rect 397132 164324 397196 164388
rect 404124 164324 404188 164388
rect 412404 164324 412468 164388
rect 429700 164324 429764 164388
rect 57284 164188 57348 164252
rect 76052 164188 76116 164252
rect 78260 164188 78324 164252
rect 80468 164188 80532 164252
rect 83044 164188 83108 164252
rect 84148 164248 84212 164252
rect 84148 164192 84198 164248
rect 84198 164192 84212 164248
rect 84148 164188 84212 164192
rect 86540 164188 86604 164252
rect 87644 164188 87708 164252
rect 88748 164188 88812 164252
rect 90036 164188 90100 164252
rect 91324 164188 91388 164252
rect 93348 164188 93412 164252
rect 94452 164188 94516 164252
rect 97028 164188 97092 164252
rect 98132 164188 98196 164252
rect 101812 164188 101876 164252
rect 102732 164188 102796 164252
rect 103836 164188 103900 164252
rect 237052 164188 237116 164252
rect 238156 164188 238220 164252
rect 240548 164188 240612 164252
rect 241652 164188 241716 164252
rect 245332 164188 245396 164252
rect 246436 164188 246500 164252
rect 248644 164188 248708 164252
rect 250116 164188 250180 164252
rect 251220 164248 251284 164252
rect 251220 164192 251234 164248
rect 251234 164192 251284 164248
rect 251220 164188 251284 164192
rect 253428 164188 253492 164252
rect 254532 164188 254596 164252
rect 255820 164188 255884 164252
rect 256924 164188 256988 164252
rect 258396 164188 258460 164252
rect 259500 164248 259564 164252
rect 259500 164192 259514 164248
rect 259514 164192 259564 164248
rect 259500 164188 259564 164192
rect 262812 164188 262876 164252
rect 263916 164188 263980 164252
rect 268700 164188 268764 164252
rect 269804 164188 269868 164252
rect 271276 164188 271340 164252
rect 274404 164188 274468 164252
rect 276980 164188 277044 164252
rect 278084 164188 278148 164252
rect 57652 164112 57716 164116
rect 57652 164056 57702 164112
rect 57702 164056 57716 164112
rect 57652 164052 57716 164056
rect 208164 164052 208228 164116
rect 318380 164188 318444 164252
rect 396028 164188 396092 164252
rect 399524 164188 399588 164252
rect 400444 164188 400508 164252
rect 403020 164248 403084 164252
rect 403020 164192 403070 164248
rect 403070 164192 403084 164248
rect 403020 164188 403084 164192
rect 406516 164188 406580 164252
rect 407620 164188 407684 164252
rect 408724 164188 408788 164252
rect 410012 164248 410076 164252
rect 410012 164192 410026 164248
rect 410026 164192 410076 164248
rect 410012 164188 410076 164192
rect 411300 164248 411364 164252
rect 411300 164192 411314 164248
rect 411314 164192 411364 164248
rect 411300 164188 411364 164192
rect 413324 164188 413388 164252
rect 414428 164188 414492 164252
rect 417004 164188 417068 164252
rect 418292 164188 418356 164252
rect 420684 164188 420748 164252
rect 422892 164188 422956 164252
rect 425284 164188 425348 164252
rect 427676 164248 427740 164252
rect 427676 164192 427726 164248
rect 427726 164192 427740 164248
rect 427676 164188 427740 164192
rect 428780 164188 428844 164252
rect 431172 164188 431236 164252
rect 432276 164188 432340 164252
rect 435772 164188 435836 164252
rect 439268 164188 439332 164252
rect 57836 163916 57900 163980
rect 377260 162964 377324 163028
rect 217548 162692 217612 162756
rect 360884 149092 360948 149156
rect 217364 146372 217428 146436
rect 377996 146236 378060 146300
rect 377628 146100 377692 146164
rect 510844 145420 510908 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 190868 144876 190932 144940
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144876 499868 144940
rect 377812 144060 377876 144124
rect 57284 140796 57348 140860
rect 57468 70348 57532 70412
rect 44956 67764 45020 67828
rect 216076 68036 216140 68100
rect 374684 68036 374748 68100
rect 218652 60616 218716 60620
rect 218652 60560 218702 60616
rect 218702 60560 218716 60616
rect 218652 60556 218716 60560
rect 219204 60616 219268 60620
rect 219204 60560 219254 60616
rect 219254 60560 219268 60616
rect 219204 60556 219268 60560
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 94550 59800 94614 59804
rect 94550 59744 94558 59800
rect 94558 59744 94614 59800
rect 94550 59740 94614 59744
rect 99446 59800 99510 59804
rect 99446 59744 99470 59800
rect 99470 59744 99510 59800
rect 99446 59740 99510 59744
rect 102846 59740 102910 59804
rect 105974 59740 106038 59804
rect 237142 59800 237206 59804
rect 237142 59744 237158 59800
rect 237158 59744 237206 59800
rect 237142 59740 237206 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 256998 59800 257062 59804
rect 256998 59744 257030 59800
rect 257030 59744 257062 59800
rect 256998 59740 257062 59744
rect 262846 59800 262910 59804
rect 262846 59744 262862 59800
rect 262862 59744 262910 59800
rect 262846 59740 262910 59744
rect 263934 59740 263998 59804
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 416046 59800 416110 59804
rect 416046 59744 416098 59800
rect 416098 59744 416110 59800
rect 416046 59740 416110 59744
rect 416998 59800 417062 59804
rect 416998 59744 417018 59800
rect 417018 59744 417062 59800
rect 416998 59740 417062 59744
rect 422846 59800 422910 59804
rect 422846 59744 422850 59800
rect 422850 59744 422906 59800
rect 422906 59744 422910 59800
rect 422846 59740 422910 59744
rect 423934 59800 423998 59804
rect 423934 59744 423954 59800
rect 423954 59744 423998 59800
rect 423934 59740 423998 59744
rect 57652 59468 57716 59532
rect 105294 59604 105358 59668
rect 107606 59664 107670 59668
rect 107606 59608 107622 59664
rect 107622 59608 107670 59664
rect 107606 59604 107670 59608
rect 258086 59664 258150 59668
rect 258086 59608 258134 59664
rect 258134 59608 258150 59664
rect 258086 59604 258150 59608
rect 260670 59664 260734 59668
rect 260670 59608 260710 59664
rect 260710 59608 260734 59664
rect 260670 59604 260734 59608
rect 261758 59664 261822 59668
rect 261758 59608 261814 59664
rect 261814 59608 261822 59664
rect 261758 59604 261822 59608
rect 308542 59664 308606 59668
rect 308542 59608 308550 59664
rect 308550 59608 308606 59664
rect 308542 59604 308606 59608
rect 315886 59664 315950 59668
rect 315886 59608 315910 59664
rect 315910 59608 315950 59664
rect 315886 59604 315950 59608
rect 403126 59604 403190 59668
rect 404214 59664 404278 59668
rect 404214 59608 404230 59664
rect 404230 59608 404278 59664
rect 404214 59604 404278 59608
rect 413462 59604 413526 59668
rect 423526 59664 423590 59668
rect 423526 59608 423550 59664
rect 423550 59608 423590 59664
rect 423526 59604 423590 59608
rect 90036 59528 90100 59532
rect 90036 59472 90050 59528
rect 90050 59472 90100 59528
rect 90036 59468 90100 59472
rect 95924 59528 95988 59532
rect 95924 59472 95938 59528
rect 95938 59472 95988 59528
rect 95924 59468 95988 59472
rect 97028 59528 97092 59532
rect 97028 59472 97042 59528
rect 97042 59472 97092 59528
rect 97028 59468 97092 59472
rect 100708 59528 100772 59532
rect 100708 59472 100758 59528
rect 100758 59472 100772 59528
rect 100708 59468 100772 59472
rect 101812 59528 101876 59532
rect 101812 59472 101826 59528
rect 101826 59472 101876 59528
rect 101812 59468 101876 59472
rect 48452 59332 48516 59396
rect 113588 59332 113652 59396
rect 200620 59332 200684 59396
rect 263548 59332 263612 59396
rect 418108 59392 418172 59396
rect 418108 59336 418158 59392
rect 418158 59336 418172 59392
rect 52316 59196 52380 59260
rect 143580 59196 143644 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 206692 59196 206756 59260
rect 279188 59256 279252 59260
rect 279188 59200 279238 59256
rect 279238 59200 279252 59256
rect 279188 59196 279252 59200
rect 418108 59332 418172 59336
rect 419396 59392 419460 59396
rect 419396 59336 419410 59392
rect 419410 59336 419460 59392
rect 419396 59332 419460 59336
rect 420684 59392 420748 59396
rect 420684 59336 420698 59392
rect 420698 59336 420748 59392
rect 420684 59332 420748 59336
rect 421788 59392 421852 59396
rect 421788 59336 421802 59392
rect 421802 59336 421852 59392
rect 421788 59332 421852 59336
rect 426020 59392 426084 59396
rect 426020 59336 426034 59392
rect 426034 59336 426084 59392
rect 426020 59332 426084 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 453436 59392 453500 59396
rect 453436 59336 453450 59392
rect 453450 59336 453500 59392
rect 453436 59332 453500 59336
rect 285996 59196 286060 59260
rect 290964 59256 291028 59260
rect 290964 59200 290978 59256
rect 290978 59200 291028 59256
rect 290964 59196 291028 59200
rect 300900 59256 300964 59260
rect 300900 59200 300914 59256
rect 300914 59200 300964 59256
rect 300900 59196 300964 59200
rect 320956 59256 321020 59260
rect 320956 59200 320970 59256
rect 320970 59200 321020 59256
rect 320956 59196 321020 59200
rect 325924 59256 325988 59260
rect 325924 59200 325938 59256
rect 325938 59200 325988 59256
rect 325924 59196 325988 59200
rect 360700 59196 360764 59260
rect 483428 59196 483492 59260
rect 54892 59060 54956 59124
rect 140820 59060 140884 59124
rect 209636 59060 209700 59124
rect 280844 59060 280908 59124
rect 371924 59060 371988 59124
rect 480852 59060 480916 59124
rect 52132 58924 52196 58988
rect 135852 58924 135916 58988
rect 138428 58984 138492 58988
rect 138428 58928 138442 58984
rect 138442 58928 138492 58984
rect 138428 58924 138492 58928
rect 198044 58924 198108 58988
rect 268332 58924 268396 58988
rect 366220 58924 366284 58988
rect 468524 58924 468588 58988
rect 475884 58984 475948 58988
rect 475884 58928 475898 58984
rect 475898 58928 475948 58984
rect 475884 58924 475948 58928
rect 48636 58788 48700 58852
rect 111012 58788 111076 58852
rect 206876 58788 206940 58852
rect 276060 58788 276124 58852
rect 373764 58788 373828 58852
rect 473492 58788 473556 58852
rect 59308 58652 59372 58716
rect 120948 58652 121012 58716
rect 197860 58652 197924 58716
rect 253612 58652 253676 58716
rect 371740 58652 371804 58716
rect 463556 58652 463620 58716
rect 47900 58516 47964 58580
rect 108252 58516 108316 58580
rect 202276 58516 202340 58580
rect 250668 58516 250732 58580
rect 370452 58516 370516 58580
rect 458404 58516 458468 58580
rect 59124 58380 59188 58444
rect 101076 58380 101140 58444
rect 217548 58380 217612 58444
rect 259500 58380 259564 58444
rect 376156 58380 376220 58444
rect 410748 58380 410812 58444
rect 85436 58108 85500 58172
rect 92428 58108 92492 58172
rect 128308 58108 128372 58172
rect 153332 58108 153396 58172
rect 235948 58108 236012 58172
rect 265204 58108 265268 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 398236 58108 398300 58172
rect 401732 58108 401796 58172
rect 405412 58108 405476 58172
rect 83964 57972 84028 58036
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57836 79612 57900
rect 80468 57896 80532 57900
rect 80468 57840 80482 57896
rect 80482 57840 80532 57896
rect 80468 57836 80532 57840
rect 81940 57836 82004 57900
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88380 57896 88444 57900
rect 88380 57840 88394 57896
rect 88394 57840 88444 57896
rect 88380 57836 88444 57840
rect 88748 57896 88812 57900
rect 88748 57840 88762 57896
rect 88762 57840 88812 57896
rect 88748 57836 88812 57840
rect 90772 57836 90836 57900
rect 91324 57836 91388 57900
rect 93348 57896 93412 57900
rect 93348 57840 93362 57896
rect 93362 57840 93412 57896
rect 93348 57836 93412 57840
rect 93716 57896 93780 57900
rect 93716 57840 93730 57896
rect 93730 57840 93780 57896
rect 93716 57836 93780 57840
rect 98132 57896 98196 57900
rect 98132 57840 98146 57896
rect 98146 57840 98196 57896
rect 98132 57836 98196 57840
rect 103836 57896 103900 57900
rect 103836 57840 103850 57896
rect 103850 57840 103900 57896
rect 103836 57836 103900 57840
rect 108620 57896 108684 57900
rect 108620 57840 108634 57896
rect 108634 57840 108684 57896
rect 108620 57836 108684 57840
rect 109540 57896 109604 57900
rect 109540 57840 109554 57896
rect 109554 57840 109604 57896
rect 109540 57836 109604 57840
rect 112116 57896 112180 57900
rect 112116 57840 112130 57896
rect 112130 57840 112180 57896
rect 112116 57836 112180 57840
rect 113220 57896 113284 57900
rect 113220 57840 113234 57896
rect 113234 57840 113284 57896
rect 113220 57836 113284 57840
rect 114324 57836 114388 57900
rect 115980 57896 116044 57900
rect 115980 57840 115994 57896
rect 115994 57840 116044 57896
rect 115980 57836 116044 57840
rect 118004 57836 118068 57900
rect 119108 57896 119172 57900
rect 119108 57840 119122 57896
rect 119122 57840 119172 57896
rect 119108 57836 119172 57840
rect 123524 57896 123588 57900
rect 123524 57840 123538 57896
rect 123538 57840 123588 57896
rect 123524 57836 123588 57840
rect 55076 57700 55140 57764
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 183508 57896 183572 57900
rect 183508 57840 183522 57896
rect 183522 57840 183572 57896
rect 183508 57836 183572 57840
rect 238156 57836 238220 57900
rect 239260 57836 239324 57900
rect 240548 57836 240612 57900
rect 241652 57896 241716 57900
rect 241652 57840 241666 57896
rect 241666 57840 241716 57896
rect 241652 57836 241716 57840
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 244228 57836 244292 57900
rect 245332 57896 245396 57900
rect 245332 57840 245346 57896
rect 245346 57840 245396 57896
rect 245332 57836 245396 57840
rect 246436 57836 246500 57900
rect 247724 57836 247788 57900
rect 248644 57896 248708 57900
rect 248644 57840 248658 57896
rect 248658 57840 248708 57896
rect 248644 57836 248708 57840
rect 250116 57836 250180 57900
rect 251220 57896 251284 57900
rect 251220 57840 251234 57896
rect 251234 57840 251284 57896
rect 251220 57836 251284 57840
rect 252324 57836 252388 57900
rect 253428 57896 253492 57900
rect 253428 57840 253442 57896
rect 253442 57840 253492 57896
rect 253428 57836 253492 57840
rect 254532 57836 254596 57900
rect 258396 57896 258460 57900
rect 258396 57840 258410 57896
rect 258410 57840 258460 57896
rect 258396 57836 258460 57840
rect 266308 57896 266372 57900
rect 266308 57840 266358 57896
rect 266358 57840 266372 57896
rect 266308 57836 266372 57840
rect 268700 57836 268764 57900
rect 271092 57896 271156 57900
rect 271092 57840 271106 57896
rect 271106 57840 271156 57896
rect 271092 57836 271156 57840
rect 273300 57896 273364 57900
rect 273300 57840 273314 57896
rect 273314 57840 273364 57896
rect 273300 57836 273364 57840
rect 283788 57836 283852 57900
rect 293356 57896 293420 57900
rect 293356 57840 293370 57896
rect 293370 57840 293420 57896
rect 293356 57836 293420 57840
rect 295932 57896 295996 57900
rect 295932 57840 295946 57896
rect 295946 57840 295996 57896
rect 295932 57836 295996 57840
rect 298508 57836 298572 57900
rect 303476 57896 303540 57900
rect 303476 57840 303490 57896
rect 303490 57840 303540 57896
rect 303476 57836 303540 57840
rect 305868 57896 305932 57900
rect 305868 57840 305882 57896
rect 305882 57840 305932 57896
rect 305868 57836 305932 57840
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 313412 57896 313476 57900
rect 313412 57840 313426 57896
rect 313426 57840 313476 57896
rect 313412 57836 313476 57840
rect 318380 57896 318444 57900
rect 318380 57840 318394 57896
rect 318394 57840 318444 57896
rect 318380 57836 318444 57840
rect 323348 57896 323412 57900
rect 323348 57840 323362 57896
rect 323362 57840 323412 57896
rect 323348 57836 323412 57840
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57836 399588 57900
rect 400444 57896 400508 57900
rect 400444 57840 400458 57896
rect 400458 57840 400508 57896
rect 400444 57836 400508 57840
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 414612 57896 414676 57900
rect 414612 57840 414626 57896
rect 414626 57840 414676 57896
rect 414612 57836 414676 57840
rect 415532 57896 415596 57900
rect 415532 57840 415546 57896
rect 415546 57840 415596 57896
rect 415532 57836 415596 57840
rect 418476 57896 418540 57900
rect 418476 57840 418490 57896
rect 418490 57840 418540 57896
rect 418476 57836 418540 57840
rect 425284 57836 425348 57900
rect 426388 57896 426452 57900
rect 426388 57840 426438 57896
rect 426438 57840 426452 57896
rect 426388 57836 426452 57840
rect 427676 57896 427740 57900
rect 427676 57840 427690 57896
rect 427690 57840 427740 57896
rect 427676 57836 427740 57840
rect 428596 57836 428660 57900
rect 429700 57836 429764 57900
rect 431172 57896 431236 57900
rect 431172 57840 431186 57896
rect 431186 57840 431236 57896
rect 431172 57836 431236 57840
rect 432276 57836 432340 57900
rect 433380 57896 433444 57900
rect 433380 57840 433394 57896
rect 433394 57840 433444 57896
rect 433380 57836 433444 57840
rect 433564 57896 433628 57900
rect 433564 57840 433578 57896
rect 433578 57840 433628 57896
rect 433564 57836 433628 57840
rect 435772 57896 435836 57900
rect 435772 57840 435786 57896
rect 435786 57840 435836 57896
rect 435772 57836 435836 57840
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 443500 57896 443564 57900
rect 443500 57840 443514 57896
rect 443514 57840 443564 57896
rect 443500 57836 443564 57840
rect 445892 57896 445956 57900
rect 445892 57840 445906 57896
rect 445906 57840 445956 57896
rect 445892 57836 445956 57840
rect 448284 57896 448348 57900
rect 448284 57840 448298 57896
rect 448298 57840 448348 57896
rect 448284 57836 448348 57840
rect 465948 57896 466012 57900
rect 465948 57840 465962 57896
rect 465962 57840 466012 57896
rect 465948 57836 466012 57840
rect 478460 57896 478524 57900
rect 478460 57840 478474 57896
rect 478474 57840 478524 57896
rect 478460 57836 478524 57840
rect 486004 57896 486068 57900
rect 486004 57840 486018 57896
rect 486018 57840 486068 57896
rect 486004 57836 486068 57840
rect 503116 57836 503180 57900
rect 503484 57896 503548 57900
rect 503484 57840 503534 57896
rect 503534 57840 503548 57896
rect 503484 57836 503548 57840
rect 183140 57760 183204 57764
rect 183140 57704 183190 57760
rect 183190 57704 183204 57760
rect 183140 57700 183204 57704
rect 210740 57700 210804 57764
rect 278452 57700 278516 57764
rect 378732 57700 378796 57764
rect 470916 57700 470980 57764
rect 60228 57564 60292 57628
rect 125916 57564 125980 57628
rect 158484 57564 158548 57628
rect 160876 57564 160940 57628
rect 165844 57564 165908 57628
rect 208900 57564 208964 57628
rect 54708 57428 54772 57492
rect 58572 57292 58636 57356
rect 103836 57292 103900 57356
rect 106412 57428 106476 57492
rect 111196 57428 111260 57492
rect 115796 57428 115860 57492
rect 116900 57428 116964 57492
rect 203196 57428 203260 57492
rect 260972 57428 261036 57492
rect 267596 57564 267660 57628
rect 269804 57564 269868 57628
rect 274404 57564 274468 57628
rect 278084 57564 278148 57628
rect 357940 57564 358004 57628
rect 434668 57564 434732 57628
rect 436876 57564 436940 57628
rect 439084 57564 439148 57628
rect 270908 57428 270972 57492
rect 379100 57428 379164 57492
rect 456380 57428 456444 57492
rect 118372 57292 118436 57356
rect 205036 57292 205100 57356
rect 256004 57292 256068 57356
rect 374500 57292 374564 57356
rect 451044 57292 451108 57356
rect 58756 57156 58820 57220
rect 98500 57156 98564 57220
rect 215892 57156 215956 57220
rect 265940 57156 266004 57220
rect 379284 57156 379348 57220
rect 430988 57156 431052 57220
rect 440924 57156 440988 57220
rect 58940 57020 59004 57084
rect 96292 57020 96356 57084
rect 214420 57020 214484 57084
rect 248276 57020 248340 57084
rect 378916 57020 378980 57084
rect 413508 57020 413572 57084
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 55444 56612 55508 56676
rect 133460 56612 133524 56676
rect 163268 56612 163332 56676
rect 214604 56612 214668 56676
rect 288204 56612 288268 56676
rect 367692 56612 367756 56676
rect 460980 56612 461044 56676
rect 50660 56476 50724 56540
rect 219940 56476 220004 56540
rect 421052 56476 421116 56540
rect 50476 56340 50540 56404
rect 201356 56340 201420 56404
rect 273484 56340 273548 56404
rect 377260 56340 377324 56404
rect 438348 56340 438412 56404
rect 55628 56204 55692 56268
rect 155908 56204 155972 56268
rect 217364 56204 217428 56268
rect 276980 56204 277044 56268
rect 57284 56068 57348 56132
rect 48084 55116 48148 55180
rect 377812 55116 377876 55180
rect 50844 54980 50908 55044
rect 377628 54980 377692 55044
rect 53604 54844 53668 54908
rect 57836 54708 57900 54772
rect 210372 3980 210436 4044
rect 202092 3844 202156 3908
rect 364932 3708 364996 3772
rect 363460 3572 363524 3636
rect 375972 3436 376036 3500
rect 365116 3300 365180 3364
rect 204852 3164 204916 3228
rect 368244 2892 368308 2956
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 44955 485348 45021 485349
rect 44955 485284 44956 485348
rect 45020 485284 45021 485348
rect 44955 485283 45021 485284
rect 44771 476780 44837 476781
rect 44771 476716 44772 476780
rect 44836 476716 44837 476780
rect 44771 476715 44837 476716
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 44774 268429 44834 476715
rect 44771 268428 44837 268429
rect 44771 268364 44772 268428
rect 44836 268364 44837 268428
rect 44771 268363 44837 268364
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 44958 67829 45018 485283
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 53051 639300 53117 639301
rect 53051 639236 53052 639300
rect 53116 639236 53117 639300
rect 53051 639235 53117 639236
rect 51579 639164 51645 639165
rect 51579 639100 51580 639164
rect 51644 639100 51645 639164
rect 51579 639099 51645 639100
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 46611 482356 46677 482357
rect 46611 482292 46612 482356
rect 46676 482292 46677 482356
rect 46611 482291 46677 482292
rect 48954 482294 49574 482378
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 46614 267749 46674 482291
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 46795 476916 46861 476917
rect 46795 476852 46796 476916
rect 46860 476852 46861 476916
rect 46795 476851 46861 476852
rect 46611 267748 46677 267749
rect 46611 267684 46612 267748
rect 46676 267684 46677 267748
rect 46611 267683 46677 267684
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 46798 251157 46858 476851
rect 47899 469164 47965 469165
rect 47899 469100 47900 469164
rect 47964 469100 47965 469164
rect 47899 469099 47965 469100
rect 46795 251156 46861 251157
rect 46795 251092 46796 251156
rect 46860 251092 46861 251156
rect 46795 251091 46861 251092
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 44955 67828 45021 67829
rect 44955 67764 44956 67828
rect 45020 67764 45021 67828
rect 44955 67763 45021 67764
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 46894 45854 82338
rect 47902 58581 47962 469099
rect 48635 469028 48701 469029
rect 48635 468964 48636 469028
rect 48700 468964 48701 469028
rect 48635 468963 48701 468964
rect 48083 467940 48149 467941
rect 48083 467876 48084 467940
rect 48148 467876 48149 467940
rect 48083 467875 48149 467876
rect 47899 58580 47965 58581
rect 47899 58516 47900 58580
rect 47964 58516 47965 58580
rect 47899 58515 47965 58516
rect 48086 55181 48146 467875
rect 48451 466172 48517 466173
rect 48451 466108 48452 466172
rect 48516 466108 48517 466172
rect 48451 466107 48517 466108
rect 48454 59397 48514 466107
rect 48451 59396 48517 59397
rect 48451 59332 48452 59396
rect 48516 59332 48517 59396
rect 48451 59331 48517 59332
rect 48638 58853 48698 468963
rect 48954 446614 49574 482058
rect 50475 468620 50541 468621
rect 50475 468556 50476 468620
rect 50540 468556 50541 468620
rect 50475 468555 50541 468556
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48635 58852 48701 58853
rect 48635 58788 48636 58852
rect 48700 58788 48701 58852
rect 48635 58787 48701 58788
rect 48083 55180 48149 55181
rect 48083 55116 48084 55180
rect 48148 55116 48149 55180
rect 48083 55115 48149 55116
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50478 56405 50538 468555
rect 50843 468484 50909 468485
rect 50843 468420 50844 468484
rect 50908 468420 50909 468484
rect 50843 468419 50909 468420
rect 50659 467940 50725 467941
rect 50659 467876 50660 467940
rect 50724 467876 50725 467940
rect 50659 467875 50725 467876
rect 50662 56541 50722 467875
rect 50659 56540 50725 56541
rect 50659 56476 50660 56540
rect 50724 56476 50725 56540
rect 50659 56475 50725 56476
rect 50475 56404 50541 56405
rect 50475 56340 50476 56404
rect 50540 56340 50541 56404
rect 50475 56339 50541 56340
rect 50846 55045 50906 468419
rect 51582 201517 51642 639099
rect 52131 465900 52197 465901
rect 52131 465836 52132 465900
rect 52196 465836 52197 465900
rect 52131 465835 52197 465836
rect 51763 465220 51829 465221
rect 51763 465156 51764 465220
rect 51828 465156 51829 465220
rect 51763 465155 51829 465156
rect 51766 379541 51826 465155
rect 51763 379540 51829 379541
rect 51763 379476 51764 379540
rect 51828 379476 51829 379540
rect 51763 379475 51829 379476
rect 51579 201516 51645 201517
rect 51579 201452 51580 201516
rect 51644 201452 51645 201516
rect 51579 201451 51645 201452
rect 52134 58989 52194 465835
rect 52315 465764 52381 465765
rect 52315 465700 52316 465764
rect 52380 465700 52381 465764
rect 52315 465699 52381 465700
rect 52318 59261 52378 465699
rect 53054 254013 53114 639235
rect 54339 639028 54405 639029
rect 54339 638964 54340 639028
rect 54404 638964 54405 639028
rect 54339 638963 54405 638964
rect 53603 468756 53669 468757
rect 53603 468692 53604 468756
rect 53668 468692 53669 468756
rect 53603 468691 53669 468692
rect 53235 466036 53301 466037
rect 53235 465972 53236 466036
rect 53300 465972 53301 466036
rect 53235 465971 53301 465972
rect 53238 378861 53298 465971
rect 53235 378860 53301 378861
rect 53235 378796 53236 378860
rect 53300 378796 53301 378860
rect 53235 378795 53301 378796
rect 53051 254012 53117 254013
rect 53051 253948 53052 254012
rect 53116 253948 53117 254012
rect 53051 253947 53117 253948
rect 52315 59260 52381 59261
rect 52315 59196 52316 59260
rect 52380 59196 52381 59260
rect 52315 59195 52381 59196
rect 52131 58988 52197 58989
rect 52131 58924 52132 58988
rect 52196 58924 52197 58988
rect 52131 58923 52197 58924
rect 50843 55044 50909 55045
rect 50843 54980 50844 55044
rect 50908 54980 50909 55044
rect 50843 54979 50909 54980
rect 53606 54909 53666 468691
rect 54342 305013 54402 638963
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 633099 60134 636618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 633099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 633099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 633099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 633099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 633099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 633099 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633099 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 633099 96134 636618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 633099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 633099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 633099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 633099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 633099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 633099 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 55794 597454 56414 632898
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 565174 60134 566000
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 550000 60134 564618
rect 63234 551834 63854 566000
rect 63234 551598 63266 551834
rect 63502 551598 63586 551834
rect 63822 551598 63854 551834
rect 63234 551514 63854 551598
rect 63234 551278 63266 551514
rect 63502 551278 63586 551514
rect 63822 551278 63854 551514
rect 63234 550000 63854 551278
rect 66954 555554 67574 566000
rect 66954 555318 66986 555554
rect 67222 555318 67306 555554
rect 67542 555318 67574 555554
rect 66954 555234 67574 555318
rect 66954 554998 66986 555234
rect 67222 554998 67306 555234
rect 67542 554998 67574 555234
rect 66954 550000 67574 554998
rect 73794 560514 74414 566000
rect 73794 560278 73826 560514
rect 74062 560278 74146 560514
rect 74382 560278 74414 560514
rect 73794 560194 74414 560278
rect 73794 559958 73826 560194
rect 74062 559958 74146 560194
rect 74382 559958 74414 560194
rect 73794 550000 74414 559958
rect 77514 564234 78134 566000
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 78134 564234
rect 77514 563914 78134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 78134 563914
rect 77514 550000 78134 563678
rect 81234 550894 81854 566000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 550000 81854 550338
rect 84954 554614 85574 566000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 550000 85574 554058
rect 91794 561454 92414 566000
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 550000 92414 560898
rect 95514 565174 96134 566000
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 550000 96134 564618
rect 99234 551834 99854 566000
rect 99234 551598 99266 551834
rect 99502 551598 99586 551834
rect 99822 551598 99854 551834
rect 99234 551514 99854 551598
rect 99234 551278 99266 551514
rect 99502 551278 99586 551514
rect 99822 551278 99854 551514
rect 99234 550000 99854 551278
rect 102954 555554 103574 566000
rect 102954 555318 102986 555554
rect 103222 555318 103306 555554
rect 103542 555318 103574 555554
rect 102954 555234 103574 555318
rect 102954 554998 102986 555234
rect 103222 554998 103306 555234
rect 103542 554998 103574 555234
rect 102954 550000 103574 554998
rect 109794 560514 110414 566000
rect 109794 560278 109826 560514
rect 110062 560278 110146 560514
rect 110382 560278 110414 560514
rect 109794 560194 110414 560278
rect 109794 559958 109826 560194
rect 110062 559958 110146 560194
rect 110382 559958 110414 560194
rect 109794 550000 110414 559958
rect 113514 564234 114134 566000
rect 113514 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 114134 564234
rect 113514 563914 114134 563998
rect 113514 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 114134 563914
rect 113514 550000 114134 563678
rect 117234 550894 117854 566000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 550000 117854 550338
rect 120954 554614 121574 566000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 550000 121574 554058
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 550000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 550000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 633099 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 633099 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 633099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 633099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 633099 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633099 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 633099 168134 636618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 633099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 633099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 633099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 633099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 633099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 633099 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633099 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 144208 615454 144528 615486
rect 144208 615218 144250 615454
rect 144486 615218 144528 615454
rect 144208 615134 144528 615218
rect 144208 614898 144250 615134
rect 144486 614898 144528 615134
rect 144208 614866 144528 614898
rect 174928 615454 175248 615486
rect 174928 615218 174970 615454
rect 175206 615218 175248 615454
rect 174928 615134 175248 615218
rect 174928 614898 174970 615134
rect 175206 614898 175248 615134
rect 174928 614866 175248 614898
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 159568 597454 159888 597486
rect 159568 597218 159610 597454
rect 159846 597218 159888 597454
rect 159568 597134 159888 597218
rect 159568 596898 159610 597134
rect 159846 596898 159888 597134
rect 159568 596866 159888 596898
rect 190288 597454 190608 597486
rect 190288 597218 190330 597454
rect 190566 597218 190608 597454
rect 190288 597134 190608 597218
rect 190288 596898 190330 597134
rect 190566 596898 190608 597134
rect 190288 596866 190608 596898
rect 144208 579454 144528 579486
rect 144208 579218 144250 579454
rect 144486 579218 144528 579454
rect 144208 579134 144528 579218
rect 144208 578898 144250 579134
rect 144486 578898 144528 579134
rect 144208 578866 144528 578898
rect 174928 579454 175248 579486
rect 174928 579218 174970 579454
rect 175206 579218 175248 579454
rect 174928 579134 175248 579218
rect 174928 578898 174970 579134
rect 175206 578898 175248 579134
rect 174928 578866 175248 578898
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 551834 135854 568338
rect 135234 551598 135266 551834
rect 135502 551598 135586 551834
rect 135822 551598 135854 551834
rect 135234 551514 135854 551598
rect 135234 551278 135266 551514
rect 135502 551278 135586 551514
rect 135822 551278 135854 551514
rect 135234 550000 135854 551278
rect 138954 555554 139574 566000
rect 138954 555318 138986 555554
rect 139222 555318 139306 555554
rect 139542 555318 139574 555554
rect 138954 555234 139574 555318
rect 138954 554998 138986 555234
rect 139222 554998 139306 555234
rect 139542 554998 139574 555234
rect 138954 550000 139574 554998
rect 145794 560514 146414 566000
rect 145794 560278 145826 560514
rect 146062 560278 146146 560514
rect 146382 560278 146414 560514
rect 145794 560194 146414 560278
rect 145794 559958 145826 560194
rect 146062 559958 146146 560194
rect 146382 559958 146414 560194
rect 145794 550000 146414 559958
rect 149514 564234 150134 566000
rect 149514 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 150134 564234
rect 149514 563914 150134 563998
rect 149514 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 150134 563914
rect 149514 550000 150134 563678
rect 153234 550894 153854 566000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 550000 153854 550338
rect 156954 554614 157574 566000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 550000 157574 554058
rect 163794 561454 164414 566000
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 550000 164414 560898
rect 167514 565174 168134 566000
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 550000 168134 564618
rect 171234 551834 171854 566000
rect 171234 551598 171266 551834
rect 171502 551598 171586 551834
rect 171822 551598 171854 551834
rect 171234 551514 171854 551598
rect 171234 551278 171266 551514
rect 171502 551278 171586 551514
rect 171822 551278 171854 551514
rect 171234 550000 171854 551278
rect 174954 555554 175574 566000
rect 174954 555318 174986 555554
rect 175222 555318 175306 555554
rect 175542 555318 175574 555554
rect 174954 555234 175574 555318
rect 174954 554998 174986 555234
rect 175222 554998 175306 555234
rect 175542 554998 175574 555234
rect 174954 550000 175574 554998
rect 181794 560514 182414 566000
rect 181794 560278 181826 560514
rect 182062 560278 182146 560514
rect 182382 560278 182414 560514
rect 181794 560194 182414 560278
rect 181794 559958 181826 560194
rect 182062 559958 182146 560194
rect 182382 559958 182414 560194
rect 181794 550000 182414 559958
rect 185514 564234 186134 566000
rect 185514 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 186134 564234
rect 185514 563914 186134 563998
rect 185514 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 186134 563914
rect 185514 550000 186134 563678
rect 189234 550894 189854 566000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 550000 189854 550338
rect 192954 554614 193574 566000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 550000 193574 554058
rect 199794 561454 200414 566000
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 550000 200414 560898
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 550000 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 551834 207854 568338
rect 207234 551598 207266 551834
rect 207502 551598 207586 551834
rect 207822 551598 207854 551834
rect 207234 551514 207854 551598
rect 207234 551278 207266 551514
rect 207502 551278 207586 551514
rect 207822 551278 207854 551514
rect 207234 550000 207854 551278
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 633099 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 633099 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 633099 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 633099 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633099 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 633099 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 633099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 633099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 633099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 633099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 633099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 633099 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633099 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 633099 276134 636618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 633099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 633099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 224208 615454 224528 615486
rect 224208 615218 224250 615454
rect 224486 615218 224528 615454
rect 224208 615134 224528 615218
rect 224208 614898 224250 615134
rect 224486 614898 224528 615134
rect 224208 614866 224528 614898
rect 254928 615454 255248 615486
rect 254928 615218 254970 615454
rect 255206 615218 255248 615454
rect 254928 615134 255248 615218
rect 254928 614898 254970 615134
rect 255206 614898 255248 615134
rect 254928 614866 255248 614898
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 239568 597454 239888 597486
rect 239568 597218 239610 597454
rect 239846 597218 239888 597454
rect 239568 597134 239888 597218
rect 239568 596898 239610 597134
rect 239846 596898 239888 597134
rect 239568 596866 239888 596898
rect 270288 597454 270608 597486
rect 270288 597218 270330 597454
rect 270566 597218 270608 597454
rect 270288 597134 270608 597218
rect 270288 596898 270330 597134
rect 270566 596898 270608 597134
rect 270288 596866 270608 596898
rect 224208 579454 224528 579486
rect 224208 579218 224250 579454
rect 224486 579218 224528 579454
rect 224208 579134 224528 579218
rect 224208 578898 224250 579134
rect 224486 578898 224528 579134
rect 224208 578866 224528 578898
rect 254928 579454 255248 579486
rect 254928 579218 254970 579454
rect 255206 579218 255248 579454
rect 254928 579134 255248 579218
rect 254928 578898 254970 579134
rect 255206 578898 255248 579134
rect 254928 578866 255248 578898
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 555554 211574 572058
rect 210954 555318 210986 555554
rect 211222 555318 211306 555554
rect 211542 555318 211574 555554
rect 210954 555234 211574 555318
rect 210954 554998 210986 555234
rect 211222 554998 211306 555234
rect 211542 554998 211574 555234
rect 210954 550000 211574 554998
rect 217794 560514 218414 566000
rect 217794 560278 217826 560514
rect 218062 560278 218146 560514
rect 218382 560278 218414 560514
rect 217794 560194 218414 560278
rect 217794 559958 217826 560194
rect 218062 559958 218146 560194
rect 218382 559958 218414 560194
rect 217794 550000 218414 559958
rect 221514 564234 222134 566000
rect 221514 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 222134 564234
rect 221514 563914 222134 563998
rect 221514 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 222134 563914
rect 221514 550000 222134 563678
rect 225234 550894 225854 566000
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 550000 225854 550338
rect 228954 554614 229574 566000
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 550000 229574 554058
rect 235794 561454 236414 566000
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 550000 236414 560898
rect 239514 565174 240134 566000
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 550000 240134 564618
rect 243234 551834 243854 566000
rect 243234 551598 243266 551834
rect 243502 551598 243586 551834
rect 243822 551598 243854 551834
rect 243234 551514 243854 551598
rect 243234 551278 243266 551514
rect 243502 551278 243586 551514
rect 243822 551278 243854 551514
rect 243234 550000 243854 551278
rect 246954 555554 247574 566000
rect 246954 555318 246986 555554
rect 247222 555318 247306 555554
rect 247542 555318 247574 555554
rect 246954 555234 247574 555318
rect 246954 554998 246986 555234
rect 247222 554998 247306 555234
rect 247542 554998 247574 555234
rect 246954 550000 247574 554998
rect 253794 560514 254414 566000
rect 253794 560278 253826 560514
rect 254062 560278 254146 560514
rect 254382 560278 254414 560514
rect 253794 560194 254414 560278
rect 253794 559958 253826 560194
rect 254062 559958 254146 560194
rect 254382 559958 254414 560194
rect 253794 550000 254414 559958
rect 257514 564234 258134 566000
rect 257514 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 258134 564234
rect 257514 563914 258134 563998
rect 257514 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 258134 563914
rect 257514 550000 258134 563678
rect 261234 550894 261854 566000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 550000 261854 550338
rect 264954 554614 265574 566000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 550000 265574 554058
rect 271794 561454 272414 566000
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 550000 272414 560898
rect 275514 565174 276134 566000
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 550000 276134 564618
rect 279234 551834 279854 566000
rect 279234 551598 279266 551834
rect 279502 551598 279586 551834
rect 279822 551598 279854 551834
rect 279234 551514 279854 551598
rect 279234 551278 279266 551514
rect 279502 551278 279586 551514
rect 279822 551278 279854 551514
rect 279234 550000 279854 551278
rect 282954 555554 283574 566000
rect 282954 555318 282986 555554
rect 283222 555318 283306 555554
rect 283542 555318 283574 555554
rect 282954 555234 283574 555318
rect 282954 554998 282986 555234
rect 283222 554998 283306 555234
rect 283542 554998 283574 555234
rect 282954 550000 283574 554998
rect 289794 550000 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 550000 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 550000 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 550000 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 64208 543454 64528 543486
rect 64208 543218 64250 543454
rect 64486 543218 64528 543454
rect 64208 543134 64528 543218
rect 64208 542898 64250 543134
rect 64486 542898 64528 543134
rect 64208 542866 64528 542898
rect 94928 543454 95248 543486
rect 94928 543218 94970 543454
rect 95206 543218 95248 543454
rect 94928 543134 95248 543218
rect 94928 542898 94970 543134
rect 95206 542898 95248 543134
rect 94928 542866 95248 542898
rect 125648 543454 125968 543486
rect 125648 543218 125690 543454
rect 125926 543218 125968 543454
rect 125648 543134 125968 543218
rect 125648 542898 125690 543134
rect 125926 542898 125968 543134
rect 125648 542866 125968 542898
rect 156368 543454 156688 543486
rect 156368 543218 156410 543454
rect 156646 543218 156688 543454
rect 156368 543134 156688 543218
rect 156368 542898 156410 543134
rect 156646 542898 156688 543134
rect 156368 542866 156688 542898
rect 187088 543454 187408 543486
rect 187088 543218 187130 543454
rect 187366 543218 187408 543454
rect 187088 543134 187408 543218
rect 187088 542898 187130 543134
rect 187366 542898 187408 543134
rect 187088 542866 187408 542898
rect 217808 543454 218128 543486
rect 217808 543218 217850 543454
rect 218086 543218 218128 543454
rect 217808 543134 218128 543218
rect 217808 542898 217850 543134
rect 218086 542898 218128 543134
rect 217808 542866 218128 542898
rect 248528 543454 248848 543486
rect 248528 543218 248570 543454
rect 248806 543218 248848 543454
rect 248528 543134 248848 543218
rect 248528 542898 248570 543134
rect 248806 542898 248848 543134
rect 248528 542866 248848 542898
rect 279248 543454 279568 543486
rect 279248 543218 279290 543454
rect 279526 543218 279568 543454
rect 279248 543134 279568 543218
rect 279248 542898 279290 543134
rect 279526 542898 279568 543134
rect 279248 542866 279568 542898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55075 485620 55141 485621
rect 55075 485556 55076 485620
rect 55140 485556 55141 485620
rect 55075 485555 55141 485556
rect 54891 485484 54957 485485
rect 54891 485420 54892 485484
rect 54956 485420 54957 485484
rect 54891 485419 54957 485420
rect 54707 466444 54773 466445
rect 54707 466380 54708 466444
rect 54772 466380 54773 466444
rect 54707 466379 54773 466380
rect 54339 305012 54405 305013
rect 54339 304948 54340 305012
rect 54404 304948 54405 305012
rect 54339 304947 54405 304948
rect 54710 57493 54770 466379
rect 54894 59125 54954 485419
rect 54891 59124 54957 59125
rect 54891 59060 54892 59124
rect 54956 59060 54957 59124
rect 54891 59059 54957 59060
rect 55078 57765 55138 485555
rect 55627 468892 55693 468893
rect 55627 468828 55628 468892
rect 55692 468828 55693 468892
rect 55627 468827 55693 468828
rect 55443 466172 55509 466173
rect 55443 466108 55444 466172
rect 55508 466108 55509 466172
rect 55443 466107 55509 466108
rect 55075 57764 55141 57765
rect 55075 57700 55076 57764
rect 55140 57700 55141 57764
rect 55075 57699 55141 57700
rect 54707 57492 54773 57493
rect 54707 57428 54708 57492
rect 54772 57428 54773 57492
rect 54707 57427 54773 57428
rect 55446 56677 55506 466107
rect 55443 56676 55509 56677
rect 55443 56612 55444 56676
rect 55508 56612 55509 56676
rect 55443 56611 55509 56612
rect 55630 56269 55690 468827
rect 55794 453454 56414 488898
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 57835 485212 57901 485213
rect 57835 485148 57836 485212
rect 57900 485148 57901 485212
rect 57835 485147 57901 485148
rect 57099 482764 57165 482765
rect 57099 482700 57100 482764
rect 57164 482700 57165 482764
rect 57099 482699 57165 482700
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57102 378997 57162 482699
rect 57467 479772 57533 479773
rect 57467 479708 57468 479772
rect 57532 479708 57533 479772
rect 57467 479707 57533 479708
rect 57099 378996 57165 378997
rect 57099 378932 57100 378996
rect 57164 378932 57165 378996
rect 57099 378931 57165 378932
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57470 270333 57530 479707
rect 57651 466308 57717 466309
rect 57651 466244 57652 466308
rect 57716 466244 57717 466308
rect 57651 466243 57717 466244
rect 57654 388653 57714 466243
rect 57651 388652 57717 388653
rect 57651 388588 57652 388652
rect 57716 388588 57717 388652
rect 57651 388587 57717 388588
rect 57651 388516 57717 388517
rect 57651 388452 57652 388516
rect 57716 388452 57717 388516
rect 57651 388451 57717 388452
rect 57467 270332 57533 270333
rect 57467 270268 57468 270332
rect 57532 270268 57533 270332
rect 57467 270267 57533 270268
rect 57467 252516 57533 252517
rect 57467 252452 57468 252516
rect 57532 252452 57533 252516
rect 57467 252451 57533 252452
rect 57283 252380 57349 252381
rect 57283 252316 57284 252380
rect 57348 252316 57349 252380
rect 57283 252315 57349 252316
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57286 164253 57346 252315
rect 57283 164252 57349 164253
rect 57283 164188 57284 164252
rect 57348 164188 57349 164252
rect 57283 164187 57349 164188
rect 57283 140860 57349 140861
rect 57283 140796 57284 140860
rect 57348 140796 57349 140860
rect 57283 140795 57349 140796
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 56268 55693 56269
rect 55627 56204 55628 56268
rect 55692 56204 55693 56268
rect 55627 56203 55693 56204
rect 53603 54908 53669 54909
rect 53603 54844 53604 54908
rect 53668 54844 53669 54908
rect 53603 54843 53669 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57286 56133 57346 140795
rect 57470 70413 57530 252451
rect 57654 175133 57714 388451
rect 57651 175132 57717 175133
rect 57651 175068 57652 175132
rect 57716 175068 57717 175132
rect 57651 175067 57717 175068
rect 57838 166973 57898 485147
rect 59123 484940 59189 484941
rect 59123 484876 59124 484940
rect 59188 484876 59189 484940
rect 59123 484875 59189 484876
rect 58939 469844 59005 469845
rect 58939 469780 58940 469844
rect 59004 469780 59005 469844
rect 58939 469779 59005 469780
rect 58755 468348 58821 468349
rect 58755 468284 58756 468348
rect 58820 468284 58821 468348
rect 58755 468283 58821 468284
rect 58571 465628 58637 465629
rect 58571 465564 58572 465628
rect 58636 465564 58637 465628
rect 58571 465563 58637 465564
rect 57835 166972 57901 166973
rect 57835 166908 57836 166972
rect 57900 166908 57901 166972
rect 57835 166907 57901 166908
rect 57651 164116 57717 164117
rect 57651 164052 57652 164116
rect 57716 164052 57717 164116
rect 57651 164051 57717 164052
rect 57467 70412 57533 70413
rect 57467 70348 57468 70412
rect 57532 70348 57533 70412
rect 57467 70347 57533 70348
rect 57654 59533 57714 164051
rect 57835 163980 57901 163981
rect 57835 163916 57836 163980
rect 57900 163916 57901 163980
rect 57835 163915 57901 163916
rect 57651 59532 57717 59533
rect 57651 59468 57652 59532
rect 57716 59468 57717 59532
rect 57651 59467 57717 59468
rect 57283 56132 57349 56133
rect 57283 56068 57284 56132
rect 57348 56068 57349 56132
rect 57283 56067 57349 56068
rect 57838 54773 57898 163915
rect 58574 57357 58634 465563
rect 58571 57356 58637 57357
rect 58571 57292 58572 57356
rect 58636 57292 58637 57356
rect 58571 57291 58637 57292
rect 58758 57221 58818 468283
rect 58755 57220 58821 57221
rect 58755 57156 58756 57220
rect 58820 57156 58821 57220
rect 58755 57155 58821 57156
rect 58942 57085 59002 469779
rect 59126 58445 59186 484875
rect 59307 484804 59373 484805
rect 59307 484740 59308 484804
rect 59372 484740 59373 484804
rect 59307 484739 59373 484740
rect 59310 58717 59370 484739
rect 59514 476114 60134 486000
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 60134 476114
rect 59514 475794 60134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 60134 475794
rect 59514 466308 60134 475558
rect 63234 477954 63854 486000
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 63854 477954
rect 63234 477634 63854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 63854 477634
rect 60227 467124 60293 467125
rect 60227 467060 60228 467124
rect 60292 467060 60293 467124
rect 60227 467059 60293 467060
rect 60230 464810 60290 467059
rect 63234 466308 63854 477398
rect 66954 481674 67574 486000
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 67574 481674
rect 66954 481354 67574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 67574 481354
rect 66954 466308 67574 481118
rect 73794 471454 74414 486000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 466308 74414 470898
rect 77514 475174 78134 486000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 466308 78134 474618
rect 81234 478894 81854 486000
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 466308 81854 478338
rect 84954 482614 85574 486000
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 466308 85574 482058
rect 91794 472394 92414 486000
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 92414 472394
rect 91794 472074 92414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 92414 472074
rect 91794 466308 92414 471838
rect 95514 476114 96134 486000
rect 95514 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 96134 476114
rect 95514 475794 96134 475878
rect 95514 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 96134 475794
rect 95514 466308 96134 475558
rect 99234 477954 99854 486000
rect 99234 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 99854 477954
rect 99234 477634 99854 477718
rect 99234 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 99854 477634
rect 99234 466308 99854 477398
rect 102954 481674 103574 486000
rect 102954 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 103574 481674
rect 102954 481354 103574 481438
rect 102954 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 103574 481354
rect 102954 466308 103574 481118
rect 109794 471454 110414 486000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 466308 110414 470898
rect 113514 475174 114134 486000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 466308 114134 474618
rect 117234 478894 117854 486000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 466308 117854 478338
rect 120954 482614 121574 486000
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 466308 121574 482058
rect 127794 472394 128414 486000
rect 127794 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 128414 472394
rect 127794 472074 128414 472158
rect 127794 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 128414 472074
rect 127794 466308 128414 471838
rect 131514 476114 132134 486000
rect 131514 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 132134 476114
rect 131514 475794 132134 475878
rect 131514 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 132134 475794
rect 131514 466308 132134 475558
rect 135234 477954 135854 486000
rect 135234 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 135854 477954
rect 135234 477634 135854 477718
rect 135234 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 135854 477634
rect 135234 466308 135854 477398
rect 138954 481674 139574 486000
rect 138954 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 139574 481674
rect 138954 481354 139574 481438
rect 138954 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 139574 481354
rect 138954 466308 139574 481118
rect 145794 471454 146414 486000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 466308 146414 470898
rect 149514 475174 150134 486000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 466308 150134 474618
rect 153234 478894 153854 486000
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 466308 153854 478338
rect 156954 482614 157574 486000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 466308 157574 482058
rect 163794 472394 164414 486000
rect 163794 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 164414 472394
rect 163794 472074 164414 472158
rect 163794 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 164414 472074
rect 163794 466308 164414 471838
rect 167514 476114 168134 486000
rect 167514 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 168134 476114
rect 167514 475794 168134 475878
rect 167514 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 168134 475794
rect 167514 466308 168134 475558
rect 171234 477954 171854 486000
rect 171234 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 171854 477954
rect 171234 477634 171854 477718
rect 171234 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 171854 477634
rect 171234 466308 171854 477398
rect 174954 481674 175574 486000
rect 174954 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 175574 481674
rect 174954 481354 175574 481438
rect 174954 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 175574 481354
rect 174954 466308 175574 481118
rect 181794 471454 182414 486000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 466988 179709 466989
rect 179643 466924 179644 466988
rect 179708 466924 179709 466988
rect 179643 466923 179709 466924
rect 178355 466580 178421 466581
rect 178355 466516 178356 466580
rect 178420 466516 178421 466580
rect 178355 466515 178421 466516
rect 59862 464750 60290 464810
rect 178358 464810 178418 466515
rect 179646 464810 179706 466923
rect 181794 466308 182414 470898
rect 185514 475174 186134 486000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 466308 186134 474618
rect 189234 478894 189854 486000
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 466308 189854 478338
rect 192954 482614 193574 486000
rect 199331 485756 199397 485757
rect 199331 485692 199332 485756
rect 199396 485692 199397 485756
rect 199331 485691 199397 485692
rect 198227 485620 198293 485621
rect 198227 485556 198228 485620
rect 198292 485556 198293 485620
rect 198227 485555 198293 485556
rect 198043 485484 198109 485485
rect 198043 485420 198044 485484
rect 198108 485420 198109 485484
rect 198043 485419 198109 485420
rect 197859 485348 197925 485349
rect 197859 485284 197860 485348
rect 197924 485284 197925 485348
rect 197859 485283 197925 485284
rect 196571 484940 196637 484941
rect 196571 484876 196572 484940
rect 196636 484876 196637 484940
rect 196571 484875 196637 484876
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190867 466580 190933 466581
rect 190867 466516 190868 466580
rect 190932 466516 190933 466580
rect 190867 466515 190933 466516
rect 190870 464810 190930 466515
rect 192954 466308 193574 482058
rect 178358 464750 178524 464810
rect 179646 464750 179748 464810
rect 59862 379810 59922 464750
rect 178464 464202 178524 464750
rect 179688 464202 179748 464750
rect 190840 464750 190930 464810
rect 190840 464202 190900 464750
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 76056 380765 76116 381106
rect 76053 380764 76119 380765
rect 76053 380700 76054 380764
rect 76118 380700 76119 380764
rect 76053 380699 76119 380700
rect 77144 380490 77204 381106
rect 78232 380490 78292 381106
rect 79592 380490 79652 381106
rect 80544 380490 80604 381106
rect 77144 380430 77218 380490
rect 78232 380430 78322 380490
rect 59862 379750 60290 379810
rect 59514 368114 60134 379000
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 60134 368114
rect 59514 367794 60134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 60134 367794
rect 59514 359308 60134 367558
rect 60230 358730 60290 379750
rect 63234 369954 63854 379000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 359308 63854 369398
rect 66954 373674 67574 379000
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 67574 373674
rect 66954 373354 67574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 67574 373354
rect 66954 359308 67574 373118
rect 73794 363454 74414 379000
rect 77158 378997 77218 380430
rect 78262 379405 78322 380430
rect 79550 380430 79652 380490
rect 80470 380430 80604 380490
rect 81768 380490 81828 381106
rect 83128 380629 83188 381106
rect 83125 380628 83191 380629
rect 83125 380564 83126 380628
rect 83190 380564 83191 380628
rect 83125 380563 83191 380564
rect 84216 380490 84276 381106
rect 84515 380492 84581 380493
rect 84515 380490 84516 380492
rect 81768 380430 82002 380490
rect 84216 380430 84516 380490
rect 78259 379404 78325 379405
rect 78259 379340 78260 379404
rect 78324 379340 78325 379404
rect 78259 379339 78325 379340
rect 77155 378996 77221 378997
rect 77155 378932 77156 378996
rect 77220 378932 77221 378996
rect 77155 378931 77221 378932
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 359308 74414 362898
rect 77514 367174 78134 379000
rect 78262 378997 78322 379339
rect 79550 379269 79610 380430
rect 80470 379405 80530 380430
rect 80467 379404 80533 379405
rect 80467 379340 80468 379404
rect 80532 379340 80533 379404
rect 80467 379339 80533 379340
rect 79547 379268 79613 379269
rect 79547 379204 79548 379268
rect 79612 379204 79613 379268
rect 79547 379203 79613 379204
rect 78259 378996 78325 378997
rect 78259 378932 78260 378996
rect 78324 378932 78325 378996
rect 78259 378931 78325 378932
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 359308 78134 366618
rect 81234 370894 81854 379000
rect 81942 378861 82002 380430
rect 84515 380428 84516 380430
rect 84580 380428 84581 380492
rect 85440 380490 85500 381106
rect 84515 380427 84581 380428
rect 85438 380430 85500 380490
rect 86528 380490 86588 381106
rect 87616 380490 87676 381106
rect 88296 380490 88356 381106
rect 88704 380490 88764 381106
rect 90064 380490 90124 381106
rect 86528 380430 86602 380490
rect 87616 380430 87706 380490
rect 88296 380430 88442 380490
rect 88704 380430 88810 380490
rect 85438 379405 85498 380430
rect 86542 379405 86602 380430
rect 87646 379405 87706 380430
rect 88382 379405 88442 380430
rect 88750 379405 88810 380430
rect 90038 380430 90124 380490
rect 90744 380490 90804 381106
rect 91288 380490 91348 381106
rect 92376 380490 92436 381106
rect 93464 380490 93524 381106
rect 90744 380430 90834 380490
rect 91288 380430 91386 380490
rect 92376 380430 92490 380490
rect 85435 379404 85501 379405
rect 85435 379340 85436 379404
rect 85500 379340 85501 379404
rect 85435 379339 85501 379340
rect 86539 379404 86605 379405
rect 86539 379340 86540 379404
rect 86604 379340 86605 379404
rect 86539 379339 86605 379340
rect 87643 379404 87709 379405
rect 87643 379340 87644 379404
rect 87708 379340 87709 379404
rect 87643 379339 87709 379340
rect 88379 379404 88445 379405
rect 88379 379340 88380 379404
rect 88444 379340 88445 379404
rect 88379 379339 88445 379340
rect 88747 379404 88813 379405
rect 88747 379340 88748 379404
rect 88812 379340 88813 379404
rect 88747 379339 88813 379340
rect 90038 379269 90098 380430
rect 90774 379405 90834 380430
rect 91326 379405 91386 380430
rect 92430 379405 92490 380430
rect 93350 380430 93524 380490
rect 93600 380490 93660 381106
rect 94552 380490 94612 381106
rect 95912 380490 95972 381106
rect 96048 380490 96108 381106
rect 97000 380490 97060 381106
rect 98088 380490 98148 381106
rect 98496 380490 98556 381106
rect 99448 380490 99508 381106
rect 93600 380430 93778 380490
rect 94552 380430 94698 380490
rect 95912 380430 95986 380490
rect 96048 380430 96170 380490
rect 97000 380430 97090 380490
rect 98088 380430 98194 380490
rect 98496 380430 98562 380490
rect 93350 379405 93410 380430
rect 90771 379404 90837 379405
rect 90771 379340 90772 379404
rect 90836 379340 90837 379404
rect 90771 379339 90837 379340
rect 91323 379404 91389 379405
rect 91323 379340 91324 379404
rect 91388 379340 91389 379404
rect 91323 379339 91389 379340
rect 92427 379404 92493 379405
rect 92427 379340 92428 379404
rect 92492 379340 92493 379404
rect 92427 379339 92493 379340
rect 93347 379404 93413 379405
rect 93347 379340 93348 379404
rect 93412 379340 93413 379404
rect 93347 379339 93413 379340
rect 93718 379269 93778 380430
rect 90035 379268 90101 379269
rect 90035 379204 90036 379268
rect 90100 379204 90101 379268
rect 90035 379203 90101 379204
rect 93715 379268 93781 379269
rect 93715 379204 93716 379268
rect 93780 379204 93781 379268
rect 93715 379203 93781 379204
rect 81939 378860 82005 378861
rect 81939 378796 81940 378860
rect 82004 378796 82005 378860
rect 81939 378795 82005 378796
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 359308 81854 370338
rect 84954 374614 85574 379000
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 359308 85574 374058
rect 91794 364394 92414 379000
rect 94638 378589 94698 380430
rect 95926 379269 95986 380430
rect 96110 379405 96170 380430
rect 96107 379404 96173 379405
rect 96107 379340 96108 379404
rect 96172 379340 96173 379404
rect 96107 379339 96173 379340
rect 95923 379268 95989 379269
rect 95923 379204 95924 379268
rect 95988 379204 95989 379268
rect 95923 379203 95989 379204
rect 94635 378588 94701 378589
rect 94635 378524 94636 378588
rect 94700 378524 94701 378588
rect 94635 378523 94701 378524
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 359308 92414 363838
rect 95514 368114 96134 379000
rect 97030 378589 97090 380430
rect 98134 379269 98194 380430
rect 98502 379405 98562 380430
rect 99422 380430 99508 380490
rect 100672 380490 100732 381106
rect 101080 380490 101140 381106
rect 100672 380430 100770 380490
rect 98499 379404 98565 379405
rect 98499 379340 98500 379404
rect 98564 379340 98565 379404
rect 98499 379339 98565 379340
rect 99422 379269 99482 380430
rect 98131 379268 98197 379269
rect 98131 379204 98132 379268
rect 98196 379204 98197 379268
rect 98131 379203 98197 379204
rect 99419 379268 99485 379269
rect 99419 379204 99420 379268
rect 99484 379204 99485 379268
rect 99419 379203 99485 379204
rect 97027 378588 97093 378589
rect 97027 378524 97028 378588
rect 97092 378524 97093 378588
rect 97027 378523 97093 378524
rect 95514 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 96134 368114
rect 95514 367794 96134 367878
rect 95514 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 96134 367794
rect 95514 359308 96134 367558
rect 99234 369954 99854 379000
rect 100710 378453 100770 380430
rect 101078 380430 101140 380490
rect 101760 380490 101820 381106
rect 102848 380490 102908 381106
rect 103528 380490 103588 381106
rect 101760 380430 101874 380490
rect 102848 380430 102978 380490
rect 101078 379405 101138 380430
rect 101075 379404 101141 379405
rect 101075 379340 101076 379404
rect 101140 379340 101141 379404
rect 101075 379339 101141 379340
rect 100707 378452 100773 378453
rect 100707 378388 100708 378452
rect 100772 378388 100773 378452
rect 100707 378387 100773 378388
rect 101814 378317 101874 380430
rect 102918 379269 102978 380430
rect 103286 380430 103588 380490
rect 103936 380490 103996 381106
rect 105296 380490 105356 381106
rect 105976 380490 106036 381106
rect 103936 380430 104082 380490
rect 105296 380430 105370 380490
rect 103286 379405 103346 380430
rect 103283 379404 103349 379405
rect 103283 379340 103284 379404
rect 103348 379340 103349 379404
rect 103283 379339 103349 379340
rect 102915 379268 102981 379269
rect 102915 379204 102916 379268
rect 102980 379204 102981 379268
rect 102915 379203 102981 379204
rect 101811 378316 101877 378317
rect 101811 378252 101812 378316
rect 101876 378252 101877 378316
rect 101811 378251 101877 378252
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 359308 99854 369398
rect 102954 373674 103574 379000
rect 104022 378453 104082 380430
rect 105310 379405 105370 380430
rect 105862 380430 106036 380490
rect 106384 380490 106444 381106
rect 107608 380490 107668 381106
rect 108288 380490 108348 381106
rect 106384 380430 106474 380490
rect 105862 380357 105922 380430
rect 105859 380356 105925 380357
rect 105859 380292 105860 380356
rect 105924 380292 105925 380356
rect 105859 380291 105925 380292
rect 105307 379404 105373 379405
rect 105307 379340 105308 379404
rect 105372 379340 105373 379404
rect 105307 379339 105373 379340
rect 104019 378452 104085 378453
rect 104019 378388 104020 378452
rect 104084 378388 104085 378452
rect 104019 378387 104085 378388
rect 106414 378181 106474 380430
rect 107518 380430 107668 380490
rect 108254 380430 108348 380490
rect 108696 380490 108756 381106
rect 109784 380490 109844 381106
rect 108696 380430 108866 380490
rect 107518 378181 107578 380430
rect 108254 379405 108314 380430
rect 108806 379405 108866 380430
rect 109726 380430 109844 380490
rect 111008 380490 111068 381106
rect 111144 380490 111204 381106
rect 112232 380490 112292 381106
rect 113320 380490 113380 381106
rect 113592 380490 113652 381106
rect 111008 380430 111074 380490
rect 111144 380430 111258 380490
rect 112232 380430 112362 380490
rect 113320 380430 113466 380490
rect 108251 379404 108317 379405
rect 108251 379340 108252 379404
rect 108316 379340 108317 379404
rect 108251 379339 108317 379340
rect 108803 379404 108869 379405
rect 108803 379340 108804 379404
rect 108868 379340 108869 379404
rect 108803 379339 108869 379340
rect 109726 379269 109786 380430
rect 111014 380357 111074 380430
rect 111011 380356 111077 380357
rect 111011 380292 111012 380356
rect 111076 380292 111077 380356
rect 111011 380291 111077 380292
rect 111198 379405 111258 380430
rect 112302 379405 112362 380430
rect 113406 379405 113466 380430
rect 113590 380430 113652 380490
rect 114408 380490 114468 381106
rect 115768 380490 115828 381106
rect 116040 380490 116100 381106
rect 114408 380430 114570 380490
rect 115768 380430 115858 380490
rect 113590 380357 113650 380430
rect 113587 380356 113653 380357
rect 113587 380292 113588 380356
rect 113652 380292 113653 380356
rect 113587 380291 113653 380292
rect 114510 379405 114570 380430
rect 115798 379405 115858 380430
rect 115982 380430 116100 380490
rect 116992 380490 117052 381106
rect 118080 380490 118140 381106
rect 118488 380490 118548 381106
rect 119168 380490 119228 381106
rect 116992 380430 117146 380490
rect 118080 380430 118250 380490
rect 115982 380357 116042 380430
rect 115979 380356 116045 380357
rect 115979 380292 115980 380356
rect 116044 380292 116045 380356
rect 115979 380291 116045 380292
rect 111195 379404 111261 379405
rect 111195 379340 111196 379404
rect 111260 379340 111261 379404
rect 111195 379339 111261 379340
rect 112299 379404 112365 379405
rect 112299 379340 112300 379404
rect 112364 379340 112365 379404
rect 112299 379339 112365 379340
rect 113403 379404 113469 379405
rect 113403 379340 113404 379404
rect 113468 379340 113469 379404
rect 113403 379339 113469 379340
rect 114507 379404 114573 379405
rect 114507 379340 114508 379404
rect 114572 379340 114573 379404
rect 114507 379339 114573 379340
rect 115795 379404 115861 379405
rect 115795 379340 115796 379404
rect 115860 379340 115861 379404
rect 115795 379339 115861 379340
rect 109723 379268 109789 379269
rect 109723 379204 109724 379268
rect 109788 379204 109789 379268
rect 109723 379203 109789 379204
rect 106411 378180 106477 378181
rect 106411 378116 106412 378180
rect 106476 378116 106477 378180
rect 106411 378115 106477 378116
rect 107515 378180 107581 378181
rect 107515 378116 107516 378180
rect 107580 378116 107581 378180
rect 107515 378115 107581 378116
rect 102954 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 103574 373674
rect 102954 373354 103574 373438
rect 102954 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 103574 373354
rect 102954 359308 103574 373118
rect 109794 363454 110414 379000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 359308 110414 362898
rect 113514 367174 114134 379000
rect 117086 378589 117146 380430
rect 117083 378588 117149 378589
rect 117083 378524 117084 378588
rect 117148 378524 117149 378588
rect 117083 378523 117149 378524
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 359308 114134 366618
rect 117234 370894 117854 379000
rect 118190 378317 118250 380430
rect 118374 380430 118548 380490
rect 119110 380430 119228 380490
rect 120936 380490 120996 381106
rect 123520 380490 123580 381106
rect 125968 380490 126028 381106
rect 120936 380430 121010 380490
rect 123520 380430 123586 380490
rect 118374 380357 118434 380430
rect 118371 380356 118437 380357
rect 118371 380292 118372 380356
rect 118436 380292 118437 380356
rect 118371 380291 118437 380292
rect 119110 380221 119170 380430
rect 120950 380357 121010 380430
rect 123526 380357 123586 380430
rect 125918 380430 126028 380490
rect 128280 380490 128340 381106
rect 131000 380490 131060 381106
rect 133448 380490 133508 381106
rect 135896 380490 135956 381106
rect 138480 380490 138540 381106
rect 128280 380430 128370 380490
rect 131000 380430 131130 380490
rect 133448 380430 133522 380490
rect 120947 380356 121013 380357
rect 120947 380292 120948 380356
rect 121012 380292 121013 380356
rect 120947 380291 121013 380292
rect 123523 380356 123589 380357
rect 123523 380292 123524 380356
rect 123588 380292 123589 380356
rect 123523 380291 123589 380292
rect 119107 380220 119173 380221
rect 119107 380156 119108 380220
rect 119172 380156 119173 380220
rect 119107 380155 119173 380156
rect 118187 378316 118253 378317
rect 118187 378252 118188 378316
rect 118252 378252 118253 378316
rect 118187 378251 118253 378252
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 359308 117854 370338
rect 120954 374614 121574 379000
rect 125918 378453 125978 380430
rect 128310 380357 128370 380430
rect 128307 380356 128373 380357
rect 128307 380292 128308 380356
rect 128372 380292 128373 380356
rect 128307 380291 128373 380292
rect 125915 378452 125981 378453
rect 125915 378388 125916 378452
rect 125980 378388 125981 378452
rect 125915 378387 125981 378388
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 359308 121574 374058
rect 127794 364394 128414 379000
rect 131070 378453 131130 380430
rect 133462 380357 133522 380430
rect 135854 380430 135956 380490
rect 138430 380430 138540 380490
rect 140928 380490 140988 381106
rect 143512 380490 143572 381106
rect 145960 380490 146020 381106
rect 148544 380490 148604 381106
rect 150992 380490 151052 381106
rect 140928 380430 141066 380490
rect 143512 380430 143642 380490
rect 145960 380430 146034 380490
rect 148544 380430 148610 380490
rect 135854 380357 135914 380430
rect 138430 380357 138490 380430
rect 133459 380356 133525 380357
rect 133459 380292 133460 380356
rect 133524 380292 133525 380356
rect 133459 380291 133525 380292
rect 135851 380356 135917 380357
rect 135851 380292 135852 380356
rect 135916 380292 135917 380356
rect 135851 380291 135917 380292
rect 138427 380356 138493 380357
rect 138427 380292 138428 380356
rect 138492 380292 138493 380356
rect 138427 380291 138493 380292
rect 141006 379405 141066 380430
rect 143582 379405 143642 380430
rect 145974 379405 146034 380430
rect 148550 380357 148610 380430
rect 150942 380430 151052 380490
rect 153440 380490 153500 381106
rect 155888 380490 155948 381106
rect 158472 380490 158532 381106
rect 160920 380490 160980 381106
rect 153440 380430 153578 380490
rect 155888 380430 155970 380490
rect 158472 380430 158546 380490
rect 148547 380356 148613 380357
rect 148547 380292 148548 380356
rect 148612 380292 148613 380356
rect 148547 380291 148613 380292
rect 150942 379405 151002 380430
rect 153518 379405 153578 380430
rect 155910 380357 155970 380430
rect 158486 380357 158546 380430
rect 160878 380430 160980 380490
rect 163368 380490 163428 381106
rect 165952 380490 166012 381106
rect 183224 380490 183284 381106
rect 163368 380430 163514 380490
rect 165952 380430 166090 380490
rect 160878 380357 160938 380430
rect 163454 380357 163514 380430
rect 166030 380357 166090 380430
rect 183142 380430 183284 380490
rect 183360 380490 183420 381106
rect 183360 380430 183570 380490
rect 155907 380356 155973 380357
rect 155907 380292 155908 380356
rect 155972 380292 155973 380356
rect 155907 380291 155973 380292
rect 158483 380356 158549 380357
rect 158483 380292 158484 380356
rect 158548 380292 158549 380356
rect 158483 380291 158549 380292
rect 160875 380356 160941 380357
rect 160875 380292 160876 380356
rect 160940 380292 160941 380356
rect 160875 380291 160941 380292
rect 163451 380356 163517 380357
rect 163451 380292 163452 380356
rect 163516 380292 163517 380356
rect 163451 380291 163517 380292
rect 166027 380356 166093 380357
rect 166027 380292 166028 380356
rect 166092 380292 166093 380356
rect 166027 380291 166093 380292
rect 141003 379404 141069 379405
rect 141003 379340 141004 379404
rect 141068 379340 141069 379404
rect 141003 379339 141069 379340
rect 143579 379404 143645 379405
rect 143579 379340 143580 379404
rect 143644 379340 143645 379404
rect 143579 379339 143645 379340
rect 145971 379404 146037 379405
rect 145971 379340 145972 379404
rect 146036 379340 146037 379404
rect 145971 379339 146037 379340
rect 150939 379404 151005 379405
rect 150939 379340 150940 379404
rect 151004 379340 151005 379404
rect 150939 379339 151005 379340
rect 153515 379404 153581 379405
rect 153515 379340 153516 379404
rect 153580 379340 153581 379404
rect 153515 379339 153581 379340
rect 131067 378452 131133 378453
rect 131067 378388 131068 378452
rect 131132 378388 131133 378452
rect 131067 378387 131133 378388
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 359308 128414 363838
rect 131514 368114 132134 379000
rect 131514 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 132134 368114
rect 131514 367794 132134 367878
rect 131514 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 132134 367794
rect 131514 359308 132134 367558
rect 135234 369954 135854 379000
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 359308 135854 369398
rect 138954 373674 139574 379000
rect 138954 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 139574 373674
rect 138954 373354 139574 373438
rect 138954 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 139574 373354
rect 138954 359308 139574 373118
rect 145794 363454 146414 379000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 359308 146414 362898
rect 149514 367174 150134 379000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 359308 150134 366618
rect 153234 370894 153854 379000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 359308 153854 370338
rect 156954 374614 157574 379000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 359308 157574 374058
rect 163794 364394 164414 379000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 359308 164414 363838
rect 167514 368114 168134 379000
rect 167514 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 168134 368114
rect 167514 367794 168134 367878
rect 167514 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 168134 367794
rect 167514 359308 168134 367558
rect 171234 369954 171854 379000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 359308 171854 369398
rect 174954 373674 175574 379000
rect 174954 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 175574 373674
rect 174954 373354 175574 373438
rect 174954 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 175574 373354
rect 174954 359308 175574 373118
rect 181794 363454 182414 379000
rect 183142 378453 183202 380430
rect 183139 378452 183205 378453
rect 183139 378388 183140 378452
rect 183204 378388 183205 378452
rect 183139 378387 183205 378388
rect 183510 378181 183570 380430
rect 183507 378180 183573 378181
rect 183507 378116 183508 378180
rect 183572 378116 183573 378180
rect 183507 378115 183573 378116
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 359308 182414 362898
rect 185514 367174 186134 379000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 359308 186134 366618
rect 189234 370894 189854 379000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 359308 189854 370338
rect 192954 374614 193574 379000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 359308 193574 374058
rect 178539 358868 178605 358869
rect 178539 358804 178540 358868
rect 178604 358804 178605 358868
rect 178539 358803 178605 358804
rect 179643 358868 179709 358869
rect 179643 358804 179644 358868
rect 179708 358804 179709 358868
rect 179643 358803 179709 358804
rect 190867 358868 190933 358869
rect 190867 358804 190868 358868
rect 190932 358804 190933 358868
rect 190867 358803 190933 358804
rect 59862 358670 60290 358730
rect 59862 272370 59922 358670
rect 178542 358050 178602 358803
rect 178464 357990 178602 358050
rect 179646 358050 179706 358803
rect 190870 358050 190930 358803
rect 179646 357990 179748 358050
rect 178464 357202 178524 357990
rect 179688 357202 179748 357990
rect 190840 357990 190930 358050
rect 190840 357202 190900 357990
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 76056 273730 76116 274040
rect 76054 273670 76116 273730
rect 77144 273730 77204 274040
rect 78232 273730 78292 274040
rect 79592 273730 79652 274040
rect 80544 273730 80604 274040
rect 77144 273670 77218 273730
rect 78232 273670 78322 273730
rect 76054 272917 76114 273670
rect 76051 272916 76117 272917
rect 76051 272852 76052 272916
rect 76116 272852 76117 272916
rect 76051 272851 76117 272852
rect 59862 272310 60290 272370
rect 59514 260114 60134 272000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 252308 60134 259558
rect 60230 251970 60290 272310
rect 63234 261954 63854 272000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 252308 63854 261398
rect 66954 265674 67574 272000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 252308 67574 265118
rect 73794 255454 74414 272000
rect 77158 271829 77218 273670
rect 77155 271828 77221 271829
rect 77155 271764 77156 271828
rect 77220 271764 77221 271828
rect 77155 271763 77221 271764
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 252308 74414 254898
rect 77514 259174 78134 272000
rect 78262 271149 78322 273670
rect 79550 273670 79652 273730
rect 80470 273670 80604 273730
rect 81768 273730 81828 274040
rect 83128 273730 83188 274040
rect 84216 273730 84276 274040
rect 85440 273730 85500 274040
rect 81768 273670 82002 273730
rect 78259 271148 78325 271149
rect 78259 271084 78260 271148
rect 78324 271084 78325 271148
rect 78259 271083 78325 271084
rect 79550 271013 79610 273670
rect 80470 271557 80530 273670
rect 80467 271556 80533 271557
rect 80467 271492 80468 271556
rect 80532 271492 80533 271556
rect 80467 271491 80533 271492
rect 79547 271012 79613 271013
rect 79547 270948 79548 271012
rect 79612 270948 79613 271012
rect 79547 270947 79613 270948
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 252308 78134 258618
rect 81234 262894 81854 272000
rect 81942 271693 82002 273670
rect 83046 273670 83188 273730
rect 83966 273670 84276 273730
rect 84702 273670 85500 273730
rect 86528 273730 86588 274040
rect 87616 273730 87676 274040
rect 88296 273730 88356 274040
rect 88704 273730 88764 274040
rect 90064 273730 90124 274040
rect 86528 273670 86602 273730
rect 87616 273670 87706 273730
rect 88296 273670 88442 273730
rect 88704 273670 88810 273730
rect 83046 271829 83106 273670
rect 83966 271829 84026 273670
rect 83043 271828 83109 271829
rect 83043 271764 83044 271828
rect 83108 271764 83109 271828
rect 83043 271763 83109 271764
rect 83963 271828 84029 271829
rect 83963 271764 83964 271828
rect 84028 271764 84029 271828
rect 83963 271763 84029 271764
rect 84702 271693 84762 273670
rect 81939 271692 82005 271693
rect 81939 271628 81940 271692
rect 82004 271628 82005 271692
rect 81939 271627 82005 271628
rect 84699 271692 84765 271693
rect 84699 271628 84700 271692
rect 84764 271628 84765 271692
rect 84699 271627 84765 271628
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 252308 81854 262338
rect 84954 266614 85574 272000
rect 86542 270877 86602 273670
rect 87646 271829 87706 273670
rect 87643 271828 87709 271829
rect 87643 271764 87644 271828
rect 87708 271764 87709 271828
rect 87643 271763 87709 271764
rect 88382 271149 88442 273670
rect 88379 271148 88445 271149
rect 88379 271084 88380 271148
rect 88444 271084 88445 271148
rect 88379 271083 88445 271084
rect 88750 271013 88810 273670
rect 90038 273670 90124 273730
rect 90744 273730 90804 274040
rect 91288 273730 91348 274040
rect 92376 273730 92436 274040
rect 93464 273730 93524 274040
rect 90744 273670 90834 273730
rect 91288 273670 91386 273730
rect 90038 271013 90098 273670
rect 90774 272917 90834 273670
rect 90771 272916 90837 272917
rect 90771 272852 90772 272916
rect 90836 272852 90837 272916
rect 90771 272851 90837 272852
rect 88747 271012 88813 271013
rect 88747 270948 88748 271012
rect 88812 270948 88813 271012
rect 88747 270947 88813 270948
rect 90035 271012 90101 271013
rect 90035 270948 90036 271012
rect 90100 270948 90101 271012
rect 90035 270947 90101 270948
rect 86539 270876 86605 270877
rect 86539 270812 86540 270876
rect 86604 270812 86605 270876
rect 86539 270811 86605 270812
rect 91326 270605 91386 273670
rect 91510 273670 92436 273730
rect 93350 273670 93524 273730
rect 93600 273730 93660 274040
rect 94552 273730 94612 274040
rect 95912 273869 95972 274040
rect 95909 273868 95975 273869
rect 95909 273804 95910 273868
rect 95974 273804 95975 273868
rect 95909 273803 95975 273804
rect 96048 273730 96108 274040
rect 93600 273670 93778 273730
rect 91323 270604 91389 270605
rect 91323 270540 91324 270604
rect 91388 270540 91389 270604
rect 91323 270539 91389 270540
rect 91510 270469 91570 273670
rect 91507 270468 91573 270469
rect 91507 270404 91508 270468
rect 91572 270404 91573 270468
rect 91507 270403 91573 270404
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 252308 85574 266058
rect 91794 256394 92414 272000
rect 93350 270877 93410 273670
rect 93718 272917 93778 273670
rect 94454 273670 94612 273730
rect 95926 273670 96108 273730
rect 97000 273730 97060 274040
rect 98088 273730 98148 274040
rect 98496 273730 98556 274040
rect 99448 273730 99508 274040
rect 97000 273670 97090 273730
rect 98088 273670 98194 273730
rect 98496 273670 98562 273730
rect 93715 272916 93781 272917
rect 93715 272852 93716 272916
rect 93780 272852 93781 272916
rect 93715 272851 93781 272852
rect 94454 271829 94514 273670
rect 95926 272917 95986 273670
rect 95923 272916 95989 272917
rect 95923 272852 95924 272916
rect 95988 272852 95989 272916
rect 95923 272851 95989 272852
rect 97030 272373 97090 273670
rect 97027 272372 97093 272373
rect 97027 272308 97028 272372
rect 97092 272308 97093 272372
rect 97027 272307 97093 272308
rect 94451 271828 94517 271829
rect 94451 271764 94452 271828
rect 94516 271764 94517 271828
rect 94451 271763 94517 271764
rect 93347 270876 93413 270877
rect 93347 270812 93348 270876
rect 93412 270812 93413 270876
rect 93347 270811 93413 270812
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 252308 92414 255838
rect 95514 260114 96134 272000
rect 98134 271829 98194 273670
rect 98502 272917 98562 273670
rect 99422 273670 99508 273730
rect 100672 273730 100732 274040
rect 101080 273730 101140 274040
rect 100672 273670 100770 273730
rect 99422 272917 99482 273670
rect 100710 273189 100770 273670
rect 101078 273670 101140 273730
rect 101760 273730 101820 274040
rect 102848 273730 102908 274040
rect 101760 273670 101874 273730
rect 100707 273188 100773 273189
rect 100707 273124 100708 273188
rect 100772 273124 100773 273188
rect 100707 273123 100773 273124
rect 98499 272916 98565 272917
rect 98499 272852 98500 272916
rect 98564 272852 98565 272916
rect 98499 272851 98565 272852
rect 99419 272916 99485 272917
rect 99419 272852 99420 272916
rect 99484 272852 99485 272916
rect 99419 272851 99485 272852
rect 98131 271828 98197 271829
rect 98131 271764 98132 271828
rect 98196 271764 98197 271828
rect 98131 271763 98197 271764
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 252308 96134 259558
rect 99234 261954 99854 272000
rect 101078 271421 101138 273670
rect 101814 271829 101874 273670
rect 102734 273670 102908 273730
rect 103528 273730 103588 274040
rect 103936 273730 103996 274040
rect 103528 273670 103714 273730
rect 102734 273053 102794 273670
rect 102731 273052 102797 273053
rect 102731 272988 102732 273052
rect 102796 272988 102797 273052
rect 102731 272987 102797 272988
rect 101811 271828 101877 271829
rect 101811 271764 101812 271828
rect 101876 271764 101877 271828
rect 101811 271763 101877 271764
rect 101075 271420 101141 271421
rect 101075 271356 101076 271420
rect 101140 271356 101141 271420
rect 101075 271355 101141 271356
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 252308 99854 261398
rect 102954 265674 103574 272000
rect 103654 271690 103714 273670
rect 103838 273670 103996 273730
rect 105296 273730 105356 274040
rect 105976 273730 106036 274040
rect 105296 273670 105370 273730
rect 103838 272781 103898 273670
rect 103835 272780 103901 272781
rect 103835 272716 103836 272780
rect 103900 272716 103901 272780
rect 103835 272715 103901 272716
rect 103835 271692 103901 271693
rect 103835 271690 103836 271692
rect 103654 271630 103836 271690
rect 103835 271628 103836 271630
rect 103900 271628 103901 271692
rect 103835 271627 103901 271628
rect 105310 270877 105370 273670
rect 105862 273670 106036 273730
rect 106384 273730 106444 274040
rect 107608 273730 107668 274040
rect 108288 273730 108348 274040
rect 108696 273730 108756 274040
rect 109784 273730 109844 274040
rect 106384 273670 106474 273730
rect 105862 271421 105922 273670
rect 105859 271420 105925 271421
rect 105859 271356 105860 271420
rect 105924 271356 105925 271420
rect 105859 271355 105925 271356
rect 106414 270877 106474 273670
rect 107518 273670 107668 273730
rect 108254 273670 108348 273730
rect 108622 273670 108756 273730
rect 109542 273670 109844 273730
rect 107518 271013 107578 273670
rect 107515 271012 107581 271013
rect 107515 270948 107516 271012
rect 107580 270948 107581 271012
rect 107515 270947 107581 270948
rect 105307 270876 105373 270877
rect 105307 270812 105308 270876
rect 105372 270812 105373 270876
rect 105307 270811 105373 270812
rect 106411 270876 106477 270877
rect 106411 270812 106412 270876
rect 106476 270812 106477 270876
rect 106411 270811 106477 270812
rect 108254 270605 108314 273670
rect 108622 271013 108682 273670
rect 108619 271012 108685 271013
rect 108619 270948 108620 271012
rect 108684 270948 108685 271012
rect 108619 270947 108685 270948
rect 109542 270605 109602 273670
rect 111008 273597 111068 274040
rect 111144 273730 111204 274040
rect 112232 273730 112292 274040
rect 113320 273730 113380 274040
rect 113592 273730 113652 274040
rect 111144 273670 111258 273730
rect 111005 273596 111071 273597
rect 111005 273532 111006 273596
rect 111070 273532 111071 273596
rect 111005 273531 111071 273532
rect 108251 270604 108317 270605
rect 108251 270540 108252 270604
rect 108316 270540 108317 270604
rect 108251 270539 108317 270540
rect 109539 270604 109605 270605
rect 109539 270540 109540 270604
rect 109604 270540 109605 270604
rect 109539 270539 109605 270540
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 252308 103574 265118
rect 109794 255454 110414 272000
rect 111198 270741 111258 273670
rect 112118 273670 112292 273730
rect 113222 273670 113380 273730
rect 113590 273670 113652 273730
rect 114408 273730 114468 274040
rect 115768 273730 115828 274040
rect 116040 273730 116100 274040
rect 114408 273670 114570 273730
rect 115768 273670 115858 273730
rect 112118 271013 112178 273670
rect 112115 271012 112181 271013
rect 112115 270948 112116 271012
rect 112180 270948 112181 271012
rect 112115 270947 112181 270948
rect 111195 270740 111261 270741
rect 111195 270676 111196 270740
rect 111260 270676 111261 270740
rect 111195 270675 111261 270676
rect 113222 270605 113282 273670
rect 113590 272237 113650 273670
rect 113587 272236 113653 272237
rect 113587 272172 113588 272236
rect 113652 272172 113653 272236
rect 113587 272171 113653 272172
rect 113219 270604 113285 270605
rect 113219 270540 113220 270604
rect 113284 270540 113285 270604
rect 113219 270539 113285 270540
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 252308 110414 254898
rect 113514 259174 114134 272000
rect 114510 271829 114570 273670
rect 114507 271828 114573 271829
rect 114507 271764 114508 271828
rect 114572 271764 114573 271828
rect 114507 271763 114573 271764
rect 115798 270605 115858 273670
rect 115982 273670 116100 273730
rect 116992 273730 117052 274040
rect 118080 273730 118140 274040
rect 118488 273730 118548 274040
rect 119168 273730 119228 274040
rect 120936 273730 120996 274040
rect 116992 273670 117146 273730
rect 115982 271557 116042 273670
rect 115979 271556 116045 271557
rect 115979 271492 115980 271556
rect 116044 271492 116045 271556
rect 115979 271491 116045 271492
rect 117086 270605 117146 273670
rect 118006 273670 118140 273730
rect 118374 273670 118548 273730
rect 119110 273670 119228 273730
rect 120766 273670 120996 273730
rect 123520 273730 123580 274040
rect 125968 273730 126028 274040
rect 123520 273670 123586 273730
rect 118006 272645 118066 273670
rect 118003 272644 118069 272645
rect 118003 272580 118004 272644
rect 118068 272580 118069 272644
rect 118003 272579 118069 272580
rect 115795 270604 115861 270605
rect 115795 270540 115796 270604
rect 115860 270540 115861 270604
rect 115795 270539 115861 270540
rect 117083 270604 117149 270605
rect 117083 270540 117084 270604
rect 117148 270540 117149 270604
rect 117083 270539 117149 270540
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 252308 114134 258618
rect 117234 262894 117854 272000
rect 118374 271557 118434 273670
rect 119110 272509 119170 273670
rect 119107 272508 119173 272509
rect 119107 272444 119108 272508
rect 119172 272444 119173 272508
rect 119107 272443 119173 272444
rect 120766 271693 120826 273670
rect 120763 271692 120829 271693
rect 120763 271628 120764 271692
rect 120828 271628 120829 271692
rect 120763 271627 120829 271628
rect 118371 271556 118437 271557
rect 118371 271492 118372 271556
rect 118436 271492 118437 271556
rect 118371 271491 118437 271492
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 252308 117854 262338
rect 120954 266614 121574 272000
rect 123526 271829 123586 273670
rect 125918 273670 126028 273730
rect 128280 273730 128340 274040
rect 131000 273730 131060 274040
rect 128280 273670 128738 273730
rect 123523 271828 123589 271829
rect 123523 271764 123524 271828
rect 123588 271764 123589 271828
rect 123523 271763 123589 271764
rect 125918 271693 125978 273670
rect 125915 271692 125981 271693
rect 125915 271628 125916 271692
rect 125980 271628 125981 271692
rect 125915 271627 125981 271628
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 252308 121574 266058
rect 127794 256394 128414 272000
rect 128678 271829 128738 273670
rect 130886 273670 131060 273730
rect 130886 271829 130946 273670
rect 133448 273597 133508 274040
rect 135896 273597 135956 274040
rect 138480 273597 138540 274040
rect 140928 273597 140988 274040
rect 143512 273730 143572 274040
rect 145960 273730 146020 274040
rect 143512 273670 143642 273730
rect 133445 273596 133511 273597
rect 133445 273532 133446 273596
rect 133510 273532 133511 273596
rect 133445 273531 133511 273532
rect 135893 273596 135959 273597
rect 135893 273532 135894 273596
rect 135958 273532 135959 273596
rect 135893 273531 135959 273532
rect 138477 273596 138543 273597
rect 138477 273532 138478 273596
rect 138542 273532 138543 273596
rect 138477 273531 138543 273532
rect 140925 273596 140991 273597
rect 140925 273532 140926 273596
rect 140990 273532 140991 273596
rect 140925 273531 140991 273532
rect 143582 272645 143642 273670
rect 145606 273670 146020 273730
rect 148544 273730 148604 274040
rect 150992 273730 151052 274040
rect 148544 273670 148610 273730
rect 143579 272644 143645 272645
rect 143579 272580 143580 272644
rect 143644 272580 143645 272644
rect 143579 272579 143645 272580
rect 128675 271828 128741 271829
rect 128675 271764 128676 271828
rect 128740 271764 128741 271828
rect 128675 271763 128741 271764
rect 130883 271828 130949 271829
rect 130883 271764 130884 271828
rect 130948 271764 130949 271828
rect 130883 271763 130949 271764
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 252308 128414 255838
rect 131514 260114 132134 272000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 252308 132134 259558
rect 135234 261954 135854 272000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 252308 135854 261398
rect 138954 265674 139574 272000
rect 145606 270605 145666 273670
rect 145603 270604 145669 270605
rect 145603 270540 145604 270604
rect 145668 270540 145669 270604
rect 145603 270539 145669 270540
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 252308 139574 265118
rect 145794 255454 146414 272000
rect 148550 270605 148610 273670
rect 150942 273670 151052 273730
rect 153440 273730 153500 274040
rect 155888 273730 155948 274040
rect 158472 273730 158532 274040
rect 160920 273730 160980 274040
rect 153440 273670 154130 273730
rect 155888 273670 155970 273730
rect 158472 273670 158546 273730
rect 148547 270604 148613 270605
rect 148547 270540 148548 270604
rect 148612 270540 148613 270604
rect 148547 270539 148613 270540
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 252308 146414 254898
rect 149514 259174 150134 272000
rect 150942 271829 151002 273670
rect 150939 271828 151005 271829
rect 150939 271764 150940 271828
rect 151004 271764 151005 271828
rect 150939 271763 151005 271764
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 252308 150134 258618
rect 153234 262894 153854 272000
rect 154070 271829 154130 273670
rect 155910 271829 155970 273670
rect 154067 271828 154133 271829
rect 154067 271764 154068 271828
rect 154132 271764 154133 271828
rect 154067 271763 154133 271764
rect 155907 271828 155973 271829
rect 155907 271764 155908 271828
rect 155972 271764 155973 271828
rect 155907 271763 155973 271764
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 252308 153854 262338
rect 156954 266614 157574 272000
rect 158486 271693 158546 273670
rect 160878 273670 160980 273730
rect 163368 273730 163428 274040
rect 165952 273730 166012 274040
rect 183224 273730 183284 274040
rect 163368 273670 163514 273730
rect 165952 273670 166090 273730
rect 160878 271693 160938 273670
rect 163454 271693 163514 273670
rect 158483 271692 158549 271693
rect 158483 271628 158484 271692
rect 158548 271628 158549 271692
rect 158483 271627 158549 271628
rect 160875 271692 160941 271693
rect 160875 271628 160876 271692
rect 160940 271628 160941 271692
rect 160875 271627 160941 271628
rect 163451 271692 163517 271693
rect 163451 271628 163452 271692
rect 163516 271628 163517 271692
rect 163451 271627 163517 271628
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 252308 157574 266058
rect 163794 256394 164414 272000
rect 166030 271693 166090 273670
rect 183142 273670 183284 273730
rect 183360 273730 183420 274040
rect 183360 273670 183570 273730
rect 166027 271692 166093 271693
rect 166027 271628 166028 271692
rect 166092 271628 166093 271692
rect 166027 271627 166093 271628
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 252308 164414 255838
rect 167514 260114 168134 272000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 252308 168134 259558
rect 171234 261954 171854 272000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 252308 171854 261398
rect 174954 265674 175574 272000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 252308 175574 265118
rect 181794 255454 182414 272000
rect 183142 271421 183202 273670
rect 183139 271420 183205 271421
rect 183139 271356 183140 271420
rect 183204 271356 183205 271420
rect 183139 271355 183205 271356
rect 183510 271149 183570 273670
rect 196574 273053 196634 484875
rect 196755 474196 196821 474197
rect 196755 474132 196756 474196
rect 196820 474132 196821 474196
rect 196755 474131 196821 474132
rect 196571 273052 196637 273053
rect 196571 272988 196572 273052
rect 196636 272988 196637 273052
rect 196571 272987 196637 272988
rect 183507 271148 183573 271149
rect 183507 271084 183508 271148
rect 183572 271084 183573 271148
rect 183507 271083 183573 271084
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 178539 253196 178605 253197
rect 178539 253132 178540 253196
rect 178604 253132 178605 253196
rect 178539 253131 178605 253132
rect 179643 253196 179709 253197
rect 179643 253132 179644 253196
rect 179708 253132 179709 253196
rect 179643 253131 179709 253132
rect 59862 251910 60290 251970
rect 59862 166290 59922 251910
rect 178542 250610 178602 253131
rect 178464 250550 178602 250610
rect 179646 250610 179706 253131
rect 181794 252308 182414 254898
rect 185514 259174 186134 272000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 252308 186134 258618
rect 189234 262894 189854 272000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252308 189854 262338
rect 192954 266614 193574 272000
rect 196758 271829 196818 474131
rect 196755 271828 196821 271829
rect 196755 271764 196756 271828
rect 196820 271764 196821 271828
rect 196755 271763 196821 271764
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 190867 253740 190933 253741
rect 190867 253676 190868 253740
rect 190932 253676 190933 253740
rect 190867 253675 190933 253676
rect 190870 250610 190930 253675
rect 192954 252308 193574 266058
rect 179646 250550 179748 250610
rect 178464 250240 178524 250550
rect 179688 250240 179748 250550
rect 190840 250550 190930 250610
rect 190840 250240 190900 250550
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 166290 76116 167106
rect 59862 166230 60290 166290
rect 59514 152114 60134 165000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 60230 145210 60290 166230
rect 76054 166230 76116 166290
rect 77144 166290 77204 167106
rect 78232 166290 78292 167106
rect 79592 166290 79652 167106
rect 80544 167010 80604 167106
rect 81768 167010 81828 167106
rect 83128 167010 83188 167106
rect 84216 167010 84276 167106
rect 85440 167010 85500 167106
rect 77144 166230 77218 166290
rect 78232 166230 78322 166290
rect 63234 155834 63854 165000
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 63854 155834
rect 63234 155514 63854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 63854 155514
rect 63234 145308 63854 155278
rect 66954 157674 67574 165000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 165000
rect 76054 164253 76114 166230
rect 77158 164389 77218 166230
rect 77155 164388 77221 164389
rect 77155 164324 77156 164388
rect 77220 164324 77221 164388
rect 77155 164323 77221 164324
rect 76051 164252 76117 164253
rect 76051 164188 76052 164252
rect 76116 164188 76117 164252
rect 76051 164187 76117 164188
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 165000
rect 78262 164253 78322 166230
rect 79550 166230 79652 166290
rect 80470 166950 80604 167010
rect 81758 166950 81828 167010
rect 83046 166950 83188 167010
rect 84150 166950 84276 167010
rect 85438 166950 85500 167010
rect 86528 167010 86588 167106
rect 87616 167010 87676 167106
rect 88296 167010 88356 167106
rect 88704 167010 88764 167106
rect 90064 167010 90124 167106
rect 86528 166950 86602 167010
rect 87616 166950 87706 167010
rect 88296 166950 88442 167010
rect 88704 166950 88810 167010
rect 79550 164933 79610 166230
rect 79547 164932 79613 164933
rect 79547 164868 79548 164932
rect 79612 164868 79613 164932
rect 79547 164867 79613 164868
rect 80470 164253 80530 166950
rect 81758 165613 81818 166950
rect 81755 165612 81821 165613
rect 81755 165548 81756 165612
rect 81820 165548 81821 165612
rect 81755 165547 81821 165548
rect 78259 164252 78325 164253
rect 78259 164188 78260 164252
rect 78324 164188 78325 164252
rect 78259 164187 78325 164188
rect 80467 164252 80533 164253
rect 80467 164188 80468 164252
rect 80532 164188 80533 164252
rect 80467 164187 80533 164188
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 165000
rect 83046 164253 83106 166950
rect 84150 164253 84210 166950
rect 85438 165613 85498 166950
rect 85435 165612 85501 165613
rect 85435 165548 85436 165612
rect 85500 165548 85501 165612
rect 85435 165547 85501 165548
rect 83043 164252 83109 164253
rect 83043 164188 83044 164252
rect 83108 164188 83109 164252
rect 83043 164187 83109 164188
rect 84147 164252 84213 164253
rect 84147 164188 84148 164252
rect 84212 164188 84213 164252
rect 84147 164187 84213 164188
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 165000
rect 86542 164253 86602 166950
rect 87646 164253 87706 166950
rect 88382 164933 88442 166950
rect 88379 164932 88445 164933
rect 88379 164868 88380 164932
rect 88444 164868 88445 164932
rect 88379 164867 88445 164868
rect 88750 164253 88810 166950
rect 90038 166950 90124 167010
rect 90744 167010 90804 167106
rect 91288 167010 91348 167106
rect 92376 167010 92436 167106
rect 93464 167010 93524 167106
rect 90744 166950 90834 167010
rect 91288 166950 91386 167010
rect 92376 166950 92490 167010
rect 90038 164253 90098 166950
rect 90774 165069 90834 166950
rect 90771 165068 90837 165069
rect 90771 165004 90772 165068
rect 90836 165004 90837 165068
rect 90771 165003 90837 165004
rect 91326 164253 91386 166950
rect 92430 165613 92490 166950
rect 93350 166950 93524 167010
rect 93600 167010 93660 167106
rect 94552 167010 94612 167106
rect 95912 167010 95972 167106
rect 93600 166950 93778 167010
rect 92427 165612 92493 165613
rect 92427 165548 92428 165612
rect 92492 165548 92493 165612
rect 92427 165547 92493 165548
rect 86539 164252 86605 164253
rect 86539 164188 86540 164252
rect 86604 164188 86605 164252
rect 86539 164187 86605 164188
rect 87643 164252 87709 164253
rect 87643 164188 87644 164252
rect 87708 164188 87709 164252
rect 87643 164187 87709 164188
rect 88747 164252 88813 164253
rect 88747 164188 88748 164252
rect 88812 164188 88813 164252
rect 88747 164187 88813 164188
rect 90035 164252 90101 164253
rect 90035 164188 90036 164252
rect 90100 164188 90101 164252
rect 90035 164187 90101 164188
rect 91323 164252 91389 164253
rect 91323 164188 91324 164252
rect 91388 164188 91389 164252
rect 91323 164187 91389 164188
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 165000
rect 93350 164253 93410 166950
rect 93718 164933 93778 166950
rect 94454 166950 94612 167010
rect 95742 166950 95972 167010
rect 96048 167010 96108 167106
rect 97000 167010 97060 167106
rect 98088 167010 98148 167106
rect 98496 167010 98556 167106
rect 96048 166950 96170 167010
rect 97000 166950 97090 167010
rect 98088 166950 98194 167010
rect 98496 166950 98562 167010
rect 93715 164932 93781 164933
rect 93715 164868 93716 164932
rect 93780 164868 93781 164932
rect 93715 164867 93781 164868
rect 94454 164253 94514 166950
rect 95742 165613 95802 166950
rect 96110 166293 96170 166950
rect 96107 166292 96173 166293
rect 96107 166228 96108 166292
rect 96172 166228 96173 166292
rect 96107 166227 96173 166228
rect 95739 165612 95805 165613
rect 95739 165548 95740 165612
rect 95804 165548 95805 165612
rect 95739 165547 95805 165548
rect 93347 164252 93413 164253
rect 93347 164188 93348 164252
rect 93412 164188 93413 164252
rect 93347 164187 93413 164188
rect 94451 164252 94517 164253
rect 94451 164188 94452 164252
rect 94516 164188 94517 164252
rect 94451 164187 94517 164188
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 165000
rect 97030 164253 97090 166950
rect 98134 164253 98194 166950
rect 98502 166293 98562 166950
rect 99448 166834 99508 167106
rect 99422 166774 99508 166834
rect 100672 166834 100732 167106
rect 101080 166837 101140 167106
rect 101077 166836 101143 166837
rect 100672 166774 100770 166834
rect 98499 166292 98565 166293
rect 98499 166228 98500 166292
rect 98564 166228 98565 166292
rect 98499 166227 98565 166228
rect 99422 165613 99482 166774
rect 100710 165613 100770 166774
rect 101077 166772 101078 166836
rect 101142 166772 101143 166836
rect 101760 166834 101820 167106
rect 102848 166834 102908 167106
rect 103528 166837 103588 167106
rect 101760 166774 101874 166834
rect 101077 166771 101143 166772
rect 99419 165612 99485 165613
rect 99419 165548 99420 165612
rect 99484 165548 99485 165612
rect 99419 165547 99485 165548
rect 100707 165612 100773 165613
rect 100707 165548 100708 165612
rect 100772 165548 100773 165612
rect 100707 165547 100773 165548
rect 97027 164252 97093 164253
rect 97027 164188 97028 164252
rect 97092 164188 97093 164252
rect 97027 164187 97093 164188
rect 98131 164252 98197 164253
rect 98131 164188 98132 164252
rect 98196 164188 98197 164252
rect 98131 164187 98197 164188
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 155834 99854 165000
rect 101814 164253 101874 166774
rect 102734 166774 102908 166834
rect 103525 166836 103591 166837
rect 102734 164253 102794 166774
rect 103525 166772 103526 166836
rect 103590 166772 103591 166836
rect 103525 166771 103591 166772
rect 103936 166290 103996 167106
rect 103838 166230 103996 166290
rect 105296 166290 105356 167106
rect 105976 166290 106036 167106
rect 105296 166230 105370 166290
rect 101811 164252 101877 164253
rect 101811 164188 101812 164252
rect 101876 164188 101877 164252
rect 101811 164187 101877 164188
rect 102731 164252 102797 164253
rect 102731 164188 102732 164252
rect 102796 164188 102797 164252
rect 102731 164187 102797 164188
rect 99234 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 99854 155834
rect 99234 155514 99854 155598
rect 99234 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 99854 155514
rect 99234 145308 99854 155278
rect 102954 157674 103574 165000
rect 103838 164253 103898 166230
rect 105310 165613 105370 166230
rect 105862 166230 106036 166290
rect 106384 166290 106444 167106
rect 107608 166565 107668 167106
rect 108288 166837 108348 167106
rect 108285 166836 108351 166837
rect 108285 166772 108286 166836
rect 108350 166772 108351 166836
rect 108285 166771 108351 166772
rect 107605 166564 107671 166565
rect 107605 166500 107606 166564
rect 107670 166500 107671 166564
rect 107605 166499 107671 166500
rect 108696 166290 108756 167106
rect 109784 166290 109844 167106
rect 106384 166230 106474 166290
rect 105862 165613 105922 166230
rect 106414 165613 106474 166230
rect 108622 166230 108756 166290
rect 109726 166230 109844 166290
rect 111008 166290 111068 167106
rect 111144 166290 111204 167106
rect 112232 166290 112292 167106
rect 113320 166290 113380 167106
rect 113592 166290 113652 167106
rect 111008 166230 111074 166290
rect 111144 166230 111258 166290
rect 108622 165613 108682 166230
rect 109726 165613 109786 166230
rect 111014 165613 111074 166230
rect 105307 165612 105373 165613
rect 105307 165548 105308 165612
rect 105372 165548 105373 165612
rect 105307 165547 105373 165548
rect 105859 165612 105925 165613
rect 105859 165548 105860 165612
rect 105924 165548 105925 165612
rect 105859 165547 105925 165548
rect 106411 165612 106477 165613
rect 106411 165548 106412 165612
rect 106476 165548 106477 165612
rect 106411 165547 106477 165548
rect 108619 165612 108685 165613
rect 108619 165548 108620 165612
rect 108684 165548 108685 165612
rect 108619 165547 108685 165548
rect 109723 165612 109789 165613
rect 109723 165548 109724 165612
rect 109788 165548 109789 165612
rect 109723 165547 109789 165548
rect 111011 165612 111077 165613
rect 111011 165548 111012 165612
rect 111076 165548 111077 165612
rect 111011 165547 111077 165548
rect 103835 164252 103901 164253
rect 103835 164188 103836 164252
rect 103900 164188 103901 164252
rect 103835 164187 103901 164188
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 165000
rect 111198 164661 111258 166230
rect 112118 166230 112292 166290
rect 113222 166230 113380 166290
rect 113590 166230 113652 166290
rect 114408 166290 114468 167106
rect 115768 166290 115828 167106
rect 116040 166290 116100 167106
rect 114408 166230 114570 166290
rect 115768 166230 115858 166290
rect 112118 165613 112178 166230
rect 112115 165612 112181 165613
rect 112115 165548 112116 165612
rect 112180 165548 112181 165612
rect 112115 165547 112181 165548
rect 113222 165069 113282 166230
rect 113590 165613 113650 166230
rect 113587 165612 113653 165613
rect 113587 165548 113588 165612
rect 113652 165548 113653 165612
rect 113587 165547 113653 165548
rect 113219 165068 113285 165069
rect 113219 165004 113220 165068
rect 113284 165004 113285 165068
rect 113219 165003 113285 165004
rect 111195 164660 111261 164661
rect 111195 164596 111196 164660
rect 111260 164596 111261 164660
rect 111195 164595 111261 164596
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 165000
rect 114510 164933 114570 166230
rect 114507 164932 114573 164933
rect 114507 164868 114508 164932
rect 114572 164868 114573 164932
rect 114507 164867 114573 164868
rect 115798 164525 115858 166230
rect 115982 166230 116100 166290
rect 116992 166290 117052 167106
rect 118080 166290 118140 167106
rect 118488 166290 118548 167106
rect 119168 166290 119228 167106
rect 116992 166230 117146 166290
rect 115982 165613 116042 166230
rect 115979 165612 116045 165613
rect 115979 165548 115980 165612
rect 116044 165548 116045 165612
rect 115979 165547 116045 165548
rect 117086 164525 117146 166230
rect 118006 166230 118140 166290
rect 118374 166230 118548 166290
rect 119110 166230 119228 166290
rect 120936 166290 120996 167106
rect 123520 166290 123580 167106
rect 125968 166290 126028 167106
rect 128280 167010 128340 167106
rect 131000 167010 131060 167106
rect 128280 166950 128554 167010
rect 128280 166910 128370 166950
rect 120936 166230 121010 166290
rect 123520 166230 123586 166290
rect 118006 165613 118066 166230
rect 118374 165613 118434 166230
rect 119110 165613 119170 166230
rect 120950 165613 121010 166230
rect 123526 165613 123586 166230
rect 125918 166230 126028 166290
rect 125918 165613 125978 166230
rect 128494 165613 128554 166950
rect 130886 166950 131060 167010
rect 133448 167010 133508 167106
rect 135896 167010 135956 167106
rect 133448 166950 133522 167010
rect 130886 165613 130946 166950
rect 133462 165613 133522 166950
rect 135854 166950 135956 167010
rect 118003 165612 118069 165613
rect 118003 165548 118004 165612
rect 118068 165548 118069 165612
rect 118003 165547 118069 165548
rect 118371 165612 118437 165613
rect 118371 165548 118372 165612
rect 118436 165548 118437 165612
rect 118371 165547 118437 165548
rect 119107 165612 119173 165613
rect 119107 165548 119108 165612
rect 119172 165548 119173 165612
rect 119107 165547 119173 165548
rect 120947 165612 121013 165613
rect 120947 165548 120948 165612
rect 121012 165548 121013 165612
rect 120947 165547 121013 165548
rect 123523 165612 123589 165613
rect 123523 165548 123524 165612
rect 123588 165548 123589 165612
rect 123523 165547 123589 165548
rect 125915 165612 125981 165613
rect 125915 165548 125916 165612
rect 125980 165548 125981 165612
rect 125915 165547 125981 165548
rect 128491 165612 128557 165613
rect 128491 165548 128492 165612
rect 128556 165548 128557 165612
rect 128491 165547 128557 165548
rect 130883 165612 130949 165613
rect 130883 165548 130884 165612
rect 130948 165548 130949 165612
rect 130883 165547 130949 165548
rect 133459 165612 133525 165613
rect 133459 165548 133460 165612
rect 133524 165548 133525 165612
rect 133459 165547 133525 165548
rect 135854 165205 135914 166950
rect 138480 166837 138540 167106
rect 140928 166837 140988 167106
rect 143512 166837 143572 167106
rect 145960 166837 146020 167106
rect 148544 167010 148604 167106
rect 150992 167010 151052 167106
rect 153440 167010 153500 167106
rect 148544 166950 148610 167010
rect 138477 166836 138543 166837
rect 138477 166772 138478 166836
rect 138542 166772 138543 166836
rect 138477 166771 138543 166772
rect 140925 166836 140991 166837
rect 140925 166772 140926 166836
rect 140990 166772 140991 166836
rect 140925 166771 140991 166772
rect 143509 166836 143575 166837
rect 143509 166772 143510 166836
rect 143574 166772 143575 166836
rect 143509 166771 143575 166772
rect 145957 166836 146023 166837
rect 145957 166772 145958 166836
rect 146022 166772 146023 166836
rect 145957 166771 146023 166772
rect 148550 166701 148610 166950
rect 150942 166950 151052 167010
rect 153334 166950 153500 167010
rect 155888 167010 155948 167106
rect 155888 166950 155970 167010
rect 148547 166700 148613 166701
rect 148547 166636 148548 166700
rect 148612 166636 148613 166700
rect 148547 166635 148613 166636
rect 150942 166565 151002 166950
rect 153334 166565 153394 166950
rect 150939 166564 151005 166565
rect 150939 166500 150940 166564
rect 151004 166500 151005 166564
rect 150939 166499 151005 166500
rect 153331 166564 153397 166565
rect 153331 166500 153332 166564
rect 153396 166500 153397 166564
rect 153331 166499 153397 166500
rect 155910 165477 155970 166950
rect 158472 166290 158532 167106
rect 160920 166290 160980 167106
rect 163368 166701 163428 167106
rect 165952 166701 166012 167106
rect 163365 166700 163431 166701
rect 163365 166636 163366 166700
rect 163430 166636 163431 166700
rect 163365 166635 163431 166636
rect 165949 166700 166015 166701
rect 165949 166636 165950 166700
rect 166014 166636 166015 166700
rect 165949 166635 166015 166636
rect 183224 166565 183284 167106
rect 183221 166564 183287 166565
rect 183221 166500 183222 166564
rect 183286 166500 183287 166564
rect 183221 166499 183287 166500
rect 183360 166290 183420 167106
rect 158472 166230 158546 166290
rect 155907 165476 155973 165477
rect 155907 165412 155908 165476
rect 155972 165412 155973 165476
rect 155907 165411 155973 165412
rect 158486 165341 158546 166230
rect 160878 166230 160980 166290
rect 183326 166230 183420 166290
rect 158483 165340 158549 165341
rect 158483 165276 158484 165340
rect 158548 165276 158549 165340
rect 158483 165275 158549 165276
rect 135851 165204 135917 165205
rect 135851 165140 135852 165204
rect 135916 165140 135917 165204
rect 135851 165139 135917 165140
rect 115795 164524 115861 164525
rect 115795 164460 115796 164524
rect 115860 164460 115861 164524
rect 115795 164459 115861 164460
rect 117083 164524 117149 164525
rect 117083 164460 117084 164524
rect 117148 164460 117149 164524
rect 117083 164459 117149 164460
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 165000
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 165000
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 165000
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 165000
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 155834 135854 165000
rect 135234 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 135854 155834
rect 135234 155514 135854 155598
rect 135234 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 135854 155514
rect 135234 145308 135854 155278
rect 138954 157674 139574 165000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 165000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 165000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 165000
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 165000
rect 160878 164797 160938 166230
rect 183326 165613 183386 166230
rect 183323 165612 183389 165613
rect 183323 165548 183324 165612
rect 183388 165548 183389 165612
rect 183323 165547 183389 165548
rect 160875 164796 160941 164797
rect 160875 164732 160876 164796
rect 160940 164732 160941 164796
rect 160875 164731 160941 164732
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 165000
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 165000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 155834 171854 165000
rect 171234 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 171854 155834
rect 171234 155514 171854 155598
rect 171234 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 171854 155514
rect 171234 145308 171854 155278
rect 174954 157674 175574 165000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 165000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 165000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 165000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 165000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 145308 193574 158058
rect 59862 145150 60290 145210
rect 59862 59530 59922 145150
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 190867 144940 190933 144941
rect 190867 144876 190868 144940
rect 190932 144876 190933 144940
rect 190867 144875 190933 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 144875
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 59862 59470 60290 59530
rect 59307 58716 59373 58717
rect 59307 58652 59308 58716
rect 59372 58652 59373 58716
rect 59307 58651 59373 58652
rect 59123 58444 59189 58445
rect 59123 58380 59124 58444
rect 59188 58380 59189 58444
rect 59123 58379 59189 58380
rect 58939 57084 59005 57085
rect 58939 57020 58940 57084
rect 59004 57020 59005 57084
rect 58939 57019 59005 57020
rect 57835 54772 57901 54773
rect 57835 54708 57836 54772
rect 57900 54708 57901 54772
rect 57835 54707 57901 54708
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 60230 57629 60290 59470
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59530 80604 60106
rect 78232 59470 78322 59530
rect 60227 57628 60293 57629
rect 60227 57564 60228 57628
rect 60292 57564 60293 57628
rect 60227 57563 60293 57564
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59470 80604 59530
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84216 59530 84276 60106
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 79550 57901 79610 59470
rect 80470 57901 80530 59470
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 83966 59470 84276 59530
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59533 90124 60106
rect 90035 59532 90124 59533
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 83966 58037 84026 59470
rect 85438 58173 85498 59470
rect 85435 58172 85501 58173
rect 85435 58108 85436 58172
rect 85500 58108 85501 58172
rect 85435 58107 85501 58108
rect 83963 58036 84029 58037
rect 83963 57972 83964 58036
rect 84028 57972 84029 58036
rect 83963 57971 84029 57972
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 88382 57901 88442 59470
rect 88750 57901 88810 59470
rect 90035 59468 90036 59532
rect 90100 59470 90124 59532
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 92376 59470 92490 59530
rect 90100 59468 90101 59470
rect 90035 59467 90101 59468
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92430 58173 92490 59470
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59805 94612 60106
rect 94549 59804 94615 59805
rect 94549 59740 94550 59804
rect 94614 59740 94615 59804
rect 94549 59739 94615 59740
rect 95912 59533 95972 60106
rect 96048 59666 96108 60106
rect 96048 59606 96354 59666
rect 95912 59532 95989 59533
rect 93600 59470 93778 59530
rect 95912 59470 95924 59532
rect 92427 58172 92493 58173
rect 92427 58108 92428 58172
rect 92492 58108 92493 58172
rect 92427 58107 92493 58108
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88379 57900 88445 57901
rect 88379 57836 88380 57900
rect 88444 57836 88445 57900
rect 88379 57835 88445 57836
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93718 57901 93778 59470
rect 95923 59468 95924 59470
rect 95988 59468 95989 59532
rect 95923 59467 95989 59468
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 93715 57900 93781 57901
rect 93715 57836 93716 57900
rect 93780 57836 93781 57900
rect 93715 57835 93781 57836
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 57085 96354 59606
rect 97000 59533 97060 60106
rect 97000 59532 97093 59533
rect 97000 59470 97028 59532
rect 97027 59468 97028 59470
rect 97092 59468 97093 59532
rect 98088 59530 98148 60106
rect 98496 59530 98556 60106
rect 99448 59805 99508 60106
rect 99445 59804 99511 59805
rect 99445 59740 99446 59804
rect 99510 59740 99511 59804
rect 99445 59739 99511 59740
rect 100672 59666 100732 60106
rect 100672 59606 100770 59666
rect 100710 59533 100770 59606
rect 100707 59532 100773 59533
rect 98088 59470 98194 59530
rect 98496 59470 98562 59530
rect 97027 59467 97093 59468
rect 98134 57901 98194 59470
rect 98131 57900 98197 57901
rect 98131 57836 98132 57900
rect 98196 57836 98197 57900
rect 98131 57835 98197 57836
rect 98502 57221 98562 59470
rect 100707 59468 100708 59532
rect 100772 59468 100773 59532
rect 101080 59530 101140 60106
rect 100707 59467 100773 59468
rect 101078 59470 101140 59530
rect 101760 59533 101820 60106
rect 102848 59805 102908 60106
rect 102845 59804 102911 59805
rect 102845 59740 102846 59804
rect 102910 59740 102911 59804
rect 102845 59739 102911 59740
rect 101760 59532 101877 59533
rect 101760 59470 101812 59532
rect 101078 58445 101138 59470
rect 101811 59468 101812 59470
rect 101876 59468 101877 59532
rect 103528 59530 103588 60106
rect 103936 59530 103996 60106
rect 105296 59669 105356 60106
rect 105976 59805 106036 60106
rect 105973 59804 106039 59805
rect 105973 59740 105974 59804
rect 106038 59740 106039 59804
rect 105973 59739 106039 59740
rect 105293 59668 105359 59669
rect 105293 59604 105294 59668
rect 105358 59604 105359 59668
rect 105293 59603 105359 59604
rect 103528 59470 103714 59530
rect 101811 59467 101877 59468
rect 101075 58444 101141 58445
rect 101075 58380 101076 58444
rect 101140 58380 101141 58444
rect 101075 58379 101141 58380
rect 98499 57220 98565 57221
rect 98499 57156 98500 57220
rect 98564 57156 98565 57220
rect 98499 57155 98565 57156
rect 96291 57084 96357 57085
rect 96291 57020 96292 57084
rect 96356 57020 96357 57084
rect 96291 57019 96357 57020
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103654 57490 103714 59470
rect 103838 59470 103996 59530
rect 106384 59530 106444 60106
rect 107608 59669 107668 60106
rect 107605 59668 107671 59669
rect 107605 59604 107606 59668
rect 107670 59604 107671 59668
rect 107605 59603 107671 59604
rect 108288 59530 108348 60106
rect 108696 59530 108756 60106
rect 109784 59530 109844 60106
rect 106384 59470 106474 59530
rect 103838 57901 103898 59470
rect 103835 57900 103901 57901
rect 103835 57836 103836 57900
rect 103900 57836 103901 57900
rect 103835 57835 103901 57836
rect 106414 57493 106474 59470
rect 108254 59470 108348 59530
rect 108622 59470 108756 59530
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59530 112292 60106
rect 113320 59530 113380 60106
rect 113592 59530 113652 60106
rect 114408 59530 114468 60106
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 108254 58581 108314 59470
rect 108251 58580 108317 58581
rect 108251 58516 108252 58580
rect 108316 58516 108317 58580
rect 108251 58515 108317 58516
rect 108622 57901 108682 59470
rect 109542 57901 109602 59470
rect 111014 58853 111074 59470
rect 111011 58852 111077 58853
rect 111011 58788 111012 58852
rect 111076 58788 111077 58852
rect 111011 58787 111077 58788
rect 108619 57900 108685 57901
rect 108619 57836 108620 57900
rect 108684 57836 108685 57900
rect 108619 57835 108685 57836
rect 109539 57900 109605 57901
rect 109539 57836 109540 57900
rect 109604 57836 109605 57900
rect 109539 57835 109605 57836
rect 106411 57492 106477 57493
rect 103654 57430 103898 57490
rect 103838 57357 103898 57430
rect 106411 57428 106412 57492
rect 106476 57428 106477 57492
rect 106411 57427 106477 57428
rect 103835 57356 103901 57357
rect 103835 57292 103836 57356
rect 103900 57292 103901 57356
rect 103835 57291 103901 57292
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 111198 57493 111258 59470
rect 112118 59470 112292 59530
rect 113222 59470 113380 59530
rect 113590 59470 113652 59530
rect 114326 59470 114468 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59530 117052 60106
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 115768 59470 115858 59530
rect 112118 57901 112178 59470
rect 113222 57901 113282 59470
rect 113590 59397 113650 59470
rect 113587 59396 113653 59397
rect 113587 59332 113588 59396
rect 113652 59332 113653 59396
rect 113587 59331 113653 59332
rect 112115 57900 112181 57901
rect 112115 57836 112116 57900
rect 112180 57836 112181 57900
rect 112115 57835 112181 57836
rect 113219 57900 113285 57901
rect 113219 57836 113220 57900
rect 113284 57836 113285 57900
rect 113219 57835 113285 57836
rect 111195 57492 111261 57493
rect 111195 57428 111196 57492
rect 111260 57428 111261 57492
rect 111195 57427 111261 57428
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 114326 57901 114386 59470
rect 114323 57900 114389 57901
rect 114323 57836 114324 57900
rect 114388 57836 114389 57900
rect 114323 57835 114389 57836
rect 115798 57493 115858 59470
rect 115982 59470 116100 59530
rect 116902 59470 117052 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 120936 59530 120996 60106
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 120936 59470 121010 59530
rect 123520 59470 123586 59530
rect 115982 57901 116042 59470
rect 115979 57900 116045 57901
rect 115979 57836 115980 57900
rect 116044 57836 116045 57900
rect 115979 57835 116045 57836
rect 116902 57493 116962 59470
rect 115795 57492 115861 57493
rect 115795 57428 115796 57492
rect 115860 57428 115861 57492
rect 115795 57427 115861 57428
rect 116899 57492 116965 57493
rect 116899 57428 116900 57492
rect 116964 57428 116965 57492
rect 116899 57427 116965 57428
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57901 118066 59470
rect 118003 57900 118069 57901
rect 118003 57836 118004 57900
rect 118068 57836 118069 57900
rect 118003 57835 118069 57836
rect 118374 57357 118434 59470
rect 119110 57901 119170 59470
rect 120950 58717 121010 59470
rect 120947 58716 121013 58717
rect 120947 58652 120948 58716
rect 121012 58652 121013 58716
rect 120947 58651 121013 58652
rect 119107 57900 119173 57901
rect 119107 57836 119108 57900
rect 119172 57836 119173 57900
rect 119107 57835 119173 57836
rect 118371 57356 118437 57357
rect 118371 57292 118372 57356
rect 118436 57292 118437 57356
rect 118371 57291 118437 57292
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57901 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128370 59530
rect 123523 57900 123589 57901
rect 123523 57836 123524 57900
rect 123588 57836 123589 57900
rect 123523 57835 123589 57836
rect 125918 57629 125978 59470
rect 128310 58173 128370 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 133448 59470 133522 59530
rect 128307 58172 128373 58173
rect 128307 58108 128308 58172
rect 128372 58108 128373 58172
rect 128307 58107 128373 58108
rect 125915 57628 125981 57629
rect 125915 57564 125916 57628
rect 125980 57564 125981 57628
rect 125915 57563 125981 57564
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 56677 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 143512 59530 143572 60106
rect 145960 59530 146020 60106
rect 143512 59470 143642 59530
rect 135854 58989 135914 59470
rect 138430 58989 138490 59470
rect 140822 59125 140882 59470
rect 143582 59261 143642 59470
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 143579 59260 143645 59261
rect 143579 59196 143580 59260
rect 143644 59196 143645 59260
rect 143579 59195 143645 59196
rect 140819 59124 140885 59125
rect 140819 59060 140820 59124
rect 140884 59060 140885 59124
rect 140819 59059 140885 59060
rect 135851 58988 135917 58989
rect 135851 58924 135852 58988
rect 135916 58924 135917 58988
rect 135851 58923 135917 58924
rect 138427 58988 138493 58989
rect 138427 58924 138428 58988
rect 138492 58924 138493 58988
rect 138427 58923 138493 58924
rect 133459 56676 133525 56677
rect 133459 56612 133460 56676
rect 133524 56612 133525 56676
rect 133459 56611 133525 56612
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 56269 155970 59470
rect 155907 56268 155973 56269
rect 155907 56204 155908 56268
rect 155972 56204 155973 56268
rect 155907 56203 155973 56204
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 57629 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 160878 57629 160938 59470
rect 158483 57628 158549 57629
rect 158483 57564 158484 57628
rect 158548 57564 158549 57628
rect 158483 57563 158549 57564
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163270 56677 163330 59470
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163267 56676 163333 56677
rect 163267 56612 163268 56676
rect 163332 56612 163333 56676
rect 163267 56611 163333 56612
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57765 183202 59470
rect 183510 57901 183570 59470
rect 197862 58717 197922 485283
rect 198046 58989 198106 485419
rect 198230 166973 198290 485555
rect 199147 485348 199213 485349
rect 199147 485284 199148 485348
rect 199212 485284 199213 485348
rect 199147 485283 199213 485284
rect 198411 484940 198477 484941
rect 198411 484876 198412 484940
rect 198476 484876 198477 484940
rect 198411 484875 198477 484876
rect 198414 381037 198474 484875
rect 198779 466172 198845 466173
rect 198779 466108 198780 466172
rect 198844 466108 198845 466172
rect 198779 466107 198845 466108
rect 198411 381036 198477 381037
rect 198411 380972 198412 381036
rect 198476 380972 198477 381036
rect 198411 380971 198477 380972
rect 198782 271693 198842 466107
rect 199150 379405 199210 485283
rect 199147 379404 199213 379405
rect 199147 379340 199148 379404
rect 199212 379340 199213 379404
rect 199147 379339 199213 379340
rect 199334 273189 199394 485691
rect 199794 472394 200414 486000
rect 200619 485212 200685 485213
rect 200619 485148 200620 485212
rect 200684 485148 200685 485212
rect 200619 485147 200685 485148
rect 199794 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 200414 472394
rect 199794 472074 200414 472158
rect 199515 471884 199581 471885
rect 199515 471820 199516 471884
rect 199580 471820 199581 471884
rect 199515 471819 199581 471820
rect 199794 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 200414 472074
rect 199331 273188 199397 273189
rect 199331 273124 199332 273188
rect 199396 273124 199397 273188
rect 199331 273123 199397 273124
rect 199518 272917 199578 471819
rect 199794 453454 200414 471838
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199515 272916 199581 272917
rect 199515 272852 199516 272916
rect 199580 272852 199581 272916
rect 199515 272851 199581 272852
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 198779 271692 198845 271693
rect 198779 271628 198780 271692
rect 198844 271628 198845 271692
rect 198779 271627 198845 271628
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198227 166972 198293 166973
rect 198227 166908 198228 166972
rect 198292 166908 198293 166972
rect 198227 166907 198293 166908
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198043 58988 198109 58989
rect 198043 58924 198044 58988
rect 198108 58924 198109 58988
rect 198043 58923 198109 58924
rect 197859 58716 197925 58717
rect 197859 58652 197860 58716
rect 197924 58652 197925 58716
rect 197859 58651 197925 58652
rect 183507 57900 183573 57901
rect 183507 57836 183508 57900
rect 183572 57836 183573 57900
rect 183507 57835 183573 57836
rect 183139 57764 183205 57765
rect 183139 57700 183140 57764
rect 183204 57700 183205 57764
rect 183139 57699 183205 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 92898
rect 200622 59397 200682 485147
rect 202275 485076 202341 485077
rect 202275 485012 202276 485076
rect 202340 485012 202341 485076
rect 202275 485011 202341 485012
rect 200987 484804 201053 484805
rect 200987 484740 200988 484804
rect 201052 484740 201053 484804
rect 200987 484739 201053 484740
rect 200803 469844 200869 469845
rect 200803 469780 200804 469844
rect 200868 469780 200869 469844
rect 200803 469779 200869 469780
rect 200806 164797 200866 469779
rect 200990 379541 201050 484739
rect 201355 484532 201421 484533
rect 201355 484468 201356 484532
rect 201420 484468 201421 484532
rect 201355 484467 201421 484468
rect 200987 379540 201053 379541
rect 200987 379476 200988 379540
rect 201052 379476 201053 379540
rect 200987 379475 201053 379476
rect 200803 164796 200869 164797
rect 200803 164732 200804 164796
rect 200868 164732 200869 164796
rect 200803 164731 200869 164732
rect 200619 59396 200685 59397
rect 200619 59332 200620 59396
rect 200684 59332 200685 59396
rect 200619 59331 200685 59332
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 201358 56405 201418 484467
rect 202091 475420 202157 475421
rect 202091 475356 202092 475420
rect 202156 475356 202157 475420
rect 202091 475355 202157 475356
rect 201355 56404 201421 56405
rect 201355 56340 201356 56404
rect 201420 56340 201421 56404
rect 201355 56339 201421 56340
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 202094 3909 202154 475355
rect 202278 58581 202338 485011
rect 202459 484940 202525 484941
rect 202459 484876 202460 484940
rect 202524 484876 202525 484940
rect 202459 484875 202525 484876
rect 202462 379541 202522 484875
rect 203195 480860 203261 480861
rect 203195 480796 203196 480860
rect 203260 480796 203261 480860
rect 203195 480795 203261 480796
rect 203011 472700 203077 472701
rect 203011 472636 203012 472700
rect 203076 472636 203077 472700
rect 203011 472635 203077 472636
rect 202459 379540 202525 379541
rect 202459 379476 202460 379540
rect 202524 379476 202525 379540
rect 202459 379475 202525 379476
rect 203014 164389 203074 472635
rect 203011 164388 203077 164389
rect 203011 164324 203012 164388
rect 203076 164324 203077 164388
rect 203011 164323 203077 164324
rect 202275 58580 202341 58581
rect 202275 58516 202276 58580
rect 202340 58516 202341 58580
rect 202275 58515 202341 58516
rect 203198 57493 203258 480795
rect 203514 476114 204134 486000
rect 206875 485620 206941 485621
rect 206875 485556 206876 485620
rect 206940 485556 206941 485620
rect 206875 485555 206941 485556
rect 206323 485212 206389 485213
rect 206323 485148 206324 485212
rect 206388 485148 206389 485212
rect 206323 485147 206389 485148
rect 205035 478412 205101 478413
rect 205035 478348 205036 478412
rect 205100 478348 205101 478412
rect 205035 478347 205101 478348
rect 204851 478140 204917 478141
rect 204851 478076 204852 478140
rect 204916 478076 204917 478140
rect 204851 478075 204917 478076
rect 203514 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 204134 476114
rect 203514 475794 204134 475878
rect 203514 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 204134 475794
rect 203514 457174 204134 475558
rect 204299 472564 204365 472565
rect 204299 472500 204300 472564
rect 204364 472500 204365 472564
rect 204299 472499 204365 472500
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 204302 413949 204362 472499
rect 204299 413948 204365 413949
rect 204299 413884 204300 413948
rect 204364 413884 204365 413948
rect 204299 413883 204365 413884
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 368114 204134 384618
rect 203514 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 204134 368114
rect 203514 367794 204134 367878
rect 203514 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 204134 367794
rect 203514 349174 204134 367558
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 152114 204134 168618
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203195 57492 203261 57493
rect 203195 57428 203196 57492
rect 203260 57428 203261 57492
rect 203195 57427 203261 57428
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 202091 3908 202157 3909
rect 202091 3844 202092 3908
rect 202156 3844 202157 3908
rect 202091 3843 202157 3844
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 24618
rect 204854 3229 204914 478075
rect 205038 57357 205098 478347
rect 206139 469980 206205 469981
rect 206139 469916 206140 469980
rect 206204 469916 206205 469980
rect 206139 469915 206205 469916
rect 205219 465900 205285 465901
rect 205219 465836 205220 465900
rect 205284 465836 205285 465900
rect 205219 465835 205285 465836
rect 205222 166701 205282 465835
rect 205219 166700 205285 166701
rect 205219 166636 205220 166700
rect 205284 166636 205285 166700
rect 205219 166635 205285 166636
rect 206142 165341 206202 469915
rect 206326 379541 206386 485147
rect 206691 484532 206757 484533
rect 206691 484468 206692 484532
rect 206756 484468 206757 484532
rect 206691 484467 206757 484468
rect 206323 379540 206389 379541
rect 206323 379476 206324 379540
rect 206388 379476 206389 379540
rect 206323 379475 206389 379476
rect 206139 165340 206205 165341
rect 206139 165276 206140 165340
rect 206204 165276 206205 165340
rect 206139 165275 206205 165276
rect 206694 59261 206754 484467
rect 206691 59260 206757 59261
rect 206691 59196 206692 59260
rect 206756 59196 206757 59260
rect 206691 59195 206757 59196
rect 206878 58853 206938 485555
rect 207234 477954 207854 486000
rect 209635 485620 209701 485621
rect 209635 485556 209636 485620
rect 209700 485556 209701 485620
rect 209635 485555 209701 485556
rect 208899 479500 208965 479501
rect 208899 479436 208900 479500
rect 208964 479436 208965 479500
rect 208899 479435 208965 479436
rect 207234 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 207854 477954
rect 207234 477634 207854 477718
rect 207234 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 207854 477634
rect 207234 460894 207854 477398
rect 207979 475692 208045 475693
rect 207979 475628 207980 475692
rect 208044 475628 208045 475692
rect 207979 475627 208045 475628
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 155834 207854 172338
rect 207982 164933 208042 475627
rect 208347 467260 208413 467261
rect 208347 467196 208348 467260
rect 208412 467196 208413 467260
rect 208347 467195 208413 467196
rect 208163 464404 208229 464405
rect 208163 464340 208164 464404
rect 208228 464340 208229 464404
rect 208163 464339 208229 464340
rect 207979 164932 208045 164933
rect 207979 164868 207980 164932
rect 208044 164868 208045 164932
rect 207979 164867 208045 164868
rect 208166 164117 208226 464339
rect 208350 390693 208410 467195
rect 208347 390692 208413 390693
rect 208347 390628 208348 390692
rect 208412 390628 208413 390692
rect 208347 390627 208413 390628
rect 208163 164116 208229 164117
rect 208163 164052 208164 164116
rect 208228 164052 208229 164116
rect 208163 164051 208229 164052
rect 207234 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 207854 155834
rect 207234 155514 207854 155598
rect 207234 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 207854 155514
rect 207234 136894 207854 155278
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 58852 206941 58853
rect 206875 58788 206876 58852
rect 206940 58788 206941 58852
rect 206875 58787 206941 58788
rect 205035 57356 205101 57357
rect 205035 57292 205036 57356
rect 205100 57292 205101 57356
rect 205035 57291 205101 57292
rect 207234 28894 207854 64338
rect 208902 57629 208962 479435
rect 209638 59125 209698 485555
rect 210954 481674 211574 486000
rect 217547 485076 217613 485077
rect 217547 485012 217548 485076
rect 217612 485012 217613 485076
rect 217547 485011 217613 485012
rect 211659 484940 211725 484941
rect 211659 484876 211660 484940
rect 211724 484876 211725 484940
rect 211659 484875 211725 484876
rect 210954 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 211574 481674
rect 210954 481354 211574 481438
rect 210954 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 211574 481354
rect 210371 479500 210437 479501
rect 210371 479436 210372 479500
rect 210436 479436 210437 479500
rect 210371 479435 210437 479436
rect 209819 476780 209885 476781
rect 209819 476716 209820 476780
rect 209884 476716 209885 476780
rect 209819 476715 209885 476716
rect 209822 379269 209882 476715
rect 210003 467124 210069 467125
rect 210003 467060 210004 467124
rect 210068 467060 210069 467124
rect 210003 467059 210069 467060
rect 209819 379268 209885 379269
rect 209819 379204 209820 379268
rect 209884 379204 209885 379268
rect 209819 379203 209885 379204
rect 210006 378589 210066 467059
rect 210003 378588 210069 378589
rect 210003 378524 210004 378588
rect 210068 378524 210069 378588
rect 210003 378523 210069 378524
rect 209635 59124 209701 59125
rect 209635 59060 209636 59124
rect 209700 59060 209701 59124
rect 209635 59059 209701 59060
rect 208899 57628 208965 57629
rect 208899 57564 208900 57628
rect 208964 57564 208965 57628
rect 208899 57563 208965 57564
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 204851 3228 204917 3229
rect 204851 3164 204852 3228
rect 204916 3164 204917 3228
rect 204851 3163 204917 3164
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 210374 4045 210434 479435
rect 210954 464614 211574 481118
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210739 381036 210805 381037
rect 210739 380972 210740 381036
rect 210804 380972 210805 381036
rect 210739 380971 210805 380972
rect 210742 57765 210802 380971
rect 210954 373674 211574 392058
rect 211662 376685 211722 484875
rect 211843 484804 211909 484805
rect 211843 484740 211844 484804
rect 211908 484740 211909 484804
rect 211843 484739 211909 484740
rect 211846 377909 211906 484739
rect 216995 484532 217061 484533
rect 216995 484468 216996 484532
rect 217060 484468 217061 484532
rect 216995 484467 217061 484468
rect 216259 483988 216325 483989
rect 216259 483924 216260 483988
rect 216324 483924 216325 483988
rect 216259 483923 216325 483924
rect 213867 483852 213933 483853
rect 213867 483788 213868 483852
rect 213932 483788 213933 483852
rect 213867 483787 213933 483788
rect 212579 482492 212645 482493
rect 212579 482428 212580 482492
rect 212644 482428 212645 482492
rect 212579 482427 212645 482428
rect 212582 377909 212642 482427
rect 213131 479772 213197 479773
rect 213131 479708 213132 479772
rect 213196 479708 213197 479772
rect 213131 479707 213197 479708
rect 211843 377908 211909 377909
rect 211843 377844 211844 377908
rect 211908 377844 211909 377908
rect 211843 377843 211909 377844
rect 212579 377908 212645 377909
rect 212579 377844 212580 377908
rect 212644 377844 212645 377908
rect 212579 377843 212645 377844
rect 211659 376684 211725 376685
rect 211659 376620 211660 376684
rect 211724 376620 211725 376684
rect 211659 376619 211725 376620
rect 210954 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 211574 373674
rect 210954 373354 211574 373438
rect 210954 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 211574 373354
rect 210954 356614 211574 373118
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 157674 211574 176058
rect 213134 165477 213194 479707
rect 213315 476916 213381 476917
rect 213315 476852 213316 476916
rect 213380 476852 213381 476916
rect 213315 476851 213381 476852
rect 213131 165476 213197 165477
rect 213131 165412 213132 165476
rect 213196 165412 213197 165476
rect 213131 165411 213197 165412
rect 213318 165205 213378 476851
rect 213499 468484 213565 468485
rect 213499 468420 213500 468484
rect 213564 468420 213565 468484
rect 213499 468419 213565 468420
rect 213502 166837 213562 468419
rect 213870 376685 213930 483787
rect 214419 483716 214485 483717
rect 214419 483652 214420 483716
rect 214484 483652 214485 483716
rect 214419 483651 214485 483652
rect 213867 376684 213933 376685
rect 213867 376620 213868 376684
rect 213932 376620 213933 376684
rect 213867 376619 213933 376620
rect 213499 166836 213565 166837
rect 213499 166772 213500 166836
rect 213564 166772 213565 166836
rect 213499 166771 213565 166772
rect 213315 165204 213381 165205
rect 213315 165140 213316 165204
rect 213380 165140 213381 165204
rect 213315 165139 213381 165140
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210739 57764 210805 57765
rect 210739 57700 210740 57764
rect 210804 57700 210805 57764
rect 210739 57699 210805 57700
rect 210954 32614 211574 68058
rect 214422 57085 214482 483651
rect 215891 482356 215957 482357
rect 215891 482292 215892 482356
rect 215956 482292 215957 482356
rect 215891 482291 215957 482292
rect 215339 479636 215405 479637
rect 215339 479572 215340 479636
rect 215404 479572 215405 479636
rect 215339 479571 215405 479572
rect 214603 478276 214669 478277
rect 214603 478212 214604 478276
rect 214668 478212 214669 478276
rect 214603 478211 214669 478212
rect 214419 57084 214485 57085
rect 214419 57020 214420 57084
rect 214484 57020 214485 57084
rect 214419 57019 214485 57020
rect 214606 56677 214666 478211
rect 215342 377909 215402 479571
rect 215339 377908 215405 377909
rect 215339 377844 215340 377908
rect 215404 377844 215405 377908
rect 215339 377843 215405 377844
rect 215894 57221 215954 482291
rect 216075 474060 216141 474061
rect 216075 473996 216076 474060
rect 216140 473996 216141 474060
rect 216075 473995 216141 473996
rect 216078 68101 216138 473995
rect 216262 165069 216322 483923
rect 216998 380493 217058 484467
rect 217179 480996 217245 480997
rect 217179 480932 217180 480996
rect 217244 480932 217245 480996
rect 217179 480931 217245 480932
rect 216627 380492 216693 380493
rect 216627 380428 216628 380492
rect 216692 380428 216693 380492
rect 216627 380427 216693 380428
rect 216995 380492 217061 380493
rect 216995 380428 216996 380492
rect 217060 380428 217061 380492
rect 216995 380427 217061 380428
rect 216630 376685 216690 380427
rect 216627 376684 216693 376685
rect 216627 376620 216628 376684
rect 216692 376620 216693 376684
rect 216627 376619 216693 376620
rect 217182 271557 217242 480931
rect 217363 471748 217429 471749
rect 217363 471684 217364 471748
rect 217428 471684 217429 471748
rect 217363 471683 217429 471684
rect 217366 272781 217426 471683
rect 217550 375325 217610 485011
rect 217794 471454 218414 486000
rect 219203 485212 219269 485213
rect 219203 485148 219204 485212
rect 219268 485148 219269 485212
rect 219203 485147 219269 485148
rect 218651 475556 218717 475557
rect 218651 475492 218652 475556
rect 218716 475492 218717 475556
rect 218651 475491 218717 475492
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 466308 218414 470898
rect 217547 375324 217613 375325
rect 217547 375260 217548 375324
rect 217612 375260 217613 375324
rect 217547 375259 217613 375260
rect 217547 375052 217613 375053
rect 217547 374988 217548 375052
rect 217612 374988 217613 375052
rect 217547 374987 217613 374988
rect 217363 272780 217429 272781
rect 217363 272716 217364 272780
rect 217428 272716 217429 272780
rect 217363 272715 217429 272716
rect 217179 271556 217245 271557
rect 217179 271492 217180 271556
rect 217244 271492 217245 271556
rect 217179 271491 217245 271492
rect 217550 268429 217610 374987
rect 217794 363454 218414 379000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 359308 218414 362898
rect 217547 268428 217613 268429
rect 217547 268364 217548 268428
rect 217612 268364 217613 268428
rect 217547 268363 217613 268364
rect 217794 255454 218414 272000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 252308 218414 254898
rect 217547 251836 217613 251837
rect 217547 251772 217548 251836
rect 217612 251772 217613 251836
rect 217547 251771 217613 251772
rect 216259 165068 216325 165069
rect 216259 165004 216260 165068
rect 216324 165004 216325 165068
rect 216259 165003 216325 165004
rect 217550 162757 217610 251771
rect 217547 162756 217613 162757
rect 217547 162692 217548 162756
rect 217612 162692 217613 162756
rect 217547 162691 217613 162692
rect 217363 146436 217429 146437
rect 217363 146372 217364 146436
rect 217428 146372 217429 146436
rect 217363 146371 217429 146372
rect 216075 68100 216141 68101
rect 216075 68036 216076 68100
rect 216140 68036 216141 68100
rect 216075 68035 216141 68036
rect 215891 57220 215957 57221
rect 215891 57156 215892 57220
rect 215956 57156 215957 57220
rect 215891 57155 215957 57156
rect 214603 56676 214669 56677
rect 214603 56612 214604 56676
rect 214668 56612 214669 56676
rect 214603 56611 214669 56612
rect 217366 56269 217426 146371
rect 217550 58445 217610 162691
rect 217794 147454 218414 165000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 145308 218414 146898
rect 218654 60621 218714 475491
rect 218835 474332 218901 474333
rect 218835 474268 218836 474332
rect 218900 474268 218901 474332
rect 218835 474267 218901 474268
rect 218838 273325 218898 474267
rect 218835 273324 218901 273325
rect 218835 273260 218836 273324
rect 218900 273260 218901 273324
rect 218835 273259 218901 273260
rect 219206 60621 219266 485147
rect 219939 484532 220005 484533
rect 219939 484468 219940 484532
rect 220004 484468 220005 484532
rect 219939 484467 220005 484468
rect 218651 60620 218717 60621
rect 218651 60556 218652 60620
rect 218716 60556 218717 60620
rect 218651 60555 218717 60556
rect 219203 60620 219269 60621
rect 219203 60556 219204 60620
rect 219268 60556 219269 60620
rect 219203 60555 219269 60556
rect 217547 58444 217613 58445
rect 217547 58380 217548 58444
rect 217612 58380 217613 58444
rect 217547 58379 217613 58380
rect 217363 56268 217429 56269
rect 217363 56204 217364 56268
rect 217428 56204 217429 56268
rect 217363 56203 217429 56204
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 210371 4044 210437 4045
rect 210371 3980 210372 4044
rect 210436 3980 210437 4044
rect 210371 3979 210437 3980
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219942 56541 220002 484467
rect 221514 475174 222134 486000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 466308 222134 474618
rect 225234 478894 225854 486000
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 466308 225854 478338
rect 228954 482614 229574 486000
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 466308 229574 482058
rect 235794 472394 236414 486000
rect 235794 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 236414 472394
rect 235794 472074 236414 472158
rect 235794 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 236414 472074
rect 235794 466308 236414 471838
rect 239514 476114 240134 486000
rect 239514 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 240134 476114
rect 239514 475794 240134 475878
rect 239514 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 240134 475794
rect 239514 466308 240134 475558
rect 243234 477954 243854 486000
rect 243234 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 243854 477954
rect 243234 477634 243854 477718
rect 243234 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 243854 477634
rect 243234 466308 243854 477398
rect 246954 481674 247574 486000
rect 246954 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 247574 481674
rect 246954 481354 247574 481438
rect 246954 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 247574 481354
rect 246954 466308 247574 481118
rect 253794 471454 254414 486000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 466308 254414 470898
rect 257514 475174 258134 486000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 466308 258134 474618
rect 261234 478894 261854 486000
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 466308 261854 478338
rect 264954 482614 265574 486000
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 466308 265574 482058
rect 271794 472394 272414 486000
rect 271794 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 271794 472074 272414 472158
rect 271794 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 271794 466308 272414 471838
rect 275514 476114 276134 486000
rect 275514 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 275514 475794 276134 475878
rect 275514 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 275514 466308 276134 475558
rect 279234 477954 279854 486000
rect 279234 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 279234 477634 279854 477718
rect 279234 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 279234 466308 279854 477398
rect 282954 481674 283574 486000
rect 282954 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 282954 481354 283574 481438
rect 282954 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 282954 466308 283574 481118
rect 289794 471454 290414 486000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 466308 290414 470898
rect 293514 475174 294134 486000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 466308 294134 474618
rect 297234 478894 297854 486000
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 466308 297854 478338
rect 300954 482614 301574 486000
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 466308 301574 482058
rect 307794 466308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 466308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 641033 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 641033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 641033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 641033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 641033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 641033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 641033 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 641033 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 641033 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 641033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 641033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 641033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 641033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 641033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 641033 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 641033 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 641033 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 641033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 641033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 641033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 641033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 641033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 641033 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 641033 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 641033 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 339568 633454 339888 633486
rect 339568 633218 339610 633454
rect 339846 633218 339888 633454
rect 339568 633134 339888 633218
rect 339568 632898 339610 633134
rect 339846 632898 339888 633134
rect 339568 632866 339888 632898
rect 370288 633454 370608 633486
rect 370288 633218 370330 633454
rect 370566 633218 370608 633454
rect 370288 633134 370608 633218
rect 370288 632898 370330 633134
rect 370566 632898 370608 633134
rect 370288 632866 370608 632898
rect 401008 633454 401328 633486
rect 401008 633218 401050 633454
rect 401286 633218 401328 633454
rect 401008 633134 401328 633218
rect 401008 632898 401050 633134
rect 401286 632898 401328 633134
rect 401008 632866 401328 632898
rect 324208 615454 324528 615486
rect 324208 615218 324250 615454
rect 324486 615218 324528 615454
rect 324208 615134 324528 615218
rect 324208 614898 324250 615134
rect 324486 614898 324528 615134
rect 324208 614866 324528 614898
rect 354928 615454 355248 615486
rect 354928 615218 354970 615454
rect 355206 615218 355248 615454
rect 354928 615134 355248 615218
rect 354928 614898 354970 615134
rect 355206 614898 355248 615134
rect 354928 614866 355248 614898
rect 385648 615454 385968 615486
rect 385648 615218 385690 615454
rect 385926 615218 385968 615454
rect 385648 615134 385968 615218
rect 385648 614898 385690 615134
rect 385926 614898 385968 615134
rect 385648 614866 385968 614898
rect 416368 615454 416688 615486
rect 416368 615218 416410 615454
rect 416646 615218 416688 615454
rect 416368 615134 416688 615218
rect 416368 614898 416410 615134
rect 416646 614898 416688 615134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 430619 615092 430685 615093
rect 430619 615028 430620 615092
rect 430684 615028 430685 615092
rect 430619 615027 430685 615028
rect 416368 614866 416688 614898
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 339568 597454 339888 597486
rect 339568 597218 339610 597454
rect 339846 597218 339888 597454
rect 339568 597134 339888 597218
rect 339568 596898 339610 597134
rect 339846 596898 339888 597134
rect 339568 596866 339888 596898
rect 370288 597454 370608 597486
rect 370288 597218 370330 597454
rect 370566 597218 370608 597454
rect 370288 597134 370608 597218
rect 370288 596898 370330 597134
rect 370566 596898 370608 597134
rect 370288 596866 370608 596898
rect 401008 597454 401328 597486
rect 401008 597218 401050 597454
rect 401286 597218 401328 597454
rect 401008 597134 401328 597218
rect 401008 596898 401050 597134
rect 401286 596898 401328 597134
rect 401008 596866 401328 596898
rect 324208 579454 324528 579486
rect 324208 579218 324250 579454
rect 324486 579218 324528 579454
rect 324208 579134 324528 579218
rect 324208 578898 324250 579134
rect 324486 578898 324528 579134
rect 324208 578866 324528 578898
rect 354928 579454 355248 579486
rect 354928 579218 354970 579454
rect 355206 579218 355248 579454
rect 354928 579134 355248 579218
rect 354928 578898 354970 579134
rect 355206 578898 355248 579134
rect 354928 578866 355248 578898
rect 385648 579454 385968 579486
rect 385648 579218 385690 579454
rect 385926 579218 385968 579454
rect 385648 579134 385968 579218
rect 385648 578898 385690 579134
rect 385926 578898 385968 579134
rect 385648 578866 385968 578898
rect 416368 579454 416688 579486
rect 416368 579218 416410 579454
rect 416646 579218 416688 579454
rect 416368 579134 416688 579218
rect 416368 578898 416410 579134
rect 416646 578898 416688 579134
rect 416368 578866 416688 578898
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 339568 561454 339888 561486
rect 339568 561218 339610 561454
rect 339846 561218 339888 561454
rect 339568 561134 339888 561218
rect 339568 560898 339610 561134
rect 339846 560898 339888 561134
rect 339568 560866 339888 560898
rect 370288 561454 370608 561486
rect 370288 561218 370330 561454
rect 370566 561218 370608 561454
rect 370288 561134 370608 561218
rect 370288 560898 370330 561134
rect 370566 560898 370608 561134
rect 370288 560866 370608 560898
rect 401008 561454 401328 561486
rect 401008 561218 401050 561454
rect 401286 561218 401328 561454
rect 401008 561134 401328 561218
rect 401008 560898 401050 561134
rect 401286 560898 401328 561134
rect 401008 560866 401328 560898
rect 324208 543454 324528 543486
rect 324208 543218 324250 543454
rect 324486 543218 324528 543454
rect 324208 543134 324528 543218
rect 324208 542898 324250 543134
rect 324486 542898 324528 543134
rect 324208 542866 324528 542898
rect 354928 543454 355248 543486
rect 354928 543218 354970 543454
rect 355206 543218 355248 543454
rect 354928 543134 355248 543218
rect 354928 542898 354970 543134
rect 355206 542898 355248 543134
rect 354928 542866 355248 542898
rect 385648 543454 385968 543486
rect 385648 543218 385690 543454
rect 385926 543218 385968 543454
rect 385648 543134 385968 543218
rect 385648 542898 385690 543134
rect 385926 542898 385968 543134
rect 385648 542866 385968 542898
rect 416368 543454 416688 543486
rect 416368 543218 416410 543454
rect 416646 543218 416688 543454
rect 416368 543134 416688 543218
rect 416368 542898 416410 543134
rect 416646 542898 416688 543134
rect 416368 542866 416688 542898
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 430622 526965 430682 615027
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 430803 600812 430869 600813
rect 430803 600748 430804 600812
rect 430868 600748 430869 600812
rect 430803 600747 430869 600748
rect 430806 527101 430866 600747
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 430803 527100 430869 527101
rect 430803 527036 430804 527100
rect 430868 527036 430869 527100
rect 430803 527035 430869 527036
rect 430619 526964 430685 526965
rect 430619 526900 430620 526964
rect 430684 526900 430685 526964
rect 430619 526899 430685 526900
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 466308 315854 496338
rect 318954 500614 319574 526000
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 466308 319574 500058
rect 325794 507454 326414 526000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 466308 326414 470898
rect 329514 511174 330134 526000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 466308 330134 474618
rect 333234 514894 333854 526000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 466308 333854 478338
rect 336954 518614 337574 526000
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 466308 337574 482058
rect 343794 525454 344414 526000
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338435 466580 338501 466581
rect 338435 466516 338436 466580
rect 338500 466516 338501 466580
rect 338435 466515 338501 466516
rect 339723 466580 339789 466581
rect 339723 466516 339724 466580
rect 339788 466516 339789 466580
rect 339723 466515 339789 466516
rect 338438 464810 338498 466515
rect 339726 464810 339786 466515
rect 343794 466308 344414 488898
rect 347514 493174 348134 526000
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 466308 348134 492618
rect 351234 496894 351854 526000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 466580 351013 466581
rect 350947 466516 350948 466580
rect 351012 466516 351013 466580
rect 350947 466515 351013 466516
rect 350950 464810 351010 466515
rect 351234 466308 351854 496338
rect 354954 500614 355574 526000
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 466308 355574 500058
rect 361794 507454 362414 526000
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 360883 489156 360949 489157
rect 360883 489092 360884 489156
rect 360948 489092 360949 489156
rect 360883 489091 360949 489092
rect 360699 484940 360765 484941
rect 360699 484876 360700 484940
rect 360764 484876 360765 484940
rect 360699 484875 360765 484876
rect 359779 482628 359845 482629
rect 359779 482564 359780 482628
rect 359844 482564 359845 482628
rect 359779 482563 359845 482564
rect 359411 479772 359477 479773
rect 359411 479708 359412 479772
rect 359476 479708 359477 479772
rect 359411 479707 359477 479708
rect 357571 478412 357637 478413
rect 357571 478348 357572 478412
rect 357636 478348 357637 478412
rect 357571 478347 357637 478348
rect 338438 464750 338524 464810
rect 338464 464202 338524 464750
rect 339688 464750 339786 464810
rect 350840 464750 351010 464810
rect 339688 464202 339748 464750
rect 350840 464202 350900 464750
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 357574 417485 357634 478347
rect 357939 476916 358005 476917
rect 357939 476852 357940 476916
rect 358004 476852 358005 476916
rect 357939 476851 358005 476852
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 357571 417484 357637 417485
rect 357571 417420 357572 417484
rect 357636 417420 357637 417484
rect 357571 417419 357637 417420
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 236056 380901 236116 381106
rect 237144 380901 237204 381106
rect 236053 380900 236119 380901
rect 236053 380836 236054 380900
rect 236118 380836 236119 380900
rect 236053 380835 236119 380836
rect 237141 380900 237207 380901
rect 237141 380836 237142 380900
rect 237206 380836 237207 380900
rect 237141 380835 237207 380836
rect 238232 380490 238292 381106
rect 239592 380490 239652 381106
rect 238158 380430 238292 380490
rect 239262 380430 239652 380490
rect 240544 380490 240604 381106
rect 241768 380490 241828 381106
rect 243128 380901 243188 381106
rect 243125 380900 243191 380901
rect 243125 380836 243126 380900
rect 243190 380836 243191 380900
rect 243125 380835 243191 380836
rect 244216 380490 244276 381106
rect 245440 380901 245500 381106
rect 245437 380900 245503 380901
rect 245437 380836 245438 380900
rect 245502 380836 245503 380900
rect 245437 380835 245503 380836
rect 246528 380490 246588 381106
rect 247616 380901 247676 381106
rect 247613 380900 247679 380901
rect 247613 380836 247614 380900
rect 247678 380836 247679 380900
rect 247613 380835 247679 380836
rect 248296 380490 248356 381106
rect 248704 380490 248764 381106
rect 240544 380430 240610 380490
rect 241768 380430 241898 380490
rect 244216 380430 244290 380490
rect 221514 367174 222134 379000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 359308 222134 366618
rect 225234 370894 225854 379000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 359308 225854 370338
rect 228954 374614 229574 379000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 359308 229574 374058
rect 235794 364394 236414 379000
rect 238158 378997 238218 380430
rect 238155 378996 238221 378997
rect 238155 378932 238156 378996
rect 238220 378932 238221 378996
rect 238155 378931 238221 378932
rect 239262 378725 239322 380430
rect 240550 379133 240610 380430
rect 240547 379132 240613 379133
rect 240547 379068 240548 379132
rect 240612 379068 240613 379132
rect 240547 379067 240613 379068
rect 241467 379132 241533 379133
rect 241467 379068 241468 379132
rect 241532 379068 241533 379132
rect 241467 379067 241533 379068
rect 239259 378724 239325 378725
rect 239259 378660 239260 378724
rect 239324 378660 239325 378724
rect 239259 378659 239325 378660
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 359308 236414 363838
rect 239514 368114 240134 379000
rect 241470 378861 241530 379067
rect 241467 378860 241533 378861
rect 241467 378796 241468 378860
rect 241532 378796 241533 378860
rect 241467 378795 241533 378796
rect 241838 378317 241898 380430
rect 244230 380357 244290 380430
rect 246438 380430 246588 380490
rect 248278 380430 248356 380490
rect 248646 380430 248764 380490
rect 250064 380490 250124 381106
rect 250744 380626 250804 381106
rect 251288 380626 251348 381106
rect 250670 380566 250804 380626
rect 251222 380566 251348 380626
rect 250064 380430 250178 380490
rect 244227 380356 244293 380357
rect 244227 380292 244228 380356
rect 244292 380292 244293 380356
rect 244227 380291 244293 380292
rect 246438 379269 246498 380430
rect 246435 379268 246501 379269
rect 246435 379204 246436 379268
rect 246500 379204 246501 379268
rect 246435 379203 246501 379204
rect 241835 378316 241901 378317
rect 241835 378252 241836 378316
rect 241900 378252 241901 378316
rect 241835 378251 241901 378252
rect 239514 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 240134 368114
rect 239514 367794 240134 367878
rect 239514 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 240134 367794
rect 239514 359308 240134 367558
rect 243234 369954 243854 379000
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 359308 243854 369398
rect 246954 373674 247574 379000
rect 248278 378453 248338 380430
rect 248646 379269 248706 380430
rect 250118 379269 250178 380430
rect 248643 379268 248709 379269
rect 248643 379204 248644 379268
rect 248708 379204 248709 379268
rect 248643 379203 248709 379204
rect 250115 379268 250181 379269
rect 250115 379204 250116 379268
rect 250180 379204 250181 379268
rect 250115 379203 250181 379204
rect 250670 378453 250730 380566
rect 251222 379269 251282 380566
rect 252376 380490 252436 381106
rect 253464 380490 253524 381106
rect 252326 380430 252436 380490
rect 253430 380430 253524 380490
rect 253600 380490 253660 381106
rect 254552 380901 254612 381106
rect 255912 380901 255972 381106
rect 254549 380900 254615 380901
rect 254549 380836 254550 380900
rect 254614 380836 254615 380900
rect 254549 380835 254615 380836
rect 255909 380900 255975 380901
rect 255909 380836 255910 380900
rect 255974 380836 255975 380900
rect 255909 380835 255975 380836
rect 256048 380490 256108 381106
rect 257000 380901 257060 381106
rect 256997 380900 257063 380901
rect 256997 380836 256998 380900
rect 257062 380836 257063 380900
rect 256997 380835 257063 380836
rect 258088 380629 258148 381106
rect 258085 380628 258151 380629
rect 258085 380564 258086 380628
rect 258150 380564 258151 380628
rect 258085 380563 258151 380564
rect 258496 380490 258556 381106
rect 259448 380629 259508 381106
rect 260672 380629 260732 381106
rect 259445 380628 259511 380629
rect 259445 380564 259446 380628
rect 259510 380564 259511 380628
rect 259445 380563 259511 380564
rect 260669 380628 260735 380629
rect 260669 380564 260670 380628
rect 260734 380564 260735 380628
rect 260669 380563 260735 380564
rect 261080 380490 261140 381106
rect 261760 380490 261820 381106
rect 262848 380490 262908 381106
rect 253600 380430 253674 380490
rect 252326 379269 252386 380430
rect 253430 379269 253490 380430
rect 251219 379268 251285 379269
rect 251219 379204 251220 379268
rect 251284 379204 251285 379268
rect 251219 379203 251285 379204
rect 252323 379268 252389 379269
rect 252323 379204 252324 379268
rect 252388 379204 252389 379268
rect 252323 379203 252389 379204
rect 253427 379268 253493 379269
rect 253427 379204 253428 379268
rect 253492 379204 253493 379268
rect 253427 379203 253493 379204
rect 253614 378453 253674 380430
rect 256006 380430 256108 380490
rect 258398 380430 258556 380490
rect 260974 380430 261140 380490
rect 261710 380430 261820 380490
rect 262814 380430 262908 380490
rect 263528 380490 263588 381106
rect 263936 380765 263996 381106
rect 263933 380764 263999 380765
rect 263933 380700 263934 380764
rect 263998 380700 263999 380764
rect 263933 380699 263999 380700
rect 265296 380629 265356 381106
rect 265293 380628 265359 380629
rect 265293 380564 265294 380628
rect 265358 380564 265359 380628
rect 265293 380563 265359 380564
rect 265976 380490 266036 381106
rect 266384 380490 266444 381106
rect 267608 380490 267668 381106
rect 263528 380430 263610 380490
rect 248275 378452 248341 378453
rect 248275 378388 248276 378452
rect 248340 378388 248341 378452
rect 248275 378387 248341 378388
rect 250667 378452 250733 378453
rect 250667 378388 250668 378452
rect 250732 378388 250733 378452
rect 250667 378387 250733 378388
rect 253611 378452 253677 378453
rect 253611 378388 253612 378452
rect 253676 378388 253677 378452
rect 253611 378387 253677 378388
rect 246954 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 247574 373674
rect 246954 373354 247574 373438
rect 246954 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 247574 373354
rect 246954 359308 247574 373118
rect 253794 363454 254414 379000
rect 256006 378453 256066 380430
rect 256003 378452 256069 378453
rect 256003 378388 256004 378452
rect 256068 378388 256069 378452
rect 256003 378387 256069 378388
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 359308 254414 362898
rect 257514 367174 258134 379000
rect 258398 378453 258458 380430
rect 260974 378453 261034 380430
rect 261710 379269 261770 380430
rect 261707 379268 261773 379269
rect 261707 379204 261708 379268
rect 261772 379204 261773 379268
rect 261707 379203 261773 379204
rect 258395 378452 258461 378453
rect 258395 378388 258396 378452
rect 258460 378388 258461 378452
rect 258395 378387 258461 378388
rect 260971 378452 261037 378453
rect 260971 378388 260972 378452
rect 261036 378388 261037 378452
rect 260971 378387 261037 378388
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 359308 258134 366618
rect 261234 370894 261854 379000
rect 262814 378317 262874 380430
rect 263550 378453 263610 380430
rect 265942 380430 266036 380490
rect 266310 380430 266444 380490
rect 267598 380430 267668 380490
rect 268288 380490 268348 381106
rect 268696 380490 268756 381106
rect 269784 380901 269844 381106
rect 269781 380900 269847 380901
rect 269781 380836 269782 380900
rect 269846 380836 269847 380900
rect 269781 380835 269847 380836
rect 271008 380629 271068 381106
rect 271005 380628 271071 380629
rect 271005 380564 271006 380628
rect 271070 380564 271071 380628
rect 271005 380563 271071 380564
rect 271144 380490 271204 381106
rect 272232 380490 272292 381106
rect 273320 380490 273380 381106
rect 273592 380490 273652 381106
rect 274408 380490 274468 381106
rect 275768 380490 275828 381106
rect 276040 380901 276100 381106
rect 276037 380900 276103 380901
rect 276037 380836 276038 380900
rect 276102 380836 276103 380900
rect 276037 380835 276103 380836
rect 276992 380490 277052 381106
rect 268288 380430 268394 380490
rect 268696 380430 268762 380490
rect 263547 378452 263613 378453
rect 263547 378388 263548 378452
rect 263612 378388 263613 378452
rect 263547 378387 263613 378388
rect 262811 378316 262877 378317
rect 262811 378252 262812 378316
rect 262876 378252 262877 378316
rect 262811 378251 262877 378252
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 359308 261854 370338
rect 264954 374614 265574 379000
rect 265942 378453 266002 380430
rect 265939 378452 266005 378453
rect 265939 378388 265940 378452
rect 266004 378388 266005 378452
rect 265939 378387 266005 378388
rect 266310 378317 266370 380430
rect 267598 378317 267658 380430
rect 268334 378453 268394 380430
rect 268702 379405 268762 380430
rect 271094 380430 271204 380490
rect 272198 380430 272292 380490
rect 273302 380430 273380 380490
rect 273486 380430 273652 380490
rect 274406 380430 274468 380490
rect 275694 380430 275828 380490
rect 276982 380430 277052 380490
rect 278080 380490 278140 381106
rect 278488 380490 278548 381106
rect 278080 380430 278146 380490
rect 271094 379405 271154 380430
rect 272198 379405 272258 380430
rect 273302 379405 273362 380430
rect 268699 379404 268765 379405
rect 268699 379340 268700 379404
rect 268764 379340 268765 379404
rect 268699 379339 268765 379340
rect 271091 379404 271157 379405
rect 271091 379340 271092 379404
rect 271156 379340 271157 379404
rect 271091 379339 271157 379340
rect 272195 379404 272261 379405
rect 272195 379340 272196 379404
rect 272260 379340 272261 379404
rect 272195 379339 272261 379340
rect 273299 379404 273365 379405
rect 273299 379340 273300 379404
rect 273364 379340 273365 379404
rect 273299 379339 273365 379340
rect 273486 379269 273546 380430
rect 274406 379405 274466 380430
rect 275694 379405 275754 380430
rect 274403 379404 274469 379405
rect 274403 379340 274404 379404
rect 274468 379340 274469 379404
rect 274403 379339 274469 379340
rect 275691 379404 275757 379405
rect 275691 379340 275692 379404
rect 275756 379340 275757 379404
rect 275691 379339 275757 379340
rect 276982 379269 277042 380430
rect 273483 379268 273549 379269
rect 273483 379204 273484 379268
rect 273548 379204 273549 379268
rect 273483 379203 273549 379204
rect 276979 379268 277045 379269
rect 276979 379204 276980 379268
rect 277044 379204 277045 379268
rect 276979 379203 277045 379204
rect 268331 378452 268397 378453
rect 268331 378388 268332 378452
rect 268396 378388 268397 378452
rect 268331 378387 268397 378388
rect 266307 378316 266373 378317
rect 266307 378252 266308 378316
rect 266372 378252 266373 378316
rect 266307 378251 266373 378252
rect 267595 378316 267661 378317
rect 267595 378252 267596 378316
rect 267660 378252 267661 378316
rect 267595 378251 267661 378252
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 359308 265574 374058
rect 271794 364394 272414 379000
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 359308 272414 363838
rect 275514 368114 276134 379000
rect 278086 378589 278146 380430
rect 278454 380430 278548 380490
rect 279168 380490 279228 381106
rect 280936 380490 280996 381106
rect 283520 380490 283580 381106
rect 279168 380430 279250 380490
rect 278454 379269 278514 380430
rect 279190 379269 279250 380430
rect 280846 380430 280996 380490
rect 283422 380430 283580 380490
rect 285968 380490 286028 381106
rect 288280 380490 288340 381106
rect 291000 380490 291060 381106
rect 293448 380490 293508 381106
rect 285968 380430 286058 380490
rect 280846 379269 280906 380430
rect 283422 379269 283482 380430
rect 285998 379405 286058 380430
rect 288206 380430 288340 380490
rect 290966 380430 291060 380490
rect 293358 380430 293508 380490
rect 295896 380490 295956 381106
rect 298480 380490 298540 381106
rect 300928 380490 300988 381106
rect 303512 380490 303572 381106
rect 305960 380490 306020 381106
rect 308544 380490 308604 381106
rect 295896 380430 295994 380490
rect 298480 380430 298570 380490
rect 288206 379405 288266 380430
rect 290966 379405 291026 380430
rect 293358 379405 293418 380430
rect 295934 379405 295994 380430
rect 298510 379405 298570 380430
rect 300902 380430 300988 380490
rect 303478 380430 303572 380490
rect 305870 380430 306020 380490
rect 308446 380430 308604 380490
rect 310992 380490 311052 381106
rect 313440 380490 313500 381106
rect 315888 380490 315948 381106
rect 318472 380490 318532 381106
rect 310992 380430 311082 380490
rect 300902 379405 300962 380430
rect 303478 379405 303538 380430
rect 305870 379405 305930 380430
rect 308446 379405 308506 380430
rect 311022 379405 311082 380430
rect 313414 380430 313500 380490
rect 315806 380430 315948 380490
rect 318382 380430 318532 380490
rect 320920 380490 320980 381106
rect 323368 380490 323428 381106
rect 325952 380490 326012 381106
rect 343224 380490 343284 381106
rect 320920 380430 321018 380490
rect 313414 379405 313474 380430
rect 315806 379405 315866 380430
rect 318382 379405 318442 380430
rect 285995 379404 286061 379405
rect 285995 379340 285996 379404
rect 286060 379340 286061 379404
rect 285995 379339 286061 379340
rect 288203 379404 288269 379405
rect 288203 379340 288204 379404
rect 288268 379340 288269 379404
rect 288203 379339 288269 379340
rect 290963 379404 291029 379405
rect 290963 379340 290964 379404
rect 291028 379340 291029 379404
rect 290963 379339 291029 379340
rect 293355 379404 293421 379405
rect 293355 379340 293356 379404
rect 293420 379340 293421 379404
rect 293355 379339 293421 379340
rect 295931 379404 295997 379405
rect 295931 379340 295932 379404
rect 295996 379340 295997 379404
rect 295931 379339 295997 379340
rect 298507 379404 298573 379405
rect 298507 379340 298508 379404
rect 298572 379340 298573 379404
rect 298507 379339 298573 379340
rect 300899 379404 300965 379405
rect 300899 379340 300900 379404
rect 300964 379340 300965 379404
rect 300899 379339 300965 379340
rect 303475 379404 303541 379405
rect 303475 379340 303476 379404
rect 303540 379340 303541 379404
rect 303475 379339 303541 379340
rect 305867 379404 305933 379405
rect 305867 379340 305868 379404
rect 305932 379340 305933 379404
rect 305867 379339 305933 379340
rect 308443 379404 308509 379405
rect 308443 379340 308444 379404
rect 308508 379340 308509 379404
rect 308443 379339 308509 379340
rect 311019 379404 311085 379405
rect 311019 379340 311020 379404
rect 311084 379340 311085 379404
rect 311019 379339 311085 379340
rect 313411 379404 313477 379405
rect 313411 379340 313412 379404
rect 313476 379340 313477 379404
rect 313411 379339 313477 379340
rect 315803 379404 315869 379405
rect 315803 379340 315804 379404
rect 315868 379340 315869 379404
rect 315803 379339 315869 379340
rect 318379 379404 318445 379405
rect 318379 379340 318380 379404
rect 318444 379340 318445 379404
rect 318379 379339 318445 379340
rect 278451 379268 278517 379269
rect 278451 379204 278452 379268
rect 278516 379204 278517 379268
rect 278451 379203 278517 379204
rect 279187 379268 279253 379269
rect 279187 379204 279188 379268
rect 279252 379204 279253 379268
rect 279187 379203 279253 379204
rect 280843 379268 280909 379269
rect 280843 379204 280844 379268
rect 280908 379204 280909 379268
rect 280843 379203 280909 379204
rect 283419 379268 283485 379269
rect 283419 379204 283420 379268
rect 283484 379204 283485 379268
rect 283419 379203 283485 379204
rect 278083 378588 278149 378589
rect 278083 378524 278084 378588
rect 278148 378524 278149 378588
rect 278083 378523 278149 378524
rect 275514 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 276134 368114
rect 275514 367794 276134 367878
rect 275514 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 276134 367794
rect 275514 359308 276134 367558
rect 279234 369954 279854 379000
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 359308 279854 369398
rect 282954 373674 283574 379000
rect 282954 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 283574 373674
rect 282954 373354 283574 373438
rect 282954 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 283574 373354
rect 282954 359308 283574 373118
rect 289794 363454 290414 379000
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 359308 290414 362898
rect 293514 367174 294134 379000
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 359308 294134 366618
rect 297234 370894 297854 379000
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 359308 297854 370338
rect 300954 374614 301574 379000
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 359308 301574 374058
rect 307794 364394 308414 379000
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 359308 308414 363838
rect 311514 368114 312134 379000
rect 311514 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 312134 368114
rect 311514 367794 312134 367878
rect 311514 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 312134 367794
rect 311514 359308 312134 367558
rect 315234 369954 315854 379000
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 359308 315854 369398
rect 318954 373674 319574 379000
rect 320958 378589 321018 380430
rect 323350 380430 323428 380490
rect 325926 380430 326012 380490
rect 343222 380430 343284 380490
rect 343360 380490 343420 381106
rect 343360 380430 343466 380490
rect 323350 379405 323410 380430
rect 323347 379404 323413 379405
rect 323347 379340 323348 379404
rect 323412 379340 323413 379404
rect 323347 379339 323413 379340
rect 325926 379269 325986 380430
rect 325923 379268 325989 379269
rect 325923 379204 325924 379268
rect 325988 379204 325989 379268
rect 325923 379203 325989 379204
rect 320955 378588 321021 378589
rect 320955 378524 320956 378588
rect 321020 378524 321021 378588
rect 320955 378523 321021 378524
rect 318954 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 319574 373674
rect 318954 373354 319574 373438
rect 318954 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 319574 373354
rect 318954 359308 319574 373118
rect 325794 363454 326414 379000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 359308 326414 362898
rect 329514 367174 330134 379000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 359308 330134 366618
rect 333234 370894 333854 379000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 359308 333854 370338
rect 336954 374614 337574 379000
rect 343222 378453 343282 380430
rect 343219 378452 343285 378453
rect 343219 378388 343220 378452
rect 343284 378388 343285 378452
rect 343219 378387 343285 378388
rect 343406 378317 343466 380430
rect 343403 378316 343469 378317
rect 343403 378252 343404 378316
rect 343468 378252 343469 378316
rect 343403 378251 343469 378252
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 359308 337574 374058
rect 343794 364394 344414 379000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 359308 344414 363838
rect 347514 368114 348134 379000
rect 347514 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 348134 368114
rect 347514 367794 348134 367878
rect 347514 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 348134 367794
rect 347514 359308 348134 367558
rect 351234 369954 351854 379000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 359308 351854 369398
rect 354954 373674 355574 379000
rect 354954 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 355574 373674
rect 354954 373354 355574 373438
rect 354954 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 355574 373354
rect 354954 359308 355574 373118
rect 338435 358868 338501 358869
rect 338435 358804 338436 358868
rect 338500 358804 338501 358868
rect 338435 358803 338501 358804
rect 339723 358868 339789 358869
rect 339723 358804 339724 358868
rect 339788 358804 339789 358868
rect 339723 358803 339789 358804
rect 350947 358868 351013 358869
rect 350947 358804 350948 358868
rect 351012 358804 351013 358868
rect 350947 358803 351013 358804
rect 338438 358050 338498 358803
rect 339726 358050 339786 358803
rect 350950 358050 351010 358803
rect 338438 357990 338524 358050
rect 338464 357202 338524 357990
rect 339688 357990 339786 358050
rect 350840 357990 351010 358050
rect 339688 357202 339748 357990
rect 350840 357202 350900 357990
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 236056 273730 236116 274040
rect 237144 273730 237204 274040
rect 238232 273730 238292 274040
rect 239592 273730 239652 274040
rect 235950 273670 236116 273730
rect 237054 273670 237204 273730
rect 238158 273670 238292 273730
rect 239262 273670 239652 273730
rect 240544 273730 240604 274040
rect 241768 273730 241828 274040
rect 243128 273730 243188 274040
rect 240544 273670 240610 273730
rect 235950 272237 236010 273670
rect 235947 272236 236013 272237
rect 235947 272172 235948 272236
rect 236012 272172 236013 272236
rect 235947 272171 236013 272172
rect 221514 259174 222134 272000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252308 222134 258618
rect 225234 262894 225854 272000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252308 225854 262338
rect 228954 266614 229574 272000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252308 229574 266058
rect 235794 256394 236414 272000
rect 237054 271421 237114 273670
rect 237051 271420 237117 271421
rect 237051 271356 237052 271420
rect 237116 271356 237117 271420
rect 237051 271355 237117 271356
rect 238158 269789 238218 273670
rect 239262 270605 239322 273670
rect 239259 270604 239325 270605
rect 239259 270540 239260 270604
rect 239324 270540 239325 270604
rect 239259 270539 239325 270540
rect 238155 269788 238221 269789
rect 238155 269724 238156 269788
rect 238220 269724 238221 269788
rect 238155 269723 238221 269724
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 252308 236414 255838
rect 239514 260114 240134 272000
rect 240550 270197 240610 273670
rect 241654 273670 241828 273730
rect 242942 273670 243188 273730
rect 244216 273730 244276 274040
rect 245440 273730 245500 274040
rect 246528 273730 246588 274040
rect 244216 273670 244290 273730
rect 241654 270333 241714 273670
rect 242942 270605 243002 273670
rect 242939 270604 243005 270605
rect 242939 270540 242940 270604
rect 243004 270540 243005 270604
rect 242939 270539 243005 270540
rect 241651 270332 241717 270333
rect 241651 270268 241652 270332
rect 241716 270268 241717 270332
rect 241651 270267 241717 270268
rect 240547 270196 240613 270197
rect 240547 270132 240548 270196
rect 240612 270132 240613 270196
rect 240547 270131 240613 270132
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 252308 240134 259558
rect 243234 261954 243854 272000
rect 244230 270741 244290 273670
rect 245334 273670 245500 273730
rect 246438 273670 246588 273730
rect 247616 273730 247676 274040
rect 248296 273730 248356 274040
rect 248704 273730 248764 274040
rect 247616 273670 247786 273730
rect 244227 270740 244293 270741
rect 244227 270676 244228 270740
rect 244292 270676 244293 270740
rect 244227 270675 244293 270676
rect 245334 270605 245394 273670
rect 246438 270605 246498 273670
rect 245331 270604 245397 270605
rect 245331 270540 245332 270604
rect 245396 270540 245397 270604
rect 245331 270539 245397 270540
rect 246435 270604 246501 270605
rect 246435 270540 246436 270604
rect 246500 270540 246501 270604
rect 246435 270539 246501 270540
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 252308 243854 261398
rect 246954 265674 247574 272000
rect 247726 270605 247786 273670
rect 248278 273670 248356 273730
rect 248646 273670 248764 273730
rect 250064 273730 250124 274040
rect 250064 273670 250178 273730
rect 248278 271149 248338 273670
rect 248275 271148 248341 271149
rect 248275 271084 248276 271148
rect 248340 271084 248341 271148
rect 248275 271083 248341 271084
rect 248646 270605 248706 273670
rect 250118 270605 250178 273670
rect 250744 273597 250804 274040
rect 251288 273730 251348 274040
rect 252376 273730 252436 274040
rect 253464 273730 253524 274040
rect 251222 273670 251348 273730
rect 252326 273670 252436 273730
rect 253430 273670 253524 273730
rect 253600 273730 253660 274040
rect 254552 273730 254612 274040
rect 255912 273730 255972 274040
rect 253600 273670 253674 273730
rect 250741 273596 250807 273597
rect 250741 273532 250742 273596
rect 250806 273532 250807 273596
rect 250741 273531 250807 273532
rect 251222 270605 251282 273670
rect 252326 270741 252386 273670
rect 252323 270740 252389 270741
rect 252323 270676 252324 270740
rect 252388 270676 252389 270740
rect 252323 270675 252389 270676
rect 253430 270605 253490 273670
rect 253614 271285 253674 273670
rect 254534 273670 254612 273730
rect 255822 273670 255972 273730
rect 256048 273730 256108 274040
rect 257000 273730 257060 274040
rect 256048 273670 256250 273730
rect 253611 271284 253677 271285
rect 253611 271220 253612 271284
rect 253676 271220 253677 271284
rect 253611 271219 253677 271220
rect 247723 270604 247789 270605
rect 247723 270540 247724 270604
rect 247788 270540 247789 270604
rect 247723 270539 247789 270540
rect 248643 270604 248709 270605
rect 248643 270540 248644 270604
rect 248708 270540 248709 270604
rect 248643 270539 248709 270540
rect 250115 270604 250181 270605
rect 250115 270540 250116 270604
rect 250180 270540 250181 270604
rect 250115 270539 250181 270540
rect 251219 270604 251285 270605
rect 251219 270540 251220 270604
rect 251284 270540 251285 270604
rect 251219 270539 251285 270540
rect 253427 270604 253493 270605
rect 253427 270540 253428 270604
rect 253492 270540 253493 270604
rect 253427 270539 253493 270540
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 252308 247574 265118
rect 253794 255454 254414 272000
rect 254534 270877 254594 273670
rect 254531 270876 254597 270877
rect 254531 270812 254532 270876
rect 254596 270812 254597 270876
rect 254531 270811 254597 270812
rect 255822 270741 255882 273670
rect 256190 271149 256250 273670
rect 256926 273670 257060 273730
rect 258088 273730 258148 274040
rect 258496 273730 258556 274040
rect 258088 273670 258274 273730
rect 256187 271148 256253 271149
rect 256187 271084 256188 271148
rect 256252 271084 256253 271148
rect 256187 271083 256253 271084
rect 255819 270740 255885 270741
rect 255819 270676 255820 270740
rect 255884 270676 255885 270740
rect 255819 270675 255885 270676
rect 256926 270605 256986 273670
rect 256923 270604 256989 270605
rect 256923 270540 256924 270604
rect 256988 270540 256989 270604
rect 256923 270539 256989 270540
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252308 254414 254898
rect 257514 259174 258134 272000
rect 258214 271010 258274 273670
rect 258398 273670 258556 273730
rect 259448 273730 259508 274040
rect 260672 273730 260732 274040
rect 261080 273730 261140 274040
rect 259448 273670 259562 273730
rect 258398 271557 258458 273670
rect 258395 271556 258461 271557
rect 258395 271492 258396 271556
rect 258460 271492 258461 271556
rect 258395 271491 258461 271492
rect 258214 270950 258458 271010
rect 258398 270605 258458 270950
rect 259502 270605 259562 273670
rect 260606 273670 260732 273730
rect 260974 273670 261140 273730
rect 261760 273730 261820 274040
rect 262848 273730 262908 274040
rect 261760 273670 262138 273730
rect 260606 270741 260666 273670
rect 260974 271285 261034 273670
rect 260971 271284 261037 271285
rect 260971 271220 260972 271284
rect 261036 271220 261037 271284
rect 260971 271219 261037 271220
rect 260603 270740 260669 270741
rect 260603 270676 260604 270740
rect 260668 270676 260669 270740
rect 260603 270675 260669 270676
rect 258395 270604 258461 270605
rect 258395 270540 258396 270604
rect 258460 270540 258461 270604
rect 258395 270539 258461 270540
rect 259499 270604 259565 270605
rect 259499 270540 259500 270604
rect 259564 270540 259565 270604
rect 259499 270539 259565 270540
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252308 258134 258618
rect 261234 262894 261854 272000
rect 262078 270605 262138 273670
rect 262814 273670 262908 273730
rect 263528 273730 263588 274040
rect 263936 273730 263996 274040
rect 265296 273730 265356 274040
rect 265976 273730 266036 274040
rect 266384 273733 266444 274040
rect 263528 273670 263610 273730
rect 262814 270605 262874 273670
rect 263550 271557 263610 273670
rect 263918 273670 263996 273730
rect 265206 273670 265356 273730
rect 265942 273670 266036 273730
rect 266381 273732 266447 273733
rect 263547 271556 263613 271557
rect 263547 271492 263548 271556
rect 263612 271492 263613 271556
rect 263547 271491 263613 271492
rect 263918 270605 263978 273670
rect 265206 272237 265266 273670
rect 265203 272236 265269 272237
rect 265203 272172 265204 272236
rect 265268 272172 265269 272236
rect 265203 272171 265269 272172
rect 262075 270604 262141 270605
rect 262075 270540 262076 270604
rect 262140 270540 262141 270604
rect 262075 270539 262141 270540
rect 262811 270604 262877 270605
rect 262811 270540 262812 270604
rect 262876 270540 262877 270604
rect 262811 270539 262877 270540
rect 263915 270604 263981 270605
rect 263915 270540 263916 270604
rect 263980 270540 263981 270604
rect 263915 270539 263981 270540
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252308 261854 262338
rect 264954 266614 265574 272000
rect 265942 271557 266002 273670
rect 266381 273668 266382 273732
rect 266446 273668 266447 273732
rect 267608 273730 267668 274040
rect 266381 273667 266447 273668
rect 267598 273670 267668 273730
rect 268288 273730 268348 274040
rect 268696 273730 268756 274040
rect 269784 273730 269844 274040
rect 271008 273730 271068 274040
rect 268288 273670 268394 273730
rect 268696 273670 268762 273730
rect 269784 273670 269866 273730
rect 265939 271556 266005 271557
rect 265939 271492 265940 271556
rect 266004 271492 266005 271556
rect 265939 271491 266005 271492
rect 267598 270605 267658 273670
rect 268334 271557 268394 273670
rect 268702 271829 268762 273670
rect 268699 271828 268765 271829
rect 268699 271764 268700 271828
rect 268764 271764 268765 271828
rect 268699 271763 268765 271764
rect 268331 271556 268397 271557
rect 268331 271492 268332 271556
rect 268396 271492 268397 271556
rect 268331 271491 268397 271492
rect 269806 270605 269866 273670
rect 270910 273670 271068 273730
rect 271144 273730 271204 274040
rect 272232 273730 272292 274040
rect 271144 273670 271338 273730
rect 272232 273670 272626 273730
rect 270910 271829 270970 273670
rect 270907 271828 270973 271829
rect 270907 271764 270908 271828
rect 270972 271764 270973 271828
rect 270907 271763 270973 271764
rect 271278 270605 271338 273670
rect 267595 270604 267661 270605
rect 267595 270540 267596 270604
rect 267660 270540 267661 270604
rect 267595 270539 267661 270540
rect 269803 270604 269869 270605
rect 269803 270540 269804 270604
rect 269868 270540 269869 270604
rect 269803 270539 269869 270540
rect 271275 270604 271341 270605
rect 271275 270540 271276 270604
rect 271340 270540 271341 270604
rect 271275 270539 271341 270540
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252308 265574 266058
rect 271794 256394 272414 272000
rect 272566 271557 272626 273670
rect 273320 273597 273380 274040
rect 273592 273730 273652 274040
rect 274408 273730 274468 274040
rect 273486 273670 273652 273730
rect 274406 273670 274468 273730
rect 273317 273596 273383 273597
rect 273317 273532 273318 273596
rect 273382 273532 273383 273596
rect 273317 273531 273383 273532
rect 272563 271556 272629 271557
rect 272563 271492 272564 271556
rect 272628 271492 272629 271556
rect 272563 271491 272629 271492
rect 273486 271421 273546 273670
rect 273483 271420 273549 271421
rect 273483 271356 273484 271420
rect 273548 271356 273549 271420
rect 273483 271355 273549 271356
rect 274406 270605 274466 273670
rect 275768 273597 275828 274040
rect 276040 273730 276100 274040
rect 276992 273730 277052 274040
rect 278080 273733 278140 274040
rect 276040 273670 276306 273730
rect 275765 273596 275831 273597
rect 275765 273532 275766 273596
rect 275830 273532 275831 273596
rect 275765 273531 275831 273532
rect 274403 270604 274469 270605
rect 274403 270540 274404 270604
rect 274468 270540 274469 270604
rect 274403 270539 274469 270540
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 252308 272414 255838
rect 275514 260114 276134 272000
rect 276246 271829 276306 273670
rect 276982 273670 277052 273730
rect 278077 273732 278143 273733
rect 276243 271828 276309 271829
rect 276243 271764 276244 271828
rect 276308 271764 276309 271828
rect 276243 271763 276309 271764
rect 276982 271557 277042 273670
rect 278077 273668 278078 273732
rect 278142 273668 278143 273732
rect 278488 273730 278548 274040
rect 279168 273730 279228 274040
rect 280936 273730 280996 274040
rect 278077 273667 278143 273668
rect 278454 273670 278548 273730
rect 279006 273670 279228 273730
rect 280846 273670 280996 273730
rect 276979 271556 277045 271557
rect 276979 271492 276980 271556
rect 277044 271492 277045 271556
rect 276979 271491 277045 271492
rect 278454 271421 278514 273670
rect 278451 271420 278517 271421
rect 278451 271356 278452 271420
rect 278516 271356 278517 271420
rect 278451 271355 278517 271356
rect 279006 270877 279066 273670
rect 279003 270876 279069 270877
rect 279003 270812 279004 270876
rect 279068 270812 279069 270876
rect 279003 270811 279069 270812
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 252308 276134 259558
rect 279234 261954 279854 272000
rect 280846 271829 280906 273670
rect 283520 273597 283580 274040
rect 285968 273730 286028 274040
rect 288280 273730 288340 274040
rect 291000 273730 291060 274040
rect 293448 273730 293508 274040
rect 285968 273670 286058 273730
rect 283517 273596 283583 273597
rect 283517 273532 283518 273596
rect 283582 273532 283583 273596
rect 283517 273531 283583 273532
rect 285998 273325 286058 273670
rect 288206 273670 288340 273730
rect 290966 273670 291060 273730
rect 293358 273670 293508 273730
rect 295896 273730 295956 274040
rect 298480 273730 298540 274040
rect 300928 273730 300988 274040
rect 303512 273730 303572 274040
rect 305960 273730 306020 274040
rect 295896 273670 295994 273730
rect 298480 273670 298570 273730
rect 285995 273324 286061 273325
rect 285995 273260 285996 273324
rect 286060 273260 286061 273324
rect 285995 273259 286061 273260
rect 288206 272917 288266 273670
rect 290966 272917 291026 273670
rect 293358 272917 293418 273670
rect 288203 272916 288269 272917
rect 288203 272852 288204 272916
rect 288268 272852 288269 272916
rect 288203 272851 288269 272852
rect 290963 272916 291029 272917
rect 290963 272852 290964 272916
rect 291028 272852 291029 272916
rect 290963 272851 291029 272852
rect 293355 272916 293421 272917
rect 293355 272852 293356 272916
rect 293420 272852 293421 272916
rect 293355 272851 293421 272852
rect 295934 272645 295994 273670
rect 298510 272781 298570 273670
rect 300902 273670 300988 273730
rect 303478 273670 303572 273730
rect 305870 273670 306020 273730
rect 308544 273730 308604 274040
rect 310992 273730 311052 274040
rect 313440 273730 313500 274040
rect 315888 273730 315948 274040
rect 318472 273730 318532 274040
rect 308544 273670 308690 273730
rect 310992 273670 311082 273730
rect 300902 272917 300962 273670
rect 300899 272916 300965 272917
rect 300899 272852 300900 272916
rect 300964 272852 300965 272916
rect 300899 272851 300965 272852
rect 298507 272780 298573 272781
rect 298507 272716 298508 272780
rect 298572 272716 298573 272780
rect 298507 272715 298573 272716
rect 303478 272645 303538 273670
rect 305870 272645 305930 273670
rect 295931 272644 295997 272645
rect 295931 272580 295932 272644
rect 295996 272580 295997 272644
rect 295931 272579 295997 272580
rect 303475 272644 303541 272645
rect 303475 272580 303476 272644
rect 303540 272580 303541 272644
rect 303475 272579 303541 272580
rect 305867 272644 305933 272645
rect 305867 272580 305868 272644
rect 305932 272580 305933 272644
rect 305867 272579 305933 272580
rect 280843 271828 280909 271829
rect 280843 271764 280844 271828
rect 280908 271764 280909 271828
rect 280843 271763 280909 271764
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 252308 279854 261398
rect 282954 265674 283574 272000
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 252308 283574 265118
rect 289794 255454 290414 272000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252308 290414 254898
rect 293514 259174 294134 272000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252308 294134 258618
rect 297234 262894 297854 272000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252308 297854 262338
rect 300954 266614 301574 272000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252308 301574 266058
rect 307794 256394 308414 272000
rect 308630 271829 308690 273670
rect 311022 273053 311082 273670
rect 313414 273670 313500 273730
rect 315070 273670 315948 273730
rect 318382 273670 318532 273730
rect 320920 273730 320980 274040
rect 323368 273730 323428 274040
rect 325952 273730 326012 274040
rect 343224 273730 343284 274040
rect 320920 273670 321018 273730
rect 311019 273052 311085 273053
rect 311019 272988 311020 273052
rect 311084 272988 311085 273052
rect 311019 272987 311085 272988
rect 308627 271828 308693 271829
rect 308627 271764 308628 271828
rect 308692 271764 308693 271828
rect 308627 271763 308693 271764
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 252308 308414 255838
rect 311514 260114 312134 272000
rect 313414 271829 313474 273670
rect 313411 271828 313477 271829
rect 313411 271764 313412 271828
rect 313476 271764 313477 271828
rect 313411 271763 313477 271764
rect 315070 271693 315130 273670
rect 318382 273189 318442 273670
rect 318379 273188 318445 273189
rect 318379 273124 318380 273188
rect 318444 273124 318445 273188
rect 318379 273123 318445 273124
rect 320958 272645 321018 273670
rect 323350 273670 323428 273730
rect 325742 273670 326012 273730
rect 343222 273670 343284 273730
rect 343360 273730 343420 274040
rect 343360 273670 343466 273730
rect 320955 272644 321021 272645
rect 320955 272580 320956 272644
rect 321020 272580 321021 272644
rect 320955 272579 321021 272580
rect 315067 271692 315133 271693
rect 315067 271628 315068 271692
rect 315132 271628 315133 271692
rect 315067 271627 315133 271628
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 252308 312134 259558
rect 315234 261954 315854 272000
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 252308 315854 261398
rect 318954 265674 319574 272000
rect 323350 270469 323410 273670
rect 325742 272370 325802 273670
rect 325558 272310 325802 272370
rect 325558 271013 325618 272310
rect 325555 271012 325621 271013
rect 325555 270948 325556 271012
rect 325620 270948 325621 271012
rect 325555 270947 325621 270948
rect 323347 270468 323413 270469
rect 323347 270404 323348 270468
rect 323412 270404 323413 270468
rect 323347 270403 323413 270404
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 252308 319574 265118
rect 325794 255454 326414 272000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252308 326414 254898
rect 329514 259174 330134 272000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252308 330134 258618
rect 333234 262894 333854 272000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252308 333854 262338
rect 336954 266614 337574 272000
rect 343222 271557 343282 273670
rect 343406 271829 343466 273670
rect 343403 271828 343469 271829
rect 343403 271764 343404 271828
rect 343468 271764 343469 271828
rect 343403 271763 343469 271764
rect 343219 271556 343285 271557
rect 343219 271492 343220 271556
rect 343284 271492 343285 271556
rect 343219 271491 343285 271492
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252308 337574 266058
rect 343794 256394 344414 272000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 339723 253468 339789 253469
rect 339723 253404 339724 253468
rect 339788 253404 339789 253468
rect 339723 253403 339789 253404
rect 338435 253060 338501 253061
rect 338435 252996 338436 253060
rect 338500 252996 338501 253060
rect 338435 252995 338501 252996
rect 338438 250610 338498 252995
rect 339726 250610 339786 253403
rect 343794 252308 344414 255838
rect 347514 260114 348134 272000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 252308 348134 259558
rect 351234 261954 351854 272000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 350947 253196 351013 253197
rect 350947 253132 350948 253196
rect 351012 253132 351013 253196
rect 350947 253131 351013 253132
rect 350950 250610 351010 253131
rect 351234 252308 351854 261398
rect 354954 265674 355574 272000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 252308 355574 265118
rect 338438 250550 338524 250610
rect 338464 250240 338524 250550
rect 339688 250550 339786 250610
rect 350840 250550 351010 250610
rect 339688 250240 339748 250550
rect 350840 250240 350900 250550
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 166290 236116 167106
rect 237144 166290 237204 167106
rect 238232 166290 238292 167106
rect 235950 166230 236116 166290
rect 237054 166230 237204 166290
rect 238158 166230 238292 166290
rect 239592 166290 239652 167106
rect 240544 166290 240604 167106
rect 241768 166290 241828 167106
rect 243128 166290 243188 167106
rect 244216 167010 244276 167106
rect 245440 167010 245500 167106
rect 246528 167010 246588 167106
rect 247616 167010 247676 167106
rect 248296 167010 248356 167106
rect 248704 167010 248764 167106
rect 244216 166950 244474 167010
rect 244216 166910 244290 166950
rect 239592 166230 239690 166290
rect 240544 166230 240610 166290
rect 235950 165613 236010 166230
rect 235947 165612 236013 165613
rect 235947 165548 235948 165612
rect 236012 165548 236013 165612
rect 235947 165547 236013 165548
rect 221514 151174 222134 165000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 165000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 165000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 165000
rect 237054 164253 237114 166230
rect 238158 164253 238218 166230
rect 239630 165613 239690 166230
rect 239627 165612 239693 165613
rect 239627 165548 239628 165612
rect 239692 165548 239693 165612
rect 239627 165547 239693 165548
rect 237051 164252 237117 164253
rect 237051 164188 237052 164252
rect 237116 164188 237117 164252
rect 237051 164187 237117 164188
rect 238155 164252 238221 164253
rect 238155 164188 238156 164252
rect 238220 164188 238221 164252
rect 238155 164187 238221 164188
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 165000
rect 240550 164253 240610 166230
rect 241654 166230 241828 166290
rect 243126 166230 243188 166290
rect 241654 164253 241714 166230
rect 243126 165613 243186 166230
rect 243123 165612 243189 165613
rect 243123 165548 243124 165612
rect 243188 165548 243189 165612
rect 243123 165547 243189 165548
rect 240547 164252 240613 164253
rect 240547 164188 240548 164252
rect 240612 164188 240613 164252
rect 240547 164187 240613 164188
rect 241651 164252 241717 164253
rect 241651 164188 241652 164252
rect 241716 164188 241717 164252
rect 241651 164187 241717 164188
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 155834 243854 165000
rect 244414 164525 244474 166950
rect 245334 166950 245500 167010
rect 246438 166950 246588 167010
rect 247542 166950 247676 167010
rect 248278 166950 248356 167010
rect 248646 166950 248764 167010
rect 250064 167010 250124 167106
rect 250744 167010 250804 167106
rect 251288 167010 251348 167106
rect 252376 167010 252436 167106
rect 253464 167010 253524 167106
rect 250064 166950 250178 167010
rect 244411 164524 244477 164525
rect 244411 164460 244412 164524
rect 244476 164460 244477 164524
rect 244411 164459 244477 164460
rect 245334 164253 245394 166950
rect 246438 164253 246498 166950
rect 247542 165613 247602 166950
rect 248278 165613 248338 166950
rect 247539 165612 247605 165613
rect 247539 165548 247540 165612
rect 247604 165548 247605 165612
rect 247539 165547 247605 165548
rect 248275 165612 248341 165613
rect 248275 165548 248276 165612
rect 248340 165548 248341 165612
rect 248275 165547 248341 165548
rect 245331 164252 245397 164253
rect 245331 164188 245332 164252
rect 245396 164188 245397 164252
rect 245331 164187 245397 164188
rect 246435 164252 246501 164253
rect 246435 164188 246436 164252
rect 246500 164188 246501 164252
rect 246435 164187 246501 164188
rect 243234 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 243854 155834
rect 243234 155514 243854 155598
rect 243234 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 243854 155514
rect 243234 145308 243854 155278
rect 246954 157674 247574 165000
rect 248646 164253 248706 166950
rect 250118 164253 250178 166950
rect 250670 166950 250804 167010
rect 251222 166950 251348 167010
rect 252326 166950 252436 167010
rect 253430 166950 253524 167010
rect 253600 167010 253660 167106
rect 254552 167010 254612 167106
rect 255912 167010 255972 167106
rect 253600 166950 253674 167010
rect 250670 165613 250730 166950
rect 250667 165612 250733 165613
rect 250667 165548 250668 165612
rect 250732 165548 250733 165612
rect 250667 165547 250733 165548
rect 251222 164253 251282 166950
rect 252326 164525 252386 166950
rect 252323 164524 252389 164525
rect 252323 164460 252324 164524
rect 252388 164460 252389 164524
rect 252323 164459 252389 164460
rect 253430 164253 253490 166950
rect 253614 165613 253674 166950
rect 254534 166950 254612 167010
rect 255822 166950 255972 167010
rect 256048 167010 256108 167106
rect 257000 167010 257060 167106
rect 256048 166950 256250 167010
rect 253611 165612 253677 165613
rect 253611 165548 253612 165612
rect 253676 165548 253677 165612
rect 253611 165547 253677 165548
rect 248643 164252 248709 164253
rect 248643 164188 248644 164252
rect 248708 164188 248709 164252
rect 248643 164187 248709 164188
rect 250115 164252 250181 164253
rect 250115 164188 250116 164252
rect 250180 164188 250181 164252
rect 250115 164187 250181 164188
rect 251219 164252 251285 164253
rect 251219 164188 251220 164252
rect 251284 164188 251285 164252
rect 251219 164187 251285 164188
rect 253427 164252 253493 164253
rect 253427 164188 253428 164252
rect 253492 164188 253493 164252
rect 253427 164187 253493 164188
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 165000
rect 254534 164253 254594 166950
rect 255822 164253 255882 166950
rect 256190 164797 256250 166950
rect 256926 166950 257060 167010
rect 258088 167010 258148 167106
rect 258496 167010 258556 167106
rect 258088 166950 258274 167010
rect 256187 164796 256253 164797
rect 256187 164732 256188 164796
rect 256252 164732 256253 164796
rect 256187 164731 256253 164732
rect 256926 164253 256986 166950
rect 254531 164252 254597 164253
rect 254531 164188 254532 164252
rect 254596 164188 254597 164252
rect 254531 164187 254597 164188
rect 255819 164252 255885 164253
rect 255819 164188 255820 164252
rect 255884 164188 255885 164252
rect 255819 164187 255885 164188
rect 256923 164252 256989 164253
rect 256923 164188 256924 164252
rect 256988 164188 256989 164252
rect 256923 164187 256989 164188
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 165000
rect 258214 164250 258274 166950
rect 258398 166950 258556 167010
rect 259448 167010 259508 167106
rect 260672 167010 260732 167106
rect 261080 167010 261140 167106
rect 261760 167010 261820 167106
rect 262848 167010 262908 167106
rect 259448 166950 259562 167010
rect 258398 165613 258458 166950
rect 258395 165612 258461 165613
rect 258395 165548 258396 165612
rect 258460 165548 258461 165612
rect 258395 165547 258461 165548
rect 259502 164253 259562 166950
rect 260606 166950 260732 167010
rect 260974 166950 261140 167010
rect 261710 166950 261820 167010
rect 262814 166950 262908 167010
rect 263528 167010 263588 167106
rect 263936 167010 263996 167106
rect 265296 167010 265356 167106
rect 265976 167010 266036 167106
rect 263528 166950 263794 167010
rect 260606 164525 260666 166950
rect 260974 166565 261034 166950
rect 260971 166564 261037 166565
rect 260971 166500 260972 166564
rect 261036 166500 261037 166564
rect 260971 166499 261037 166500
rect 261710 165613 261770 166950
rect 261707 165612 261773 165613
rect 261707 165548 261708 165612
rect 261772 165548 261773 165612
rect 261707 165547 261773 165548
rect 260603 164524 260669 164525
rect 260603 164460 260604 164524
rect 260668 164460 260669 164524
rect 260603 164459 260669 164460
rect 258395 164252 258461 164253
rect 258395 164250 258396 164252
rect 258214 164190 258396 164250
rect 258395 164188 258396 164190
rect 258460 164188 258461 164252
rect 258395 164187 258461 164188
rect 259499 164252 259565 164253
rect 259499 164188 259500 164252
rect 259564 164188 259565 164252
rect 259499 164187 259565 164188
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 165000
rect 262814 164253 262874 166950
rect 263734 164933 263794 166950
rect 263918 166950 263996 167010
rect 265206 166950 265356 167010
rect 265942 166950 266036 167010
rect 266384 167010 266444 167106
rect 267608 167010 267668 167106
rect 266384 166950 266554 167010
rect 263731 164932 263797 164933
rect 263731 164868 263732 164932
rect 263796 164868 263797 164932
rect 263731 164867 263797 164868
rect 263918 164253 263978 166950
rect 265206 165613 265266 166950
rect 265942 166565 266002 166950
rect 265939 166564 266005 166565
rect 265939 166500 265940 166564
rect 266004 166500 266005 166564
rect 265939 166499 266005 166500
rect 266494 165613 266554 166950
rect 267598 166950 267668 167010
rect 268288 167010 268348 167106
rect 268696 167010 268756 167106
rect 269784 167010 269844 167106
rect 271008 167010 271068 167106
rect 268288 166950 268394 167010
rect 268696 166950 268762 167010
rect 269784 166950 269866 167010
rect 265203 165612 265269 165613
rect 265203 165548 265204 165612
rect 265268 165548 265269 165612
rect 265203 165547 265269 165548
rect 266491 165612 266557 165613
rect 266491 165548 266492 165612
rect 266556 165548 266557 165612
rect 266491 165547 266557 165548
rect 262811 164252 262877 164253
rect 262811 164188 262812 164252
rect 262876 164188 262877 164252
rect 262811 164187 262877 164188
rect 263915 164252 263981 164253
rect 263915 164188 263916 164252
rect 263980 164188 263981 164252
rect 263915 164187 263981 164188
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 165000
rect 267598 164525 267658 166950
rect 268334 165613 268394 166950
rect 268331 165612 268397 165613
rect 268331 165548 268332 165612
rect 268396 165548 268397 165612
rect 268331 165547 268397 165548
rect 267595 164524 267661 164525
rect 267595 164460 267596 164524
rect 267660 164460 267661 164524
rect 267595 164459 267661 164460
rect 268702 164253 268762 166950
rect 269806 164253 269866 166950
rect 270910 166950 271068 167010
rect 271144 167010 271204 167106
rect 272232 167010 272292 167106
rect 273320 167010 273380 167106
rect 273592 167010 273652 167106
rect 274408 167010 274468 167106
rect 271144 166950 271338 167010
rect 270910 166565 270970 166950
rect 270907 166564 270973 166565
rect 270907 166500 270908 166564
rect 270972 166500 270973 166564
rect 270907 166499 270973 166500
rect 271278 164253 271338 166950
rect 272198 166950 272292 167010
rect 273302 166950 273380 167010
rect 273486 166950 273652 167010
rect 274406 166950 274468 167010
rect 275768 167010 275828 167106
rect 276040 167010 276100 167106
rect 276992 167010 277052 167106
rect 275768 166950 275938 167010
rect 276040 166950 276122 167010
rect 272198 165205 272258 166950
rect 272195 165204 272261 165205
rect 272195 165140 272196 165204
rect 272260 165140 272261 165204
rect 272195 165139 272261 165140
rect 268699 164252 268765 164253
rect 268699 164188 268700 164252
rect 268764 164188 268765 164252
rect 268699 164187 268765 164188
rect 269803 164252 269869 164253
rect 269803 164188 269804 164252
rect 269868 164188 269869 164252
rect 269803 164187 269869 164188
rect 271275 164252 271341 164253
rect 271275 164188 271276 164252
rect 271340 164188 271341 164252
rect 271275 164187 271341 164188
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 165000
rect 273302 164525 273362 166950
rect 273486 165069 273546 166950
rect 273483 165068 273549 165069
rect 273483 165004 273484 165068
rect 273548 165004 273549 165068
rect 273483 165003 273549 165004
rect 273299 164524 273365 164525
rect 273299 164460 273300 164524
rect 273364 164460 273365 164524
rect 273299 164459 273365 164460
rect 274406 164253 274466 166950
rect 275878 165205 275938 166950
rect 276062 165205 276122 166950
rect 276982 166950 277052 167010
rect 278080 167010 278140 167106
rect 278488 167010 278548 167106
rect 278080 166950 278146 167010
rect 275875 165204 275941 165205
rect 275875 165140 275876 165204
rect 275940 165140 275941 165204
rect 275875 165139 275941 165140
rect 276059 165204 276125 165205
rect 276059 165140 276060 165204
rect 276124 165140 276125 165204
rect 276059 165139 276125 165140
rect 274403 164252 274469 164253
rect 274403 164188 274404 164252
rect 274468 164188 274469 164252
rect 274403 164187 274469 164188
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 165000
rect 276982 164253 277042 166950
rect 278086 164253 278146 166950
rect 278454 166950 278548 167010
rect 279168 167010 279228 167106
rect 280936 167010 280996 167106
rect 279168 166950 279250 167010
rect 278454 165205 278514 166950
rect 279190 165205 279250 166950
rect 280846 166950 280996 167010
rect 280846 165613 280906 166950
rect 283520 166290 283580 167106
rect 285968 166701 286028 167106
rect 285965 166700 286031 166701
rect 285965 166636 285966 166700
rect 286030 166636 286031 166700
rect 285965 166635 286031 166636
rect 288280 166565 288340 167106
rect 291000 166701 291060 167106
rect 293448 166701 293508 167106
rect 295896 166701 295956 167106
rect 298480 166701 298540 167106
rect 290997 166700 291063 166701
rect 290997 166636 290998 166700
rect 291062 166636 291063 166700
rect 290997 166635 291063 166636
rect 293445 166700 293511 166701
rect 293445 166636 293446 166700
rect 293510 166636 293511 166700
rect 293445 166635 293511 166636
rect 295893 166700 295959 166701
rect 295893 166636 295894 166700
rect 295958 166636 295959 166700
rect 295893 166635 295959 166636
rect 298477 166700 298543 166701
rect 298477 166636 298478 166700
rect 298542 166636 298543 166700
rect 298477 166635 298543 166636
rect 288277 166564 288343 166565
rect 288277 166500 288278 166564
rect 288342 166500 288343 166564
rect 288277 166499 288343 166500
rect 300928 166290 300988 167106
rect 303512 166837 303572 167106
rect 303509 166836 303575 166837
rect 303509 166772 303510 166836
rect 303574 166772 303575 166836
rect 303509 166771 303575 166772
rect 305960 166701 306020 167106
rect 305957 166700 306023 166701
rect 305957 166636 305958 166700
rect 306022 166636 306023 166700
rect 308544 166698 308604 167106
rect 305957 166635 306023 166636
rect 308446 166638 308604 166698
rect 310992 166698 311052 167106
rect 313440 166837 313500 167106
rect 313437 166836 313503 166837
rect 313437 166772 313438 166836
rect 313502 166772 313503 166836
rect 313437 166771 313503 166772
rect 315888 166698 315948 167106
rect 318472 166698 318532 167106
rect 310992 166638 311082 166698
rect 283422 166230 283580 166290
rect 300902 166230 300988 166290
rect 283422 165613 283482 166230
rect 300902 165613 300962 166230
rect 308446 165613 308506 166638
rect 280843 165612 280909 165613
rect 280843 165548 280844 165612
rect 280908 165548 280909 165612
rect 280843 165547 280909 165548
rect 283419 165612 283485 165613
rect 283419 165548 283420 165612
rect 283484 165548 283485 165612
rect 283419 165547 283485 165548
rect 300899 165612 300965 165613
rect 300899 165548 300900 165612
rect 300964 165548 300965 165612
rect 300899 165547 300965 165548
rect 308443 165612 308509 165613
rect 308443 165548 308444 165612
rect 308508 165548 308509 165612
rect 308443 165547 308509 165548
rect 311022 165341 311082 166638
rect 315070 166638 315948 166698
rect 318382 166638 318532 166698
rect 320920 166698 320980 167106
rect 323368 166698 323428 167106
rect 320920 166638 321018 166698
rect 311019 165340 311085 165341
rect 311019 165276 311020 165340
rect 311084 165276 311085 165340
rect 311019 165275 311085 165276
rect 278451 165204 278517 165205
rect 278451 165140 278452 165204
rect 278516 165140 278517 165204
rect 278451 165139 278517 165140
rect 279187 165204 279253 165205
rect 279187 165140 279188 165204
rect 279252 165140 279253 165204
rect 279187 165139 279253 165140
rect 276979 164252 277045 164253
rect 276979 164188 276980 164252
rect 277044 164188 277045 164252
rect 276979 164187 277045 164188
rect 278083 164252 278149 164253
rect 278083 164188 278084 164252
rect 278148 164188 278149 164252
rect 278083 164187 278149 164188
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 155834 279854 165000
rect 279234 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 279854 155834
rect 279234 155514 279854 155598
rect 279234 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 279854 155514
rect 279234 145308 279854 155278
rect 282954 157674 283574 165000
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 165000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 165000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 165000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 165000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 165000
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 165000
rect 315070 164389 315130 166638
rect 315067 164388 315133 164389
rect 315067 164324 315068 164388
rect 315132 164324 315133 164388
rect 315067 164323 315133 164324
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 155834 315854 165000
rect 318382 164253 318442 166638
rect 320958 165477 321018 166638
rect 323350 166638 323428 166698
rect 323350 165613 323410 166638
rect 325952 166290 326012 167106
rect 343224 166290 343284 167106
rect 325926 166230 326012 166290
rect 343222 166230 343284 166290
rect 343360 166290 343420 167106
rect 343360 166230 343466 166290
rect 325926 165613 325986 166230
rect 343222 165613 343282 166230
rect 343406 165613 343466 166230
rect 323347 165612 323413 165613
rect 323347 165548 323348 165612
rect 323412 165548 323413 165612
rect 323347 165547 323413 165548
rect 325923 165612 325989 165613
rect 325923 165548 325924 165612
rect 325988 165548 325989 165612
rect 325923 165547 325989 165548
rect 343219 165612 343285 165613
rect 343219 165548 343220 165612
rect 343284 165548 343285 165612
rect 343219 165547 343285 165548
rect 343403 165612 343469 165613
rect 343403 165548 343404 165612
rect 343468 165548 343469 165612
rect 343403 165547 343469 165548
rect 320955 165476 321021 165477
rect 320955 165412 320956 165476
rect 321020 165412 321021 165476
rect 320955 165411 321021 165412
rect 318379 164252 318445 164253
rect 318379 164188 318380 164252
rect 318444 164188 318445 164252
rect 318379 164187 318445 164188
rect 315234 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 315854 155834
rect 315234 155514 315854 155598
rect 315234 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 315854 155514
rect 315234 145308 315854 155278
rect 318954 157674 319574 165000
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 165000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 165000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 165000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 165000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 165000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 165000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 155834 351854 165000
rect 351234 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 351854 155834
rect 351234 155514 351854 155598
rect 351234 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 351854 155514
rect 351234 145308 351854 155278
rect 354954 157674 355574 165000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59530 236116 60106
rect 237144 59805 237204 60106
rect 237141 59804 237207 59805
rect 237141 59740 237142 59804
rect 237206 59740 237207 59804
rect 237141 59739 237207 59740
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 235950 59470 236116 59530
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 235950 58173 236010 59470
rect 235947 58172 236013 58173
rect 235947 58108 235948 58172
rect 236012 58108 236013 58172
rect 235947 58107 236013 58108
rect 219939 56540 220005 56541
rect 219939 56476 219940 56540
rect 220004 56476 220005 56540
rect 219939 56475 220005 56476
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57901 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57901 241714 59470
rect 242942 57901 243002 59470
rect 240547 57900 240613 57901
rect 240547 57836 240548 57900
rect 240612 57836 240613 57900
rect 240547 57835 240613 57836
rect 241651 57900 241717 57901
rect 241651 57836 241652 57900
rect 241716 57836 241717 57900
rect 241651 57835 241717 57836
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57901 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 244227 57900 244293 57901
rect 244227 57836 244228 57900
rect 244292 57836 244293 57900
rect 244227 57835 244293 57836
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57901 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59666 250804 60106
rect 251288 59666 251348 60106
rect 250670 59606 250804 59666
rect 251222 59606 251348 59666
rect 250064 59470 250178 59530
rect 247723 57900 247789 57901
rect 247723 57836 247724 57900
rect 247788 57836 247789 57900
rect 247723 57835 247789 57836
rect 248278 57085 248338 59470
rect 248646 57901 248706 59470
rect 250118 57901 250178 59470
rect 250670 58581 250730 59606
rect 250667 58580 250733 58581
rect 250667 58516 250668 58580
rect 250732 58516 250733 58580
rect 250667 58515 250733 58516
rect 251222 57901 251282 59606
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59805 257060 60106
rect 256997 59804 257063 59805
rect 256997 59740 256998 59804
rect 257062 59740 257063 59804
rect 256997 59739 257063 59740
rect 258088 59669 258148 60106
rect 258085 59668 258151 59669
rect 258085 59604 258086 59668
rect 258150 59604 258151 59668
rect 258085 59603 258151 59604
rect 258496 59530 258556 60106
rect 253600 59470 253674 59530
rect 252326 57901 252386 59470
rect 253430 57901 253490 59470
rect 253614 58717 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 258398 59470 258556 59530
rect 259448 59530 259508 60106
rect 260672 59669 260732 60106
rect 260669 59668 260735 59669
rect 260669 59604 260670 59668
rect 260734 59604 260735 59668
rect 260669 59603 260735 59604
rect 261080 59530 261140 60106
rect 261760 59669 261820 60106
rect 262848 59805 262908 60106
rect 262845 59804 262911 59805
rect 262845 59740 262846 59804
rect 262910 59740 262911 59804
rect 262845 59739 262911 59740
rect 261757 59668 261823 59669
rect 261757 59604 261758 59668
rect 261822 59604 261823 59668
rect 261757 59603 261823 59604
rect 259448 59470 259562 59530
rect 253611 58716 253677 58717
rect 253611 58652 253612 58716
rect 253676 58652 253677 58716
rect 253611 58651 253677 58652
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250115 57900 250181 57901
rect 250115 57836 250116 57900
rect 250180 57836 250181 57900
rect 250115 57835 250181 57836
rect 251219 57900 251285 57901
rect 251219 57836 251220 57900
rect 251284 57836 251285 57900
rect 251219 57835 251285 57836
rect 252323 57900 252389 57901
rect 252323 57836 252324 57900
rect 252388 57836 252389 57900
rect 252323 57835 252389 57836
rect 253427 57900 253493 57901
rect 253427 57836 253428 57900
rect 253492 57836 253493 57900
rect 253427 57835 253493 57836
rect 248275 57084 248341 57085
rect 248275 57020 248276 57084
rect 248340 57020 248341 57084
rect 248275 57019 248341 57020
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57901 254594 59470
rect 254531 57900 254597 57901
rect 254531 57836 254532 57900
rect 254596 57836 254597 57900
rect 254531 57835 254597 57836
rect 256006 57357 256066 59470
rect 256003 57356 256069 57357
rect 256003 57292 256004 57356
rect 256068 57292 256069 57356
rect 256003 57291 256069 57292
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 258398 57901 258458 59470
rect 259502 58445 259562 59470
rect 260974 59470 261140 59530
rect 263528 59530 263588 60106
rect 263936 59805 263996 60106
rect 263933 59804 263999 59805
rect 263933 59740 263934 59804
rect 263998 59740 263999 59804
rect 263933 59739 263999 59740
rect 265296 59530 265356 60106
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263528 59470 263610 59530
rect 259499 58444 259565 58445
rect 259499 58380 259500 58444
rect 259564 58380 259565 58444
rect 259499 58379 259565 58380
rect 258395 57900 258461 57901
rect 258395 57836 258396 57900
rect 258460 57836 258461 57900
rect 258395 57835 258461 57836
rect 260974 57493 261034 59470
rect 263550 59397 263610 59470
rect 265206 59470 265356 59530
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59666 271068 60106
rect 270910 59606 271068 59666
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 263547 59396 263613 59397
rect 263547 59332 263548 59396
rect 263612 59332 263613 59396
rect 263547 59331 263613 59332
rect 265206 58173 265266 59470
rect 265203 58172 265269 58173
rect 265203 58108 265204 58172
rect 265268 58108 265269 58172
rect 265203 58107 265269 58108
rect 260971 57492 261037 57493
rect 260971 57428 260972 57492
rect 261036 57428 261037 57492
rect 260971 57427 261037 57428
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57221 266002 59470
rect 266310 57901 266370 59470
rect 266307 57900 266373 57901
rect 266307 57836 266308 57900
rect 266372 57836 266373 57900
rect 266307 57835 266373 57836
rect 267598 57629 267658 59470
rect 268334 58989 268394 59470
rect 268331 58988 268397 58989
rect 268331 58924 268332 58988
rect 268396 58924 268397 58988
rect 268331 58923 268397 58924
rect 268702 57901 268762 59470
rect 268699 57900 268765 57901
rect 268699 57836 268700 57900
rect 268764 57836 268765 57900
rect 268699 57835 268765 57836
rect 269806 57629 269866 59470
rect 267595 57628 267661 57629
rect 267595 57564 267596 57628
rect 267660 57564 267661 57628
rect 267595 57563 267661 57564
rect 269803 57628 269869 57629
rect 269803 57564 269804 57628
rect 269868 57564 269869 57628
rect 269803 57563 269869 57564
rect 270910 57493 270970 59606
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59666 273652 60106
rect 271094 59470 271204 59530
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59606 273652 59666
rect 271094 57901 271154 59470
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 271091 57900 271157 57901
rect 271091 57836 271092 57900
rect 271156 57836 271157 57900
rect 271091 57835 271157 57836
rect 270907 57492 270973 57493
rect 270907 57428 270908 57492
rect 270972 57428 270973 57492
rect 270907 57427 270973 57428
rect 271794 57454 272414 58000
rect 273302 57901 273362 59470
rect 273299 57900 273365 57901
rect 273299 57836 273300 57900
rect 273364 57836 273365 57900
rect 273299 57835 273365 57836
rect 265939 57220 266005 57221
rect 265939 57156 265940 57220
rect 266004 57156 266005 57220
rect 265939 57155 266005 57156
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 273486 56405 273546 59606
rect 274408 59530 274468 60106
rect 275768 59666 275828 60106
rect 274406 59470 274468 59530
rect 275694 59606 275828 59666
rect 274406 57629 274466 59470
rect 275694 58173 275754 59606
rect 276040 59530 276100 60106
rect 276992 59530 277052 60106
rect 276040 59470 276122 59530
rect 276062 58853 276122 59470
rect 276982 59470 277052 59530
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 278080 59470 278146 59530
rect 276059 58852 276125 58853
rect 276059 58788 276060 58852
rect 276124 58788 276125 58852
rect 276059 58787 276125 58788
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57628 274469 57629
rect 274403 57564 274404 57628
rect 274468 57564 274469 57628
rect 274403 57563 274469 57564
rect 273483 56404 273549 56405
rect 273483 56340 273484 56404
rect 273548 56340 273549 56404
rect 273483 56339 273549 56340
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 56269 277042 59470
rect 278086 57629 278146 59470
rect 278454 59470 278548 59530
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 279168 59470 279250 59530
rect 278454 57765 278514 59470
rect 279190 59261 279250 59470
rect 280846 59470 280996 59530
rect 283520 59530 283580 60106
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 283520 59470 283850 59530
rect 285968 59470 286058 59530
rect 279187 59260 279253 59261
rect 279187 59196 279188 59260
rect 279252 59196 279253 59260
rect 279187 59195 279253 59196
rect 280846 59125 280906 59470
rect 280843 59124 280909 59125
rect 280843 59060 280844 59124
rect 280908 59060 280909 59124
rect 280843 59059 280909 59060
rect 278451 57764 278517 57765
rect 278451 57700 278452 57764
rect 278516 57700 278517 57764
rect 278451 57699 278517 57700
rect 278083 57628 278149 57629
rect 278083 57564 278084 57628
rect 278148 57564 278149 57628
rect 278083 57563 278149 57564
rect 276979 56268 277045 56269
rect 276979 56204 276980 56268
rect 277044 56204 277045 56268
rect 276979 56203 277045 56204
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 283790 57901 283850 59470
rect 285998 59261 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59530 306020 60106
rect 308544 59669 308604 60106
rect 308541 59668 308607 59669
rect 308541 59604 308542 59668
rect 308606 59604 308607 59668
rect 308541 59603 308607 59604
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 285995 59260 286061 59261
rect 285995 59196 285996 59260
rect 286060 59196 286061 59260
rect 285995 59195 286061 59196
rect 283787 57900 283853 57901
rect 283787 57836 283788 57900
rect 283852 57836 283853 57900
rect 283787 57835 283853 57836
rect 288206 56677 288266 59470
rect 290966 59261 291026 59470
rect 290963 59260 291029 59261
rect 290963 59196 290964 59260
rect 291028 59196 291029 59260
rect 290963 59195 291029 59196
rect 288203 56676 288269 56677
rect 288203 56612 288204 56676
rect 288268 56612 288269 56676
rect 288203 56611 288269 56612
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 57901 293418 59470
rect 293355 57900 293421 57901
rect 293355 57836 293356 57900
rect 293420 57836 293421 57900
rect 293355 57835 293421 57836
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 295934 57901 295994 59470
rect 295931 57900 295997 57901
rect 295931 57836 295932 57900
rect 295996 57836 295997 57900
rect 295931 57835 295997 57836
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 298510 57901 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 305870 59470 306020 59530
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59669 315948 60106
rect 315885 59668 315951 59669
rect 315885 59604 315886 59668
rect 315950 59604 315951 59668
rect 318472 59666 318532 60106
rect 315885 59603 315951 59604
rect 318382 59606 318532 59666
rect 310992 59470 311082 59530
rect 300902 59261 300962 59470
rect 300899 59260 300965 59261
rect 300899 59196 300900 59260
rect 300964 59196 300965 59260
rect 300899 59195 300965 59196
rect 298507 57900 298573 57901
rect 298507 57836 298508 57900
rect 298572 57836 298573 57900
rect 298507 57835 298573 57836
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 303478 57901 303538 59470
rect 305870 57901 305930 59470
rect 303475 57900 303541 57901
rect 303475 57836 303476 57900
rect 303540 57836 303541 57900
rect 303475 57835 303541 57836
rect 305867 57900 305933 57901
rect 305867 57836 305868 57900
rect 305932 57836 305933 57900
rect 305867 57835 305933 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 313414 57901 313474 59470
rect 313411 57900 313477 57901
rect 313411 57836 313412 57900
rect 313476 57836 313477 57900
rect 313411 57835 313477 57836
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 318382 57901 318442 59606
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 320958 59261 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 320955 59260 321021 59261
rect 320955 59196 320956 59260
rect 321020 59196 321021 59260
rect 320955 59195 321021 59196
rect 318379 57900 318445 57901
rect 318379 57836 318380 57900
rect 318444 57836 318445 57900
rect 318379 57835 318445 57836
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 323350 57901 323410 59470
rect 325926 59261 325986 59470
rect 325923 59260 325989 59261
rect 325923 59196 325924 59260
rect 325988 59196 325989 59260
rect 325923 59195 325989 59196
rect 323347 57900 323413 57901
rect 323347 57836 323348 57900
rect 323412 57836 323413 57900
rect 323347 57835 323413 57836
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 357942 57629 358002 476851
rect 359414 273325 359474 479707
rect 359595 468484 359661 468485
rect 359595 468420 359596 468484
rect 359660 468420 359661 468484
rect 359595 468419 359661 468420
rect 359411 273324 359477 273325
rect 359411 273260 359412 273324
rect 359476 273260 359477 273324
rect 359411 273259 359477 273260
rect 359598 273189 359658 468419
rect 359782 378045 359842 482563
rect 359963 465764 360029 465765
rect 359963 465700 359964 465764
rect 360028 465700 360029 465764
rect 359963 465699 360029 465700
rect 359779 378044 359845 378045
rect 359779 377980 359780 378044
rect 359844 377980 359845 378044
rect 359779 377979 359845 377980
rect 359966 374645 360026 465699
rect 359963 374644 360029 374645
rect 359963 374580 359964 374644
rect 360028 374580 360029 374644
rect 359963 374579 360029 374580
rect 359595 273188 359661 273189
rect 359595 273124 359596 273188
rect 359660 273124 359661 273188
rect 359595 273123 359661 273124
rect 360702 59261 360762 484875
rect 360886 149157 360946 489091
rect 361794 471454 362414 506898
rect 365514 511174 366134 526000
rect 368243 518124 368309 518125
rect 368243 518060 368244 518124
rect 368308 518060 368309 518124
rect 368243 518059 368309 518060
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 364931 487796 364997 487797
rect 364931 487732 364932 487796
rect 364996 487732 364997 487796
rect 364931 487731 364997 487732
rect 363459 486436 363525 486437
rect 363459 486372 363460 486436
rect 363524 486372 363525 486436
rect 363459 486371 363525 486372
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360883 149156 360949 149157
rect 360883 149092 360884 149156
rect 360948 149092 360949 149156
rect 360883 149091 360949 149092
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 360699 59260 360765 59261
rect 360699 59196 360700 59260
rect 360764 59196 360765 59260
rect 360699 59195 360765 59196
rect 357939 57628 358005 57629
rect 357939 57564 357940 57628
rect 358004 57564 358005 57628
rect 357939 57563 358005 57564
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 363462 3637 363522 486371
rect 364934 3773 364994 487731
rect 365514 475174 366134 510618
rect 366219 485756 366285 485757
rect 366219 485692 366220 485756
rect 366284 485692 366285 485756
rect 366219 485691 366285 485692
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365115 472564 365181 472565
rect 365115 472500 365116 472564
rect 365180 472500 365181 472564
rect 365115 472499 365181 472500
rect 364931 3772 364997 3773
rect 364931 3708 364932 3772
rect 364996 3708 364997 3772
rect 364931 3707 364997 3708
rect 363459 3636 363525 3637
rect 363459 3572 363460 3636
rect 363524 3572 363525 3636
rect 363459 3571 363525 3572
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 365118 3365 365178 472499
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 366222 58989 366282 485691
rect 367691 475828 367757 475829
rect 367691 475764 367692 475828
rect 367756 475764 367757 475828
rect 367691 475763 367757 475764
rect 366219 58988 366285 58989
rect 366219 58924 366220 58988
rect 366284 58924 366285 58988
rect 366219 58923 366285 58924
rect 367694 56677 367754 475763
rect 367691 56676 367757 56677
rect 367691 56612 367692 56676
rect 367756 56612 367757 56676
rect 367691 56611 367757 56612
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365115 3364 365181 3365
rect 365115 3300 365116 3364
rect 365180 3300 365181 3364
rect 365115 3299 365181 3300
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 6618
rect 368246 2957 368306 518059
rect 369234 514894 369854 526000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 372954 518614 373574 526000
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 371923 485620 371989 485621
rect 371923 485556 371924 485620
rect 371988 485556 371989 485620
rect 371923 485555 371989 485556
rect 371739 485484 371805 485485
rect 371739 485420 371740 485484
rect 371804 485420 371805 485484
rect 371739 485419 371805 485420
rect 370451 485348 370517 485349
rect 370451 485284 370452 485348
rect 370516 485284 370517 485348
rect 370451 485283 370517 485284
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 370454 58581 370514 485283
rect 371742 58717 371802 485419
rect 371926 59125 371986 485555
rect 372954 482614 373574 518058
rect 379794 525454 380414 526000
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 373763 485212 373829 485213
rect 373763 485148 373764 485212
rect 373828 485148 373829 485212
rect 373763 485147 373829 485148
rect 375971 485212 376037 485213
rect 375971 485148 375972 485212
rect 376036 485148 376037 485212
rect 375971 485147 376037 485148
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 371923 59124 371989 59125
rect 371923 59060 371924 59124
rect 371988 59060 371989 59124
rect 371923 59059 371989 59060
rect 371739 58716 371805 58717
rect 371739 58652 371740 58716
rect 371804 58652 371805 58716
rect 371739 58651 371805 58652
rect 370451 58580 370517 58581
rect 370451 58516 370452 58580
rect 370516 58516 370517 58580
rect 370451 58515 370517 58516
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 368243 2956 368309 2957
rect 368243 2892 368244 2956
rect 368308 2892 368309 2956
rect 368243 2891 368309 2892
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 86058
rect 373766 58853 373826 485147
rect 375419 482492 375485 482493
rect 375419 482428 375420 482492
rect 375484 482428 375485 482492
rect 375419 482427 375485 482428
rect 374683 482356 374749 482357
rect 374683 482292 374684 482356
rect 374748 482292 374749 482356
rect 374683 482291 374749 482292
rect 374499 479636 374565 479637
rect 374499 479572 374500 479636
rect 374564 479572 374565 479636
rect 374499 479571 374565 479572
rect 373763 58852 373829 58853
rect 373763 58788 373764 58852
rect 373828 58788 373829 58852
rect 373763 58787 373829 58788
rect 374502 57357 374562 479571
rect 374686 68101 374746 482291
rect 374867 480996 374933 480997
rect 374867 480932 374868 480996
rect 374932 480932 374933 480996
rect 374867 480931 374933 480932
rect 374870 165205 374930 480931
rect 375422 269109 375482 482427
rect 375419 269108 375485 269109
rect 375419 269044 375420 269108
rect 375484 269044 375485 269108
rect 375419 269043 375485 269044
rect 374867 165204 374933 165205
rect 374867 165140 374868 165204
rect 374932 165140 374933 165204
rect 374867 165139 374933 165140
rect 374683 68100 374749 68101
rect 374683 68036 374684 68100
rect 374748 68036 374749 68100
rect 374683 68035 374749 68036
rect 374499 57356 374565 57357
rect 374499 57292 374500 57356
rect 374564 57292 374565 57356
rect 374499 57291 374565 57292
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 375974 3501 376034 485147
rect 376155 485076 376221 485077
rect 376155 485012 376156 485076
rect 376220 485012 376221 485076
rect 376155 485011 376221 485012
rect 376158 58445 376218 485011
rect 377259 481132 377325 481133
rect 377259 481068 377260 481132
rect 377324 481068 377325 481132
rect 377259 481067 377325 481068
rect 376891 475964 376957 475965
rect 376891 475900 376892 475964
rect 376956 475900 376957 475964
rect 376891 475899 376957 475900
rect 376894 381037 376954 475899
rect 376891 381036 376957 381037
rect 376891 380972 376892 381036
rect 376956 380972 376957 381036
rect 376891 380971 376957 380972
rect 376891 379540 376957 379541
rect 376891 379476 376892 379540
rect 376956 379476 376957 379540
rect 376891 379475 376957 379476
rect 376894 274685 376954 379475
rect 377262 376685 377322 481067
rect 378731 480860 378797 480861
rect 378731 480796 378732 480860
rect 378796 480796 378797 480860
rect 378731 480795 378797 480796
rect 377443 478548 377509 478549
rect 377443 478484 377444 478548
rect 377508 478484 377509 478548
rect 377443 478483 377509 478484
rect 377446 379405 377506 478483
rect 377627 471204 377693 471205
rect 377627 471140 377628 471204
rect 377692 471140 377693 471204
rect 377627 471139 377693 471140
rect 377443 379404 377509 379405
rect 377443 379340 377444 379404
rect 377508 379340 377509 379404
rect 377443 379339 377509 379340
rect 377630 378725 377690 471139
rect 377627 378724 377693 378725
rect 377627 378660 377628 378724
rect 377692 378660 377693 378724
rect 377627 378659 377693 378660
rect 377995 378180 378061 378181
rect 377995 378116 377996 378180
rect 378060 378116 378061 378180
rect 377995 378115 378061 378116
rect 377259 376684 377325 376685
rect 377259 376620 377260 376684
rect 377324 376620 377325 376684
rect 377259 376619 377325 376620
rect 377998 277410 378058 378115
rect 377814 277350 378058 277410
rect 376891 274684 376957 274685
rect 376891 274620 376892 274684
rect 376956 274620 376957 274684
rect 376891 274619 376957 274620
rect 376894 273461 376954 274619
rect 376891 273460 376957 273461
rect 376891 273396 376892 273460
rect 376956 273396 376957 273460
rect 376891 273395 376957 273396
rect 377814 271421 377874 277350
rect 377811 271420 377877 271421
rect 377811 271356 377812 271420
rect 377876 271356 377877 271420
rect 377811 271355 377877 271356
rect 377995 251836 378061 251837
rect 377995 251772 377996 251836
rect 378060 251772 378061 251836
rect 377995 251771 378061 251772
rect 377259 163028 377325 163029
rect 377259 162964 377260 163028
rect 377324 162964 377325 163028
rect 377259 162963 377325 162964
rect 376155 58444 376221 58445
rect 376155 58380 376156 58444
rect 376220 58380 376221 58444
rect 376155 58379 376221 58380
rect 377262 56405 377322 162963
rect 377998 146301 378058 251771
rect 377995 146300 378061 146301
rect 377995 146236 377996 146300
rect 378060 146236 378061 146300
rect 377995 146235 378061 146236
rect 377627 146164 377693 146165
rect 377627 146100 377628 146164
rect 377692 146100 377693 146164
rect 377627 146099 377693 146100
rect 377259 56404 377325 56405
rect 377259 56340 377260 56404
rect 377324 56340 377325 56404
rect 377259 56339 377325 56340
rect 377630 55045 377690 146099
rect 377811 144124 377877 144125
rect 377811 144060 377812 144124
rect 377876 144060 377877 144124
rect 377811 144059 377877 144060
rect 377814 55181 377874 144059
rect 378734 57765 378794 480795
rect 378915 478276 378981 478277
rect 378915 478212 378916 478276
rect 378980 478212 378981 478276
rect 378915 478211 378981 478212
rect 378731 57764 378797 57765
rect 378731 57700 378732 57764
rect 378796 57700 378797 57764
rect 378731 57699 378797 57700
rect 378918 57085 378978 478211
rect 379099 476780 379165 476781
rect 379099 476716 379100 476780
rect 379164 476716 379165 476780
rect 379099 476715 379165 476716
rect 379102 57493 379162 476715
rect 379467 475692 379533 475693
rect 379467 475628 379468 475692
rect 379532 475690 379533 475692
rect 379532 475630 379714 475690
rect 379532 475628 379533 475630
rect 379467 475627 379533 475628
rect 379283 475556 379349 475557
rect 379283 475492 379284 475556
rect 379348 475492 379349 475556
rect 379283 475491 379349 475492
rect 379099 57492 379165 57493
rect 379099 57428 379100 57492
rect 379164 57428 379165 57492
rect 379099 57427 379165 57428
rect 379286 57221 379346 475491
rect 379654 171150 379714 475630
rect 379794 466308 380414 488898
rect 383514 493174 384134 526000
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 466308 384134 492618
rect 387234 496894 387854 526000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 466308 387854 496338
rect 390954 500614 391574 526000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 466308 391574 500058
rect 397794 507454 398414 526000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 466308 398414 470898
rect 401514 511174 402134 526000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 466308 402134 474618
rect 405234 514894 405854 526000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 466308 405854 478338
rect 408954 518614 409574 526000
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 466308 409574 482058
rect 415794 525454 416414 526000
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 466308 416414 488898
rect 419514 493174 420134 526000
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 466308 420134 492618
rect 423234 496894 423854 526000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 466308 423854 496338
rect 426954 500614 427574 526000
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 466308 427574 500058
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 466308 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 466308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 466308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 466308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 466308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 630000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 630000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 630000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 630000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 630000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 630000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 630000 488414 632898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 630000 492134 636618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 630000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 630000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 630000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 630000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 476067 627876 476133 627877
rect 476067 627812 476068 627876
rect 476132 627812 476133 627876
rect 476067 627811 476133 627812
rect 488579 627876 488645 627877
rect 488579 627812 488580 627876
rect 488644 627812 488645 627876
rect 488579 627811 488645 627812
rect 506611 627876 506677 627877
rect 506611 627812 506612 627876
rect 506676 627812 506677 627876
rect 506611 627811 506677 627812
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 466308 456134 492618
rect 459234 568894 459854 576000
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 466308 459854 496338
rect 462954 572614 463574 576000
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 466308 463574 500058
rect 469794 543454 470414 576000
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 466308 470414 470898
rect 473514 547174 474134 576000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 466308 474134 474618
rect 476070 472565 476130 627811
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 477234 550894 477854 576000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 476067 472564 476133 472565
rect 476067 472500 476068 472564
rect 476132 472500 476133 472564
rect 476067 472499 476133 472500
rect 477234 466308 477854 478338
rect 480954 554614 481574 576000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 466308 481574 482058
rect 487794 561454 488414 576000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 466308 488414 488898
rect 488582 486437 488642 627811
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 491514 565174 492134 576000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 488579 486436 488645 486437
rect 488579 486372 488580 486436
rect 488644 486372 488645 486436
rect 488579 486371 488645 486372
rect 491514 466308 492134 492618
rect 495234 568894 495854 576000
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 466308 495854 496338
rect 498954 572614 499574 576000
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498515 466580 498581 466581
rect 498515 466516 498516 466580
rect 498580 466516 498581 466580
rect 498515 466515 498581 466516
rect 498518 464810 498578 466515
rect 498954 466308 499574 500058
rect 505794 543454 506414 576000
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 506614 518125 506674 627811
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 509514 547174 510134 576000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 506611 518124 506677 518125
rect 506611 518060 506612 518124
rect 506676 518060 506677 518124
rect 506611 518059 506677 518060
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 466580 499869 466581
rect 499803 466516 499804 466580
rect 499868 466516 499869 466580
rect 499803 466515 499869 466516
rect 499806 464810 499866 466515
rect 505794 466308 506414 470898
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 466308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 466580 510909 466581
rect 510843 466516 510844 466580
rect 510908 466516 510909 466580
rect 510843 466515 510909 466516
rect 510846 464810 510906 466515
rect 513234 466308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 466308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 464750 498578 464810
rect 499688 464750 499866 464810
rect 510840 464750 510906 464810
rect 498464 464202 498524 464750
rect 499688 464202 499748 464750
rect 510840 464202 510900 464750
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 396056 380490 396116 381106
rect 397144 380490 397204 381106
rect 398232 380490 398292 381106
rect 399592 380490 399652 381106
rect 400544 380490 400604 381106
rect 401768 380490 401828 381106
rect 403128 380490 403188 381106
rect 404216 380490 404276 381106
rect 405440 380490 405500 381106
rect 406528 380490 406588 381106
rect 396030 380430 396116 380490
rect 397134 380430 397204 380490
rect 397502 380430 398292 380490
rect 399526 380430 399652 380490
rect 400446 380430 400604 380490
rect 401734 380430 401828 380490
rect 403022 380430 403188 380490
rect 404126 380430 404276 380490
rect 405414 380430 405500 380490
rect 406518 380430 406588 380490
rect 407616 380490 407676 381106
rect 408296 380490 408356 381106
rect 408704 380629 408764 381106
rect 408701 380628 408767 380629
rect 408701 380564 408702 380628
rect 408766 380564 408767 380628
rect 408701 380563 408767 380564
rect 410064 380490 410124 381106
rect 407616 380430 407682 380490
rect 408296 380430 408418 380490
rect 379794 364394 380414 379000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 359308 380414 363838
rect 383514 368114 384134 379000
rect 383514 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 384134 368114
rect 383514 367794 384134 367878
rect 383514 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 384134 367794
rect 383514 359308 384134 367558
rect 387234 369954 387854 379000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 359308 387854 369398
rect 390954 373674 391574 379000
rect 396030 378589 396090 380430
rect 397134 379405 397194 380430
rect 397131 379404 397197 379405
rect 397131 379340 397132 379404
rect 397196 379340 397197 379404
rect 397131 379339 397197 379340
rect 397502 378997 397562 380430
rect 397499 378996 397565 378997
rect 397499 378932 397500 378996
rect 397564 378932 397565 378996
rect 397499 378931 397565 378932
rect 396027 378588 396093 378589
rect 396027 378524 396028 378588
rect 396092 378524 396093 378588
rect 396027 378523 396093 378524
rect 390954 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 391574 373674
rect 390954 373354 391574 373438
rect 390954 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 391574 373354
rect 390954 359308 391574 373118
rect 397794 363454 398414 379000
rect 399526 378453 399586 380430
rect 400446 379405 400506 380430
rect 400443 379404 400509 379405
rect 400443 379340 400444 379404
rect 400508 379340 400509 379404
rect 400443 379339 400509 379340
rect 401734 379269 401794 380430
rect 403022 379269 403082 380430
rect 401731 379268 401797 379269
rect 401731 379204 401732 379268
rect 401796 379204 401797 379268
rect 401731 379203 401797 379204
rect 403019 379268 403085 379269
rect 403019 379204 403020 379268
rect 403084 379204 403085 379268
rect 403019 379203 403085 379204
rect 399523 378452 399589 378453
rect 399523 378388 399524 378452
rect 399588 378388 399589 378452
rect 399523 378387 399589 378388
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 359308 398414 362898
rect 401514 367174 402134 379000
rect 404126 378589 404186 380430
rect 405414 379269 405474 380430
rect 406518 379405 406578 380430
rect 407622 379405 407682 380430
rect 408358 379405 408418 380430
rect 410014 380430 410124 380490
rect 410744 380490 410804 381106
rect 411288 380490 411348 381106
rect 412376 380490 412436 381106
rect 413464 380629 413524 381106
rect 413461 380628 413527 380629
rect 413461 380564 413462 380628
rect 413526 380564 413527 380628
rect 413461 380563 413527 380564
rect 413600 380490 413660 381106
rect 410744 380430 410810 380490
rect 411288 380430 411362 380490
rect 412376 380430 412466 380490
rect 406515 379404 406581 379405
rect 406515 379340 406516 379404
rect 406580 379340 406581 379404
rect 406515 379339 406581 379340
rect 407619 379404 407685 379405
rect 407619 379340 407620 379404
rect 407684 379340 407685 379404
rect 407619 379339 407685 379340
rect 408355 379404 408421 379405
rect 408355 379340 408356 379404
rect 408420 379340 408421 379404
rect 408355 379339 408421 379340
rect 410014 379269 410074 380430
rect 410750 379405 410810 380430
rect 411302 379405 411362 380430
rect 412406 379405 412466 380430
rect 413510 380430 413660 380490
rect 414552 380490 414612 381106
rect 415912 380490 415972 381106
rect 414552 380430 414674 380490
rect 413510 379405 413570 380430
rect 410747 379404 410813 379405
rect 410747 379340 410748 379404
rect 410812 379340 410813 379404
rect 410747 379339 410813 379340
rect 411299 379404 411365 379405
rect 411299 379340 411300 379404
rect 411364 379340 411365 379404
rect 411299 379339 411365 379340
rect 412403 379404 412469 379405
rect 412403 379340 412404 379404
rect 412468 379340 412469 379404
rect 412403 379339 412469 379340
rect 413507 379404 413573 379405
rect 413507 379340 413508 379404
rect 413572 379340 413573 379404
rect 413507 379339 413573 379340
rect 414614 379269 414674 380430
rect 415902 380430 415972 380490
rect 416048 380490 416108 381106
rect 417000 380490 417060 381106
rect 418088 380490 418148 381106
rect 418496 380490 418556 381106
rect 419448 380490 419508 381106
rect 416048 380430 416146 380490
rect 417000 380430 417066 380490
rect 418088 380430 418170 380490
rect 415902 379269 415962 380430
rect 416086 379269 416146 380430
rect 405411 379268 405477 379269
rect 405411 379204 405412 379268
rect 405476 379204 405477 379268
rect 405411 379203 405477 379204
rect 410011 379268 410077 379269
rect 410011 379204 410012 379268
rect 410076 379204 410077 379268
rect 410011 379203 410077 379204
rect 414611 379268 414677 379269
rect 414611 379204 414612 379268
rect 414676 379204 414677 379268
rect 414611 379203 414677 379204
rect 415899 379268 415965 379269
rect 415899 379204 415900 379268
rect 415964 379204 415965 379268
rect 415899 379203 415965 379204
rect 416083 379268 416149 379269
rect 416083 379204 416084 379268
rect 416148 379204 416149 379268
rect 416083 379203 416149 379204
rect 404123 378588 404189 378589
rect 404123 378524 404124 378588
rect 404188 378524 404189 378588
rect 404123 378523 404189 378524
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 359308 402134 366618
rect 405234 370894 405854 379000
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 359308 405854 370338
rect 408954 374614 409574 379000
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 359308 409574 374058
rect 415794 364394 416414 379000
rect 417006 378181 417066 380430
rect 418110 378181 418170 380430
rect 418478 380430 418556 380490
rect 419398 380430 419508 380490
rect 420672 380490 420732 381106
rect 421080 380765 421140 381106
rect 421760 380765 421820 381106
rect 421077 380764 421143 380765
rect 421077 380700 421078 380764
rect 421142 380700 421143 380764
rect 421077 380699 421143 380700
rect 421757 380764 421823 380765
rect 421757 380700 421758 380764
rect 421822 380700 421823 380764
rect 421757 380699 421823 380700
rect 422848 380629 422908 381106
rect 422845 380628 422911 380629
rect 422845 380564 422846 380628
rect 422910 380564 422911 380628
rect 422845 380563 422911 380564
rect 423528 380490 423588 381106
rect 420672 380430 420746 380490
rect 418478 378861 418538 380430
rect 419398 379269 419458 380430
rect 419395 379268 419461 379269
rect 419395 379204 419396 379268
rect 419460 379204 419461 379268
rect 419395 379203 419461 379204
rect 418475 378860 418541 378861
rect 418475 378796 418476 378860
rect 418540 378796 418541 378860
rect 418475 378795 418541 378796
rect 417003 378180 417069 378181
rect 417003 378116 417004 378180
rect 417068 378116 417069 378180
rect 417003 378115 417069 378116
rect 418107 378180 418173 378181
rect 418107 378116 418108 378180
rect 418172 378116 418173 378180
rect 418107 378115 418173 378116
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 359308 416414 363838
rect 419514 368114 420134 379000
rect 420686 378181 420746 380430
rect 423446 380430 423588 380490
rect 423936 380490 423996 381106
rect 425296 380629 425356 381106
rect 425976 380765 426036 381106
rect 425973 380764 426039 380765
rect 425973 380700 425974 380764
rect 426038 380700 426039 380764
rect 425973 380699 426039 380700
rect 425293 380628 425359 380629
rect 425293 380564 425294 380628
rect 425358 380564 425359 380628
rect 425293 380563 425359 380564
rect 426384 380490 426444 381106
rect 427608 380490 427668 381106
rect 428288 380490 428348 381106
rect 428696 380490 428756 381106
rect 429784 380490 429844 381106
rect 431008 380490 431068 381106
rect 423936 380430 424058 380490
rect 426384 380430 426450 380490
rect 423446 379405 423506 380430
rect 423443 379404 423509 379405
rect 423443 379340 423444 379404
rect 423508 379340 423509 379404
rect 423443 379339 423509 379340
rect 420683 378180 420749 378181
rect 420683 378116 420684 378180
rect 420748 378116 420749 378180
rect 420683 378115 420749 378116
rect 419514 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 420134 368114
rect 419514 367794 420134 367878
rect 419514 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 420134 367794
rect 419514 359308 420134 367558
rect 423234 369954 423854 379000
rect 423998 378181 424058 380430
rect 426390 378181 426450 380430
rect 427494 380430 427668 380490
rect 428230 380430 428348 380490
rect 428598 380430 428756 380490
rect 429702 380430 429844 380490
rect 430990 380430 431068 380490
rect 431144 380490 431204 381106
rect 432232 380490 432292 381106
rect 433320 380490 433380 381106
rect 433592 380765 433652 381106
rect 434408 380765 434468 381106
rect 433589 380764 433655 380765
rect 433589 380700 433590 380764
rect 433654 380700 433655 380764
rect 433589 380699 433655 380700
rect 434405 380764 434471 380765
rect 434405 380700 434406 380764
rect 434470 380700 434471 380764
rect 434405 380699 434471 380700
rect 435768 380490 435828 381106
rect 436040 380765 436100 381106
rect 436037 380764 436103 380765
rect 436037 380700 436038 380764
rect 436102 380700 436103 380764
rect 436037 380699 436103 380700
rect 436992 380629 437052 381106
rect 436989 380628 437055 380629
rect 436989 380564 436990 380628
rect 437054 380564 437055 380628
rect 436989 380563 437055 380564
rect 438080 380490 438140 381106
rect 438488 380765 438548 381106
rect 438485 380764 438551 380765
rect 438485 380700 438486 380764
rect 438550 380700 438551 380764
rect 438485 380699 438551 380700
rect 439168 380490 439228 381106
rect 440936 380765 440996 381106
rect 443520 380765 443580 381106
rect 440933 380764 440999 380765
rect 440933 380700 440934 380764
rect 440998 380700 440999 380764
rect 440933 380699 440999 380700
rect 443517 380764 443583 380765
rect 443517 380700 443518 380764
rect 443582 380700 443583 380764
rect 443517 380699 443583 380700
rect 445968 380490 446028 381106
rect 431144 380430 431234 380490
rect 432232 380430 432338 380490
rect 433320 380430 433442 380490
rect 435768 380430 435834 380490
rect 427494 379405 427554 380430
rect 427491 379404 427557 379405
rect 427491 379340 427492 379404
rect 427556 379340 427557 379404
rect 427491 379339 427557 379340
rect 423995 378180 424061 378181
rect 423995 378116 423996 378180
rect 424060 378116 424061 378180
rect 423995 378115 424061 378116
rect 426387 378180 426453 378181
rect 426387 378116 426388 378180
rect 426452 378116 426453 378180
rect 426387 378115 426453 378116
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 359308 423854 369398
rect 426954 373674 427574 379000
rect 428230 378589 428290 380430
rect 428227 378588 428293 378589
rect 428227 378524 428228 378588
rect 428292 378524 428293 378588
rect 428227 378523 428293 378524
rect 428598 378317 428658 380430
rect 428595 378316 428661 378317
rect 428595 378252 428596 378316
rect 428660 378252 428661 378316
rect 428595 378251 428661 378252
rect 429702 378181 429762 380430
rect 430990 378589 431050 380430
rect 430987 378588 431053 378589
rect 430987 378524 430988 378588
rect 431052 378524 431053 378588
rect 430987 378523 431053 378524
rect 431174 378181 431234 380430
rect 432278 378181 432338 380430
rect 433382 379133 433442 380430
rect 433379 379132 433445 379133
rect 433379 379068 433380 379132
rect 433444 379068 433445 379132
rect 433379 379067 433445 379068
rect 429699 378180 429765 378181
rect 429699 378116 429700 378180
rect 429764 378116 429765 378180
rect 429699 378115 429765 378116
rect 431171 378180 431237 378181
rect 431171 378116 431172 378180
rect 431236 378116 431237 378180
rect 431171 378115 431237 378116
rect 432275 378180 432341 378181
rect 432275 378116 432276 378180
rect 432340 378116 432341 378180
rect 432275 378115 432341 378116
rect 426954 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 427574 373674
rect 426954 373354 427574 373438
rect 426954 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 427574 373354
rect 426954 359308 427574 373118
rect 433794 363454 434414 379000
rect 435774 378725 435834 380430
rect 437982 380430 438140 380490
rect 439086 380430 439228 380490
rect 445894 380430 446028 380490
rect 448280 380490 448340 381106
rect 451000 380490 451060 381106
rect 453448 380490 453508 381106
rect 455896 380490 455956 381106
rect 458480 380490 458540 381106
rect 448280 380430 448346 380490
rect 451000 380430 451106 380490
rect 437982 379269 438042 380430
rect 439086 379405 439146 380430
rect 445894 379405 445954 380430
rect 448286 379405 448346 380430
rect 451046 379405 451106 380430
rect 453438 380430 453508 380490
rect 455830 380430 455956 380490
rect 458406 380430 458540 380490
rect 460928 380490 460988 381106
rect 463512 380490 463572 381106
rect 465960 380629 466020 381106
rect 465957 380628 466023 380629
rect 465957 380564 465958 380628
rect 466022 380564 466023 380628
rect 465957 380563 466023 380564
rect 468544 380490 468604 381106
rect 470992 380490 471052 381106
rect 460928 380430 461042 380490
rect 463512 380430 463618 380490
rect 453438 379405 453498 380430
rect 455830 379405 455890 380430
rect 458406 379405 458466 380430
rect 439083 379404 439149 379405
rect 439083 379340 439084 379404
rect 439148 379340 439149 379404
rect 439083 379339 439149 379340
rect 445891 379404 445957 379405
rect 445891 379340 445892 379404
rect 445956 379340 445957 379404
rect 445891 379339 445957 379340
rect 448283 379404 448349 379405
rect 448283 379340 448284 379404
rect 448348 379340 448349 379404
rect 448283 379339 448349 379340
rect 451043 379404 451109 379405
rect 451043 379340 451044 379404
rect 451108 379340 451109 379404
rect 451043 379339 451109 379340
rect 453435 379404 453501 379405
rect 453435 379340 453436 379404
rect 453500 379340 453501 379404
rect 453435 379339 453501 379340
rect 455827 379404 455893 379405
rect 455827 379340 455828 379404
rect 455892 379340 455893 379404
rect 455827 379339 455893 379340
rect 458403 379404 458469 379405
rect 458403 379340 458404 379404
rect 458468 379340 458469 379404
rect 458403 379339 458469 379340
rect 437979 379268 438045 379269
rect 437979 379204 437980 379268
rect 438044 379204 438045 379268
rect 437979 379203 438045 379204
rect 435771 378724 435837 378725
rect 435771 378660 435772 378724
rect 435836 378660 435837 378724
rect 435771 378659 435837 378660
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 359308 434414 362898
rect 437514 367174 438134 379000
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 359308 438134 366618
rect 441234 370894 441854 379000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 359308 441854 370338
rect 444954 374614 445574 379000
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 359308 445574 374058
rect 451794 364394 452414 379000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 359308 452414 363838
rect 455514 368114 456134 379000
rect 455514 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 456134 368114
rect 455514 367794 456134 367878
rect 455514 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 456134 367794
rect 455514 359308 456134 367558
rect 459234 369954 459854 379000
rect 460982 378181 461042 380430
rect 463558 379269 463618 380430
rect 468526 380430 468604 380490
rect 470918 380430 471052 380490
rect 473440 380490 473500 381106
rect 475888 380490 475948 381106
rect 478472 380490 478532 381106
rect 480920 380490 480980 381106
rect 473440 380430 473554 380490
rect 463555 379268 463621 379269
rect 463555 379204 463556 379268
rect 463620 379204 463621 379268
rect 463555 379203 463621 379204
rect 460979 378180 461045 378181
rect 460979 378116 460980 378180
rect 461044 378116 461045 378180
rect 460979 378115 461045 378116
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 359308 459854 369398
rect 462954 373674 463574 379000
rect 468526 378861 468586 380430
rect 468523 378860 468589 378861
rect 468523 378796 468524 378860
rect 468588 378796 468589 378860
rect 468523 378795 468589 378796
rect 462954 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 463574 373674
rect 462954 373354 463574 373438
rect 462954 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 463574 373354
rect 462954 359308 463574 373118
rect 469794 363454 470414 379000
rect 470918 378861 470978 380430
rect 473494 379269 473554 380430
rect 475886 380430 475948 380490
rect 478462 380430 478532 380490
rect 480854 380430 480980 380490
rect 483368 380490 483428 381106
rect 485952 380901 486012 381106
rect 485949 380900 486015 380901
rect 485949 380836 485950 380900
rect 486014 380836 486015 380900
rect 485949 380835 486015 380836
rect 503224 380490 503284 381106
rect 483368 380430 483490 380490
rect 475886 379269 475946 380430
rect 473491 379268 473557 379269
rect 473491 379204 473492 379268
rect 473556 379204 473557 379268
rect 473491 379203 473557 379204
rect 475883 379268 475949 379269
rect 475883 379204 475884 379268
rect 475948 379204 475949 379268
rect 475883 379203 475949 379204
rect 470915 378860 470981 378861
rect 470915 378796 470916 378860
rect 470980 378796 470981 378860
rect 470915 378795 470981 378796
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 359308 470414 362898
rect 473514 367174 474134 379000
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 359308 474134 366618
rect 477234 370894 477854 379000
rect 478462 378861 478522 380430
rect 480854 379269 480914 380430
rect 480851 379268 480917 379269
rect 480851 379204 480852 379268
rect 480916 379204 480917 379268
rect 480851 379203 480917 379204
rect 478459 378860 478525 378861
rect 478459 378796 478460 378860
rect 478524 378796 478525 378860
rect 478459 378795 478525 378796
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 359308 477854 370338
rect 480954 374614 481574 379000
rect 483430 378861 483490 380430
rect 503118 380430 503284 380490
rect 503360 380490 503420 381106
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 503360 380430 503546 380490
rect 503118 379269 503178 380430
rect 503486 379269 503546 380430
rect 503115 379268 503181 379269
rect 503115 379204 503116 379268
rect 503180 379204 503181 379268
rect 503115 379203 503181 379204
rect 503483 379268 503549 379269
rect 503483 379204 503484 379268
rect 503548 379204 503549 379268
rect 503483 379203 503549 379204
rect 483427 378860 483493 378861
rect 483427 378796 483428 378860
rect 483492 378796 483493 378860
rect 483427 378795 483493 378796
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 359308 481574 374058
rect 487794 364394 488414 379000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 359308 488414 363838
rect 491514 368114 492134 379000
rect 491514 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 491514 367794 492134 367878
rect 491514 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 491514 359308 492134 367558
rect 495234 369954 495854 379000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 359308 495854 369398
rect 498954 373674 499574 379000
rect 498954 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 498954 373354 499574 373438
rect 498954 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 498954 359308 499574 373118
rect 505794 363454 506414 379000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 359308 506414 362898
rect 509514 367174 510134 379000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 359308 510134 366618
rect 513234 370894 513854 379000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 359308 513854 370338
rect 516954 374614 517574 379000
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 359308 517574 374058
rect 498515 358868 498581 358869
rect 498515 358804 498516 358868
rect 498580 358804 498581 358868
rect 498515 358803 498581 358804
rect 499803 358868 499869 358869
rect 499803 358804 499804 358868
rect 499868 358804 499869 358868
rect 499803 358803 499869 358804
rect 510843 358868 510909 358869
rect 510843 358804 510844 358868
rect 510908 358804 510909 358868
rect 510843 358803 510909 358804
rect 498518 358050 498578 358803
rect 499806 358050 499866 358803
rect 510846 358050 510906 358803
rect 498464 357990 498578 358050
rect 499688 357990 499866 358050
rect 510840 357990 510906 358050
rect 498464 357202 498524 357990
rect 499688 357202 499748 357990
rect 510840 357202 510900 357990
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 396056 273730 396116 274040
rect 397144 273730 397204 274040
rect 398232 273730 398292 274040
rect 399592 273730 399652 274040
rect 400544 273730 400604 274040
rect 401768 273730 401828 274040
rect 403128 273730 403188 274040
rect 404216 273730 404276 274040
rect 405440 273730 405500 274040
rect 406528 273730 406588 274040
rect 396030 273670 396116 273730
rect 397134 273670 397204 273730
rect 397502 273670 398292 273730
rect 399526 273670 399652 273730
rect 400446 273670 400604 273730
rect 401734 273670 401828 273730
rect 403022 273670 403188 273730
rect 404126 273670 404276 273730
rect 405046 273670 405500 273730
rect 406518 273670 406588 273730
rect 407616 273730 407676 274040
rect 408296 273730 408356 274040
rect 407616 273670 407682 273730
rect 379794 256394 380414 272000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 252308 380414 255838
rect 383514 260114 384134 272000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 252308 384134 259558
rect 387234 261954 387854 272000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 252308 387854 261398
rect 390954 265674 391574 272000
rect 396030 271285 396090 273670
rect 396027 271284 396093 271285
rect 396027 271220 396028 271284
rect 396092 271220 396093 271284
rect 396027 271219 396093 271220
rect 397134 270605 397194 273670
rect 397502 270605 397562 273670
rect 397131 270604 397197 270605
rect 397131 270540 397132 270604
rect 397196 270540 397197 270604
rect 397131 270539 397197 270540
rect 397499 270604 397565 270605
rect 397499 270540 397500 270604
rect 397564 270540 397565 270604
rect 397499 270539 397565 270540
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 252308 391574 265118
rect 397794 255454 398414 272000
rect 399526 270605 399586 273670
rect 400446 270605 400506 273670
rect 401734 272237 401794 273670
rect 401731 272236 401797 272237
rect 401731 272172 401732 272236
rect 401796 272172 401797 272236
rect 401731 272171 401797 272172
rect 399523 270604 399589 270605
rect 399523 270540 399524 270604
rect 399588 270540 399589 270604
rect 399523 270539 399589 270540
rect 400443 270604 400509 270605
rect 400443 270540 400444 270604
rect 400508 270540 400509 270604
rect 400443 270539 400509 270540
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252308 398414 254898
rect 401514 259174 402134 272000
rect 403022 271829 403082 273670
rect 403019 271828 403085 271829
rect 403019 271764 403020 271828
rect 403084 271764 403085 271828
rect 403019 271763 403085 271764
rect 404126 270605 404186 273670
rect 405046 271013 405106 273670
rect 405043 271012 405109 271013
rect 405043 270948 405044 271012
rect 405108 270948 405109 271012
rect 405043 270947 405109 270948
rect 404123 270604 404189 270605
rect 404123 270540 404124 270604
rect 404188 270540 404189 270604
rect 404123 270539 404189 270540
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252308 402134 258618
rect 405234 262894 405854 272000
rect 406518 270605 406578 273670
rect 407622 270605 407682 273670
rect 408174 273670 408356 273730
rect 408704 273730 408764 274040
rect 410064 273730 410124 274040
rect 408704 273670 408786 273730
rect 408174 271013 408234 273670
rect 408171 271012 408237 271013
rect 408171 270948 408172 271012
rect 408236 270948 408237 271012
rect 408171 270947 408237 270948
rect 408726 270605 408786 273670
rect 410014 273670 410124 273730
rect 410744 273730 410804 274040
rect 411288 273730 411348 274040
rect 412376 273730 412436 274040
rect 413464 273730 413524 274040
rect 410744 273670 410810 273730
rect 411288 273670 411362 273730
rect 412376 273670 412466 273730
rect 406515 270604 406581 270605
rect 406515 270540 406516 270604
rect 406580 270540 406581 270604
rect 406515 270539 406581 270540
rect 407619 270604 407685 270605
rect 407619 270540 407620 270604
rect 407684 270540 407685 270604
rect 407619 270539 407685 270540
rect 408723 270604 408789 270605
rect 408723 270540 408724 270604
rect 408788 270540 408789 270604
rect 408723 270539 408789 270540
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252308 405854 262338
rect 408954 266614 409574 272000
rect 410014 270605 410074 273670
rect 410750 271149 410810 273670
rect 410747 271148 410813 271149
rect 410747 271084 410748 271148
rect 410812 271084 410813 271148
rect 410747 271083 410813 271084
rect 411302 270605 411362 273670
rect 412406 271013 412466 273670
rect 413326 273670 413524 273730
rect 413600 273730 413660 274040
rect 414552 273730 414612 274040
rect 415912 273730 415972 274040
rect 413600 273670 413754 273730
rect 412403 271012 412469 271013
rect 412403 270948 412404 271012
rect 412468 270948 412469 271012
rect 412403 270947 412469 270948
rect 413326 270741 413386 273670
rect 413694 271285 413754 273670
rect 414430 273670 414612 273730
rect 415534 273670 415972 273730
rect 416048 273730 416108 274040
rect 417000 273730 417060 274040
rect 418088 273730 418148 274040
rect 418496 273730 418556 274040
rect 419448 273730 419508 274040
rect 416048 273670 416146 273730
rect 417000 273670 417066 273730
rect 418088 273670 418170 273730
rect 413691 271284 413757 271285
rect 413691 271220 413692 271284
rect 413756 271220 413757 271284
rect 413691 271219 413757 271220
rect 414430 271149 414490 273670
rect 415534 271421 415594 273670
rect 416086 272237 416146 273670
rect 416083 272236 416149 272237
rect 416083 272172 416084 272236
rect 416148 272172 416149 272236
rect 416083 272171 416149 272172
rect 415531 271420 415597 271421
rect 415531 271356 415532 271420
rect 415596 271356 415597 271420
rect 415531 271355 415597 271356
rect 414427 271148 414493 271149
rect 414427 271084 414428 271148
rect 414492 271084 414493 271148
rect 414427 271083 414493 271084
rect 413323 270740 413389 270741
rect 413323 270676 413324 270740
rect 413388 270676 413389 270740
rect 413323 270675 413389 270676
rect 410011 270604 410077 270605
rect 410011 270540 410012 270604
rect 410076 270540 410077 270604
rect 410011 270539 410077 270540
rect 411299 270604 411365 270605
rect 411299 270540 411300 270604
rect 411364 270540 411365 270604
rect 411299 270539 411365 270540
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252308 409574 266058
rect 415794 256394 416414 272000
rect 417006 271149 417066 273670
rect 417003 271148 417069 271149
rect 417003 271084 417004 271148
rect 417068 271084 417069 271148
rect 417003 271083 417069 271084
rect 418110 270605 418170 273670
rect 418478 273670 418556 273730
rect 419214 273670 419508 273730
rect 420672 273730 420732 274040
rect 420672 273670 420746 273730
rect 418478 271829 418538 273670
rect 418475 271828 418541 271829
rect 418475 271764 418476 271828
rect 418540 271764 418541 271828
rect 418475 271763 418541 271764
rect 419214 270741 419274 273670
rect 419211 270740 419277 270741
rect 419211 270676 419212 270740
rect 419276 270676 419277 270740
rect 419211 270675 419277 270676
rect 418107 270604 418173 270605
rect 418107 270540 418108 270604
rect 418172 270540 418173 270604
rect 418107 270539 418173 270540
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 252308 416414 255838
rect 419514 260114 420134 272000
rect 420686 270605 420746 273670
rect 421080 273597 421140 274040
rect 421760 273730 421820 274040
rect 422848 273730 422908 274040
rect 423528 273730 423588 274040
rect 423936 273730 423996 274040
rect 425296 273730 425356 274040
rect 421760 273670 421850 273730
rect 422848 273670 422954 273730
rect 421077 273596 421143 273597
rect 421077 273532 421078 273596
rect 421142 273532 421143 273596
rect 421077 273531 421143 273532
rect 421790 270605 421850 273670
rect 422894 273461 422954 273670
rect 423446 273670 423588 273730
rect 423814 273670 423996 273730
rect 425286 273670 425356 273730
rect 425976 273730 426036 274040
rect 426384 273730 426444 274040
rect 427608 273730 427668 274040
rect 428288 273730 428348 274040
rect 428696 273730 428756 274040
rect 429784 273730 429844 274040
rect 431008 273730 431068 274040
rect 425976 273670 426082 273730
rect 426384 273670 426450 273730
rect 427608 273670 427738 273730
rect 422891 273460 422957 273461
rect 422891 273396 422892 273460
rect 422956 273396 422957 273460
rect 422891 273395 422957 273396
rect 423446 273325 423506 273670
rect 423814 273325 423874 273670
rect 423443 273324 423509 273325
rect 423443 273260 423444 273324
rect 423508 273260 423509 273324
rect 423443 273259 423509 273260
rect 423811 273324 423877 273325
rect 423811 273260 423812 273324
rect 423876 273260 423877 273324
rect 423811 273259 423877 273260
rect 420683 270604 420749 270605
rect 420683 270540 420684 270604
rect 420748 270540 420749 270604
rect 420683 270539 420749 270540
rect 421787 270604 421853 270605
rect 421787 270540 421788 270604
rect 421852 270540 421853 270604
rect 421787 270539 421853 270540
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 252308 420134 259558
rect 423234 261954 423854 272000
rect 425286 270333 425346 273670
rect 426022 272781 426082 273670
rect 426390 273325 426450 273670
rect 426387 273324 426453 273325
rect 426387 273260 426388 273324
rect 426452 273260 426453 273324
rect 426387 273259 426453 273260
rect 426019 272780 426085 272781
rect 426019 272716 426020 272780
rect 426084 272716 426085 272780
rect 426019 272715 426085 272716
rect 425283 270332 425349 270333
rect 425283 270268 425284 270332
rect 425348 270268 425349 270332
rect 425283 270267 425349 270268
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 252308 423854 261398
rect 426954 265674 427574 272000
rect 427678 270741 427738 273670
rect 428230 273670 428348 273730
rect 428598 273670 428756 273730
rect 429702 273670 429844 273730
rect 430990 273670 431068 273730
rect 431144 273730 431204 274040
rect 432232 273730 432292 274040
rect 433320 273730 433380 274040
rect 433592 273730 433652 274040
rect 431144 273670 431234 273730
rect 432232 273670 432338 273730
rect 433320 273670 433442 273730
rect 428230 272781 428290 273670
rect 428227 272780 428293 272781
rect 428227 272716 428228 272780
rect 428292 272716 428293 272780
rect 428227 272715 428293 272716
rect 428598 271013 428658 273670
rect 429702 271013 429762 273670
rect 430990 273461 431050 273670
rect 430987 273460 431053 273461
rect 430987 273396 430988 273460
rect 431052 273396 431053 273460
rect 430987 273395 431053 273396
rect 431174 272781 431234 273670
rect 431171 272780 431237 272781
rect 431171 272716 431172 272780
rect 431236 272716 431237 272780
rect 431171 272715 431237 272716
rect 428595 271012 428661 271013
rect 428595 270948 428596 271012
rect 428660 270948 428661 271012
rect 428595 270947 428661 270948
rect 429699 271012 429765 271013
rect 429699 270948 429700 271012
rect 429764 270948 429765 271012
rect 429699 270947 429765 270948
rect 427675 270740 427741 270741
rect 427675 270676 427676 270740
rect 427740 270676 427741 270740
rect 427675 270675 427741 270676
rect 432278 270469 432338 273670
rect 433382 271013 433442 273670
rect 433566 273670 433652 273730
rect 434408 273730 434468 274040
rect 435768 273730 435828 274040
rect 436040 273730 436100 274040
rect 436992 273730 437052 274040
rect 438080 273730 438140 274040
rect 434408 273670 434730 273730
rect 435768 273670 435834 273730
rect 433566 271829 433626 273670
rect 433563 271828 433629 271829
rect 433563 271764 433564 271828
rect 433628 271764 433629 271828
rect 433563 271763 433629 271764
rect 433379 271012 433445 271013
rect 433379 270948 433380 271012
rect 433444 270948 433445 271012
rect 433379 270947 433445 270948
rect 432275 270468 432341 270469
rect 432275 270404 432276 270468
rect 432340 270404 432341 270468
rect 432275 270403 432341 270404
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 252308 427574 265118
rect 433794 255454 434414 272000
rect 434670 271149 434730 273670
rect 434667 271148 434733 271149
rect 434667 271084 434668 271148
rect 434732 271084 434733 271148
rect 434667 271083 434733 271084
rect 435774 271013 435834 273670
rect 435958 273670 436100 273730
rect 436878 273670 437052 273730
rect 437982 273670 438140 273730
rect 438488 273730 438548 274040
rect 439168 273730 439228 274040
rect 440936 273730 440996 274040
rect 443520 273730 443580 274040
rect 445968 273730 446028 274040
rect 438488 273670 438594 273730
rect 439168 273670 439330 273730
rect 435958 271829 436018 273670
rect 435955 271828 436021 271829
rect 435955 271764 435956 271828
rect 436020 271764 436021 271828
rect 435955 271763 436021 271764
rect 435771 271012 435837 271013
rect 435771 270948 435772 271012
rect 435836 270948 435837 271012
rect 435771 270947 435837 270948
rect 436878 270605 436938 273670
rect 437982 272237 438042 273670
rect 437979 272236 438045 272237
rect 437979 272172 437980 272236
rect 438044 272172 438045 272236
rect 437979 272171 438045 272172
rect 436875 270604 436941 270605
rect 436875 270540 436876 270604
rect 436940 270540 436941 270604
rect 436875 270539 436941 270540
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 252308 434414 254898
rect 437514 259174 438134 272000
rect 438534 271829 438594 273670
rect 438531 271828 438597 271829
rect 438531 271764 438532 271828
rect 438596 271764 438597 271828
rect 438531 271763 438597 271764
rect 439270 271285 439330 273670
rect 440926 273670 440996 273730
rect 443502 273670 443580 273730
rect 445894 273670 446028 273730
rect 448280 273730 448340 274040
rect 448280 273670 448346 273730
rect 440926 271421 440986 273670
rect 440923 271420 440989 271421
rect 440923 271356 440924 271420
rect 440988 271356 440989 271420
rect 440923 271355 440989 271356
rect 439267 271284 439333 271285
rect 439267 271220 439268 271284
rect 439332 271220 439333 271284
rect 439267 271219 439333 271220
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 252308 438134 258618
rect 441234 262894 441854 272000
rect 443502 271285 443562 273670
rect 443499 271284 443565 271285
rect 443499 271220 443500 271284
rect 443564 271220 443565 271284
rect 443499 271219 443565 271220
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 252308 441854 262338
rect 444954 266614 445574 272000
rect 445894 271829 445954 273670
rect 448286 271829 448346 273670
rect 451000 273597 451060 274040
rect 450997 273596 451063 273597
rect 450997 273532 450998 273596
rect 451062 273532 451063 273596
rect 453448 273594 453508 274040
rect 455896 273594 455956 274040
rect 458480 273594 458540 274040
rect 460928 273730 460988 274040
rect 463512 273730 463572 274040
rect 465960 273730 466020 274040
rect 468544 273730 468604 274040
rect 470992 273730 471052 274040
rect 460928 273670 461042 273730
rect 450997 273531 451063 273532
rect 453438 273534 453508 273594
rect 455830 273534 455956 273594
rect 458406 273534 458540 273594
rect 445891 271828 445957 271829
rect 445891 271764 445892 271828
rect 445956 271764 445957 271828
rect 445891 271763 445957 271764
rect 448283 271828 448349 271829
rect 448283 271764 448284 271828
rect 448348 271764 448349 271828
rect 448283 271763 448349 271764
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 252308 445574 266058
rect 451794 256394 452414 272000
rect 453438 271829 453498 273534
rect 455830 272237 455890 273534
rect 455827 272236 455893 272237
rect 455827 272172 455828 272236
rect 455892 272172 455893 272236
rect 455827 272171 455893 272172
rect 453435 271828 453501 271829
rect 453435 271764 453436 271828
rect 453500 271764 453501 271828
rect 453435 271763 453501 271764
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 252308 452414 255838
rect 455514 260114 456134 272000
rect 458406 271829 458466 273534
rect 458403 271828 458469 271829
rect 458403 271764 458404 271828
rect 458468 271764 458469 271828
rect 458403 271763 458469 271764
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 252308 456134 259558
rect 459234 261954 459854 272000
rect 460982 271557 461042 273670
rect 462638 273670 463572 273730
rect 465950 273670 466020 273730
rect 468526 273670 468604 273730
rect 470918 273670 471052 273730
rect 473440 273730 473500 274040
rect 475888 273730 475948 274040
rect 478472 273730 478532 274040
rect 480920 273730 480980 274040
rect 483368 273730 483428 274040
rect 473440 273670 473554 273730
rect 460979 271556 461045 271557
rect 460979 271492 460980 271556
rect 461044 271492 461045 271556
rect 460979 271491 461045 271492
rect 462638 270877 462698 273670
rect 462635 270876 462701 270877
rect 462635 270812 462636 270876
rect 462700 270812 462701 270876
rect 462635 270811 462701 270812
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 252308 459854 261398
rect 462954 265674 463574 272000
rect 465950 271693 466010 273670
rect 468526 272781 468586 273670
rect 470918 272781 470978 273670
rect 473494 272781 473554 273670
rect 475886 273670 475948 273730
rect 478462 273670 478532 273730
rect 480854 273670 480980 273730
rect 483246 273670 483428 273730
rect 485952 273730 486012 274040
rect 503224 273730 503284 274040
rect 485952 273670 486066 273730
rect 468523 272780 468589 272781
rect 468523 272716 468524 272780
rect 468588 272716 468589 272780
rect 468523 272715 468589 272716
rect 470915 272780 470981 272781
rect 470915 272716 470916 272780
rect 470980 272716 470981 272780
rect 470915 272715 470981 272716
rect 473491 272780 473557 272781
rect 473491 272716 473492 272780
rect 473556 272716 473557 272780
rect 473491 272715 473557 272716
rect 475886 272645 475946 273670
rect 478462 272645 478522 273670
rect 480854 272917 480914 273670
rect 483246 273053 483306 273670
rect 486006 273189 486066 273670
rect 503118 273670 503284 273730
rect 503360 273730 503420 274040
rect 503360 273670 503546 273730
rect 486003 273188 486069 273189
rect 486003 273124 486004 273188
rect 486068 273124 486069 273188
rect 486003 273123 486069 273124
rect 483243 273052 483309 273053
rect 483243 272988 483244 273052
rect 483308 272988 483309 273052
rect 483243 272987 483309 272988
rect 480851 272916 480917 272917
rect 480851 272852 480852 272916
rect 480916 272852 480917 272916
rect 480851 272851 480917 272852
rect 475883 272644 475949 272645
rect 475883 272580 475884 272644
rect 475948 272580 475949 272644
rect 475883 272579 475949 272580
rect 478459 272644 478525 272645
rect 478459 272580 478460 272644
rect 478524 272580 478525 272644
rect 478459 272579 478525 272580
rect 465947 271692 466013 271693
rect 465947 271628 465948 271692
rect 466012 271628 466013 271692
rect 465947 271627 466013 271628
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 252308 463574 265118
rect 469794 255454 470414 272000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 252308 470414 254898
rect 473514 259174 474134 272000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 252308 474134 258618
rect 477234 262894 477854 272000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 252308 477854 262338
rect 480954 266614 481574 272000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 252308 481574 266058
rect 487794 256394 488414 272000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 252308 488414 255838
rect 491514 260114 492134 272000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 252308 492134 259558
rect 495234 261954 495854 272000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 252308 495854 261398
rect 498954 265674 499574 272000
rect 503118 271693 503178 273670
rect 503115 271692 503181 271693
rect 503115 271628 503116 271692
rect 503180 271628 503181 271692
rect 503115 271627 503181 271628
rect 503486 271285 503546 273670
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 503483 271284 503549 271285
rect 503483 271220 503484 271284
rect 503548 271220 503549 271284
rect 503483 271219 503549 271220
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498515 252788 498581 252789
rect 498515 252724 498516 252788
rect 498580 252724 498581 252788
rect 498515 252723 498581 252724
rect 498518 250610 498578 252723
rect 498954 252308 499574 265118
rect 505794 255454 506414 272000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 499803 253332 499869 253333
rect 499803 253268 499804 253332
rect 499868 253268 499869 253332
rect 499803 253267 499869 253268
rect 499806 250610 499866 253267
rect 505794 252308 506414 254898
rect 509514 259174 510134 272000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 252308 510134 258618
rect 513234 262894 513854 272000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 510843 252652 510909 252653
rect 510843 252588 510844 252652
rect 510908 252588 510909 252652
rect 510843 252587 510909 252588
rect 510846 250610 510906 252587
rect 513234 252308 513854 262338
rect 516954 266614 517574 272000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 252308 517574 266058
rect 498464 250550 498578 250610
rect 499688 250550 499866 250610
rect 510840 250550 510906 250610
rect 498464 250240 498524 250550
rect 499688 250240 499748 250550
rect 510840 250240 510900 250550
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 379470 171090 379714 171150
rect 379470 165069 379530 171090
rect 396056 167010 396116 167106
rect 397144 167010 397204 167106
rect 396030 166950 396116 167010
rect 397134 166950 397204 167010
rect 398232 167010 398292 167106
rect 399592 167010 399652 167106
rect 400544 167010 400604 167106
rect 401768 167010 401828 167106
rect 403128 167010 403188 167106
rect 404216 167010 404276 167106
rect 405440 167010 405500 167106
rect 406528 167010 406588 167106
rect 398232 166950 398298 167010
rect 379467 165068 379533 165069
rect 379467 165004 379468 165068
rect 379532 165004 379533 165068
rect 379467 165003 379533 165004
rect 379794 148394 380414 165000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379794 145308 380414 147838
rect 383514 152114 384134 165000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 155834 387854 165000
rect 387234 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 387854 155834
rect 387234 155514 387854 155598
rect 387234 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 387854 155514
rect 387234 145308 387854 155278
rect 390954 157674 391574 165000
rect 396030 164253 396090 166950
rect 397134 164389 397194 166950
rect 398238 165613 398298 166950
rect 399526 166950 399652 167010
rect 400446 166950 400604 167010
rect 401734 166950 401828 167010
rect 403022 166950 403188 167010
rect 404126 166950 404276 167010
rect 405414 166950 405500 167010
rect 406518 166950 406588 167010
rect 407616 167010 407676 167106
rect 408296 167010 408356 167106
rect 407616 166950 407682 167010
rect 398235 165612 398301 165613
rect 398235 165548 398236 165612
rect 398300 165548 398301 165612
rect 398235 165547 398301 165548
rect 397131 164388 397197 164389
rect 397131 164324 397132 164388
rect 397196 164324 397197 164388
rect 397131 164323 397197 164324
rect 396027 164252 396093 164253
rect 396027 164188 396028 164252
rect 396092 164188 396093 164252
rect 396027 164187 396093 164188
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 165000
rect 399526 164253 399586 166950
rect 400446 164253 400506 166950
rect 401734 165613 401794 166950
rect 401731 165612 401797 165613
rect 401731 165548 401732 165612
rect 401796 165548 401797 165612
rect 401731 165547 401797 165548
rect 399523 164252 399589 164253
rect 399523 164188 399524 164252
rect 399588 164188 399589 164252
rect 399523 164187 399589 164188
rect 400443 164252 400509 164253
rect 400443 164188 400444 164252
rect 400508 164188 400509 164252
rect 400443 164187 400509 164188
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 165000
rect 403022 164253 403082 166950
rect 404126 164389 404186 166950
rect 405414 165613 405474 166950
rect 405411 165612 405477 165613
rect 405411 165548 405412 165612
rect 405476 165548 405477 165612
rect 405411 165547 405477 165548
rect 404123 164388 404189 164389
rect 404123 164324 404124 164388
rect 404188 164324 404189 164388
rect 404123 164323 404189 164324
rect 403019 164252 403085 164253
rect 403019 164188 403020 164252
rect 403084 164188 403085 164252
rect 403019 164187 403085 164188
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 165000
rect 406518 164253 406578 166950
rect 407622 164253 407682 166950
rect 408174 166950 408356 167010
rect 408704 167010 408764 167106
rect 410064 167010 410124 167106
rect 408704 166950 408786 167010
rect 408174 165613 408234 166950
rect 408171 165612 408237 165613
rect 408171 165548 408172 165612
rect 408236 165548 408237 165612
rect 408171 165547 408237 165548
rect 408726 164253 408786 166950
rect 410014 166950 410124 167010
rect 410744 167010 410804 167106
rect 411288 167010 411348 167106
rect 412376 167010 412436 167106
rect 413464 167010 413524 167106
rect 410744 166950 410810 167010
rect 411288 166950 411362 167010
rect 412376 166950 412466 167010
rect 406515 164252 406581 164253
rect 406515 164188 406516 164252
rect 406580 164188 406581 164252
rect 406515 164187 406581 164188
rect 407619 164252 407685 164253
rect 407619 164188 407620 164252
rect 407684 164188 407685 164252
rect 407619 164187 407685 164188
rect 408723 164252 408789 164253
rect 408723 164188 408724 164252
rect 408788 164188 408789 164252
rect 408723 164187 408789 164188
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 165000
rect 410014 164253 410074 166950
rect 410750 165613 410810 166950
rect 410747 165612 410813 165613
rect 410747 165548 410748 165612
rect 410812 165548 410813 165612
rect 410747 165547 410813 165548
rect 411302 164253 411362 166950
rect 412406 164389 412466 166950
rect 413326 166950 413524 167010
rect 413600 167010 413660 167106
rect 414552 167010 414612 167106
rect 415912 167010 415972 167106
rect 413600 166950 413754 167010
rect 412403 164388 412469 164389
rect 412403 164324 412404 164388
rect 412468 164324 412469 164388
rect 412403 164323 412469 164324
rect 413326 164253 413386 166950
rect 413694 164797 413754 166950
rect 414430 166950 414612 167010
rect 415902 166950 415972 167010
rect 416048 167010 416108 167106
rect 417000 167010 417060 167106
rect 418088 167010 418148 167106
rect 418496 167010 418556 167106
rect 419448 167010 419508 167106
rect 416048 166950 416146 167010
rect 417000 166950 417066 167010
rect 418088 166950 418354 167010
rect 413691 164796 413757 164797
rect 413691 164732 413692 164796
rect 413756 164732 413757 164796
rect 413691 164731 413757 164732
rect 414430 164253 414490 166950
rect 415902 165613 415962 166950
rect 416086 165613 416146 166950
rect 415899 165612 415965 165613
rect 415899 165548 415900 165612
rect 415964 165548 415965 165612
rect 415899 165547 415965 165548
rect 416083 165612 416149 165613
rect 416083 165548 416084 165612
rect 416148 165548 416149 165612
rect 416083 165547 416149 165548
rect 410011 164252 410077 164253
rect 410011 164188 410012 164252
rect 410076 164188 410077 164252
rect 410011 164187 410077 164188
rect 411299 164252 411365 164253
rect 411299 164188 411300 164252
rect 411364 164188 411365 164252
rect 411299 164187 411365 164188
rect 413323 164252 413389 164253
rect 413323 164188 413324 164252
rect 413388 164188 413389 164252
rect 413323 164187 413389 164188
rect 414427 164252 414493 164253
rect 414427 164188 414428 164252
rect 414492 164188 414493 164252
rect 414427 164187 414493 164188
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 165000
rect 417006 164253 417066 166950
rect 418294 164253 418354 166950
rect 418478 166950 418556 167010
rect 419398 166950 419508 167010
rect 420672 167010 420732 167106
rect 421080 167010 421140 167106
rect 420672 166950 420746 167010
rect 418478 166837 418538 166950
rect 418475 166836 418541 166837
rect 418475 166772 418476 166836
rect 418540 166772 418541 166836
rect 418475 166771 418541 166772
rect 419398 165613 419458 166950
rect 419395 165612 419461 165613
rect 419395 165548 419396 165612
rect 419460 165548 419461 165612
rect 419395 165547 419461 165548
rect 417003 164252 417069 164253
rect 417003 164188 417004 164252
rect 417068 164188 417069 164252
rect 417003 164187 417069 164188
rect 418291 164252 418357 164253
rect 418291 164188 418292 164252
rect 418356 164188 418357 164252
rect 418291 164187 418357 164188
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 165000
rect 420686 164253 420746 166950
rect 421054 166950 421140 167010
rect 421760 167010 421820 167106
rect 422848 167010 422908 167106
rect 423528 167010 423588 167106
rect 423936 167010 423996 167106
rect 425296 167010 425356 167106
rect 421760 166950 421850 167010
rect 422848 166950 422954 167010
rect 421054 166837 421114 166950
rect 421051 166836 421117 166837
rect 421051 166772 421052 166836
rect 421116 166772 421117 166836
rect 421051 166771 421117 166772
rect 421790 164797 421850 166950
rect 421787 164796 421853 164797
rect 421787 164732 421788 164796
rect 421852 164732 421853 164796
rect 421787 164731 421853 164732
rect 422894 164253 422954 166950
rect 423446 166950 423588 167010
rect 423814 166950 423996 167010
rect 425286 166950 425356 167010
rect 425976 167010 426036 167106
rect 426384 167010 426444 167106
rect 427608 167010 427668 167106
rect 428288 167010 428348 167106
rect 425976 166950 426082 167010
rect 426384 166950 426450 167010
rect 427608 166950 427738 167010
rect 423446 166837 423506 166950
rect 423443 166836 423509 166837
rect 423443 166772 423444 166836
rect 423508 166772 423509 166836
rect 423443 166771 423509 166772
rect 423814 165613 423874 166950
rect 423811 165612 423877 165613
rect 423811 165548 423812 165612
rect 423876 165548 423877 165612
rect 423811 165547 423877 165548
rect 420683 164252 420749 164253
rect 420683 164188 420684 164252
rect 420748 164188 420749 164252
rect 420683 164187 420749 164188
rect 422891 164252 422957 164253
rect 422891 164188 422892 164252
rect 422956 164188 422957 164252
rect 422891 164187 422957 164188
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 155834 423854 165000
rect 425286 164253 425346 166950
rect 426022 165069 426082 166950
rect 426390 165613 426450 166950
rect 426387 165612 426453 165613
rect 426387 165548 426388 165612
rect 426452 165548 426453 165612
rect 426387 165547 426453 165548
rect 426019 165068 426085 165069
rect 426019 165004 426020 165068
rect 426084 165004 426085 165068
rect 426019 165003 426085 165004
rect 425283 164252 425349 164253
rect 425283 164188 425284 164252
rect 425348 164188 425349 164252
rect 425283 164187 425349 164188
rect 423234 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 423854 155834
rect 423234 155514 423854 155598
rect 423234 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 423854 155514
rect 423234 145308 423854 155278
rect 426954 157674 427574 165000
rect 427678 164253 427738 166950
rect 428230 166950 428348 167010
rect 428696 167010 428756 167106
rect 429784 167010 429844 167106
rect 431008 167010 431068 167106
rect 428696 166950 428842 167010
rect 428230 166293 428290 166950
rect 428227 166292 428293 166293
rect 428227 166228 428228 166292
rect 428292 166228 428293 166292
rect 428227 166227 428293 166228
rect 428782 164253 428842 166950
rect 429702 166950 429844 167010
rect 430990 166950 431068 167010
rect 431144 167010 431204 167106
rect 432232 167010 432292 167106
rect 433320 167010 433380 167106
rect 433592 167010 433652 167106
rect 434408 167010 434468 167106
rect 431144 166950 431234 167010
rect 432232 166950 432338 167010
rect 433320 166950 433442 167010
rect 429702 164389 429762 166950
rect 430990 166293 431050 166950
rect 430987 166292 431053 166293
rect 430987 166228 430988 166292
rect 431052 166228 431053 166292
rect 430987 166227 431053 166228
rect 429699 164388 429765 164389
rect 429699 164324 429700 164388
rect 429764 164324 429765 164388
rect 429699 164323 429765 164324
rect 431174 164253 431234 166950
rect 432278 164253 432338 166950
rect 433382 165613 433442 166950
rect 433566 166950 433652 167010
rect 434302 166950 434468 167010
rect 435768 167010 435828 167106
rect 436040 167010 436100 167106
rect 436992 167010 437052 167106
rect 438080 167010 438140 167106
rect 435768 166950 435834 167010
rect 433379 165612 433445 165613
rect 433379 165548 433380 165612
rect 433444 165548 433445 165612
rect 433379 165547 433445 165548
rect 433566 165069 433626 166950
rect 434302 165613 434362 166950
rect 434299 165612 434365 165613
rect 434299 165548 434300 165612
rect 434364 165548 434365 165612
rect 434299 165547 434365 165548
rect 433563 165068 433629 165069
rect 433563 165004 433564 165068
rect 433628 165004 433629 165068
rect 433563 165003 433629 165004
rect 427675 164252 427741 164253
rect 427675 164188 427676 164252
rect 427740 164188 427741 164252
rect 427675 164187 427741 164188
rect 428779 164252 428845 164253
rect 428779 164188 428780 164252
rect 428844 164188 428845 164252
rect 428779 164187 428845 164188
rect 431171 164252 431237 164253
rect 431171 164188 431172 164252
rect 431236 164188 431237 164252
rect 431171 164187 431237 164188
rect 432275 164252 432341 164253
rect 432275 164188 432276 164252
rect 432340 164188 432341 164252
rect 432275 164187 432341 164188
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 165000
rect 435774 164253 435834 166950
rect 435958 166950 436100 167010
rect 436878 166950 437052 167010
rect 437798 166950 438140 167010
rect 438488 167010 438548 167106
rect 439168 167010 439228 167106
rect 440936 167010 440996 167106
rect 443520 167010 443580 167106
rect 445968 167010 446028 167106
rect 438488 166950 438594 167010
rect 439168 166950 439330 167010
rect 435958 165613 436018 166950
rect 435955 165612 436021 165613
rect 435955 165548 435956 165612
rect 436020 165548 436021 165612
rect 435955 165547 436021 165548
rect 436878 164525 436938 166950
rect 437798 165613 437858 166950
rect 438534 165613 438594 166950
rect 437795 165612 437861 165613
rect 437795 165548 437796 165612
rect 437860 165548 437861 165612
rect 437795 165547 437861 165548
rect 438531 165612 438597 165613
rect 438531 165548 438532 165612
rect 438596 165548 438597 165612
rect 438531 165547 438597 165548
rect 436875 164524 436941 164525
rect 436875 164460 436876 164524
rect 436940 164460 436941 164524
rect 436875 164459 436941 164460
rect 435771 164252 435837 164253
rect 435771 164188 435772 164252
rect 435836 164188 435837 164252
rect 435771 164187 435837 164188
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 165000
rect 439270 164253 439330 166950
rect 440926 166950 440996 167010
rect 443502 166950 443580 167010
rect 445894 166950 446028 167010
rect 448280 167010 448340 167106
rect 451000 167010 451060 167106
rect 453448 167010 453508 167106
rect 455896 167010 455956 167106
rect 448280 166950 448346 167010
rect 451000 166950 451106 167010
rect 440926 164933 440986 166950
rect 443502 165613 443562 166950
rect 445894 166837 445954 166950
rect 445891 166836 445957 166837
rect 445891 166772 445892 166836
rect 445956 166772 445957 166836
rect 445891 166771 445957 166772
rect 448286 165613 448346 166950
rect 451046 165613 451106 166950
rect 453438 166950 453508 167010
rect 455830 166950 455956 167010
rect 453438 165613 453498 166950
rect 455830 165613 455890 166950
rect 458480 166290 458540 167106
rect 458406 166230 458540 166290
rect 460928 166290 460988 167106
rect 463512 166290 463572 167106
rect 465960 166290 466020 167106
rect 468544 166290 468604 167106
rect 470992 166837 471052 167106
rect 473440 166837 473500 167106
rect 475888 166837 475948 167106
rect 478472 166837 478532 167106
rect 480920 166837 480980 167106
rect 470989 166836 471055 166837
rect 470989 166772 470990 166836
rect 471054 166772 471055 166836
rect 470989 166771 471055 166772
rect 473437 166836 473503 166837
rect 473437 166772 473438 166836
rect 473502 166772 473503 166836
rect 473437 166771 473503 166772
rect 475885 166836 475951 166837
rect 475885 166772 475886 166836
rect 475950 166772 475951 166836
rect 475885 166771 475951 166772
rect 478469 166836 478535 166837
rect 478469 166772 478470 166836
rect 478534 166772 478535 166836
rect 478469 166771 478535 166772
rect 480917 166836 480983 166837
rect 480917 166772 480918 166836
rect 480982 166772 480983 166836
rect 480917 166771 480983 166772
rect 483368 166701 483428 167106
rect 485952 166701 486012 167106
rect 483365 166700 483431 166701
rect 483365 166636 483366 166700
rect 483430 166636 483431 166700
rect 483365 166635 483431 166636
rect 485949 166700 486015 166701
rect 485949 166636 485950 166700
rect 486014 166636 486015 166700
rect 485949 166635 486015 166636
rect 503224 166565 503284 167106
rect 503221 166564 503287 166565
rect 503221 166500 503222 166564
rect 503286 166500 503287 166564
rect 503221 166499 503287 166500
rect 503360 166290 503420 167106
rect 460928 166230 461042 166290
rect 463512 166230 463618 166290
rect 458406 165613 458466 166230
rect 443499 165612 443565 165613
rect 443499 165548 443500 165612
rect 443564 165548 443565 165612
rect 443499 165547 443565 165548
rect 448283 165612 448349 165613
rect 448283 165548 448284 165612
rect 448348 165548 448349 165612
rect 448283 165547 448349 165548
rect 451043 165612 451109 165613
rect 451043 165548 451044 165612
rect 451108 165548 451109 165612
rect 451043 165547 451109 165548
rect 453435 165612 453501 165613
rect 453435 165548 453436 165612
rect 453500 165548 453501 165612
rect 453435 165547 453501 165548
rect 455827 165612 455893 165613
rect 455827 165548 455828 165612
rect 455892 165548 455893 165612
rect 455827 165547 455893 165548
rect 458403 165612 458469 165613
rect 458403 165548 458404 165612
rect 458468 165548 458469 165612
rect 458403 165547 458469 165548
rect 440923 164932 440989 164933
rect 440923 164868 440924 164932
rect 440988 164868 440989 164932
rect 440923 164867 440989 164868
rect 439267 164252 439333 164253
rect 439267 164188 439268 164252
rect 439332 164188 439333 164252
rect 439267 164187 439333 164188
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 165000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 165000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 165000
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 165000
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 155834 459854 165000
rect 460982 164661 461042 166230
rect 463558 165205 463618 166230
rect 465950 166230 466020 166290
rect 468526 166230 468604 166290
rect 503302 166230 503420 166290
rect 465950 165341 466010 166230
rect 468526 165477 468586 166230
rect 503302 165613 503362 166230
rect 503299 165612 503365 165613
rect 503299 165548 503300 165612
rect 503364 165548 503365 165612
rect 503299 165547 503365 165548
rect 468523 165476 468589 165477
rect 468523 165412 468524 165476
rect 468588 165412 468589 165476
rect 468523 165411 468589 165412
rect 523794 165454 524414 200898
rect 465947 165340 466013 165341
rect 465947 165276 465948 165340
rect 466012 165276 466013 165340
rect 465947 165275 466013 165276
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 463555 165204 463621 165205
rect 463555 165140 463556 165204
rect 463620 165140 463621 165204
rect 463555 165139 463621 165140
rect 523794 165134 524414 165218
rect 460979 164660 461045 164661
rect 460979 164596 460980 164660
rect 461044 164596 461045 164660
rect 460979 164595 461045 164596
rect 459234 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 459854 155834
rect 459234 155514 459854 155598
rect 459234 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 459854 155514
rect 459234 145308 459854 155278
rect 462954 157674 463574 165000
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 165000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 165000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 165000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 165000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 165000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 165000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 155834 495854 165000
rect 495234 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 495234 155514 495854 155598
rect 495234 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 495234 145308 495854 155278
rect 498954 157674 499574 165000
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 165000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 165000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 165000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 145484 510909 145485
rect 510843 145420 510844 145484
rect 510908 145420 510909 145484
rect 510843 145419 510909 145420
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 145419
rect 513234 145308 513854 154338
rect 516954 158614 517574 165000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 397141 59739 397207 59740
rect 398232 59530 398292 60106
rect 399592 59666 399652 60106
rect 400544 59666 400604 60106
rect 399526 59606 399652 59666
rect 400446 59606 400604 59666
rect 398232 59470 398298 59530
rect 398238 58173 398298 59470
rect 398235 58172 398301 58173
rect 398235 58108 398236 58172
rect 398300 58108 398301 58172
rect 398235 58107 398301 58108
rect 379794 57454 380414 58000
rect 379283 57220 379349 57221
rect 379283 57156 379284 57220
rect 379348 57156 379349 57220
rect 379283 57155 379349 57156
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 378915 57084 378981 57085
rect 378915 57020 378916 57084
rect 378980 57020 378981 57084
rect 378915 57019 378981 57020
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 377811 55180 377877 55181
rect 377811 55116 377812 55180
rect 377876 55116 377877 55180
rect 377811 55115 377877 55116
rect 377627 55044 377693 55045
rect 377627 54980 377628 55044
rect 377692 54980 377693 55044
rect 377627 54979 377693 54980
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 375971 3500 376037 3501
rect 375971 3436 375972 3500
rect 376036 3436 376037 3500
rect 375971 3435 376037 3436
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59606
rect 400446 57901 400506 59606
rect 401768 59530 401828 60106
rect 403128 59669 403188 60106
rect 404216 59669 404276 60106
rect 403125 59668 403191 59669
rect 403125 59604 403126 59668
rect 403190 59604 403191 59668
rect 403125 59603 403191 59604
rect 404213 59668 404279 59669
rect 404213 59604 404214 59668
rect 404278 59604 404279 59668
rect 404213 59603 404279 59604
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 405414 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 405414 58173 405474 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 405411 58172 405477 58173
rect 405411 58108 405412 58172
rect 405476 58108 405477 58172
rect 405411 58107 405477 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59530 410804 60106
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59669 413524 60106
rect 413461 59668 413527 59669
rect 413461 59604 413462 59668
rect 413526 59604 413527 59668
rect 413461 59603 413527 59604
rect 413600 59530 413660 60106
rect 410744 59470 410810 59530
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410750 58445 410810 59470
rect 410747 58444 410813 58445
rect 410747 58380 410748 58444
rect 410812 58380 410813 58444
rect 410747 58379 410813 58380
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 59470 413660 59530
rect 414552 59530 414612 60106
rect 415912 59530 415972 60106
rect 416048 59805 416108 60106
rect 417000 59805 417060 60106
rect 416045 59804 416111 59805
rect 416045 59740 416046 59804
rect 416110 59740 416111 59804
rect 416045 59739 416111 59740
rect 416997 59804 417063 59805
rect 416997 59740 416998 59804
rect 417062 59740 417063 59804
rect 416997 59739 417063 59740
rect 414552 59470 414674 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413510 57085 413570 59470
rect 414614 57901 414674 59470
rect 415534 59470 415972 59530
rect 418088 59530 418148 60106
rect 418496 59530 418556 60106
rect 419448 59530 419508 60106
rect 418088 59470 418170 59530
rect 415534 57901 415594 59470
rect 418110 59397 418170 59470
rect 418478 59470 418556 59530
rect 419398 59470 419508 59530
rect 420672 59530 420732 60106
rect 421080 59530 421140 60106
rect 420672 59470 420746 59530
rect 418107 59396 418173 59397
rect 418107 59332 418108 59396
rect 418172 59332 418173 59396
rect 418107 59331 418173 59332
rect 414611 57900 414677 57901
rect 414611 57836 414612 57900
rect 414676 57836 414677 57900
rect 414611 57835 414677 57836
rect 415531 57900 415597 57901
rect 415531 57836 415532 57900
rect 415596 57836 415597 57900
rect 415531 57835 415597 57836
rect 415794 57454 416414 58000
rect 418478 57901 418538 59470
rect 419398 59397 419458 59470
rect 420686 59397 420746 59470
rect 421054 59470 421140 59530
rect 421760 59530 421820 60106
rect 422848 59805 422908 60106
rect 422845 59804 422911 59805
rect 422845 59740 422846 59804
rect 422910 59740 422911 59804
rect 422845 59739 422911 59740
rect 423528 59669 423588 60106
rect 423936 59805 423996 60106
rect 423933 59804 423999 59805
rect 423933 59740 423934 59804
rect 423998 59740 423999 59804
rect 423933 59739 423999 59740
rect 423525 59668 423591 59669
rect 423525 59604 423526 59668
rect 423590 59604 423591 59668
rect 423525 59603 423591 59604
rect 425296 59530 425356 60106
rect 421760 59470 421850 59530
rect 419395 59396 419461 59397
rect 419395 59332 419396 59396
rect 419460 59332 419461 59396
rect 419395 59331 419461 59332
rect 420683 59396 420749 59397
rect 420683 59332 420684 59396
rect 420748 59332 420749 59396
rect 420683 59331 420749 59332
rect 418475 57900 418541 57901
rect 418475 57836 418476 57900
rect 418540 57836 418541 57900
rect 418475 57835 418541 57836
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 413507 57084 413573 57085
rect 413507 57020 413508 57084
rect 413572 57020 413573 57084
rect 413507 57019 413573 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 421054 56541 421114 59470
rect 421790 59397 421850 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 421787 59396 421853 59397
rect 421787 59332 421788 59396
rect 421852 59332 421853 59396
rect 421787 59331 421853 59332
rect 421051 56540 421117 56541
rect 421051 56476 421052 56540
rect 421116 56476 421117 56540
rect 421051 56475 421117 56476
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 425286 57901 425346 59470
rect 426022 59397 426082 59470
rect 426019 59396 426085 59397
rect 426019 59332 426020 59396
rect 426084 59332 426085 59396
rect 426019 59331 426085 59332
rect 426390 57901 426450 59470
rect 425283 57900 425349 57901
rect 425283 57836 425284 57900
rect 425348 57836 425349 57900
rect 425283 57835 425349 57836
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57901 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 427675 57900 427741 57901
rect 427675 57836 427676 57900
rect 427740 57836 427741 57900
rect 427675 57835 427741 57836
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430990 57221 431050 59470
rect 431174 57901 431234 59470
rect 432278 57901 432338 59470
rect 433382 57901 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433566 57901 433626 59470
rect 431171 57900 431237 57901
rect 431171 57836 431172 57900
rect 431236 57836 431237 57900
rect 431171 57835 431237 57836
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433379 57900 433445 57901
rect 433379 57836 433380 57900
rect 433444 57836 433445 57900
rect 433379 57835 433445 57836
rect 433563 57900 433629 57901
rect 433563 57836 433564 57900
rect 433628 57836 433629 57900
rect 433563 57835 433629 57836
rect 430987 57220 431053 57221
rect 430987 57156 430988 57220
rect 431052 57156 431053 57220
rect 430987 57155 431053 57156
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57629 434730 59470
rect 435774 57901 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 435771 57900 435837 57901
rect 435771 57836 435772 57900
rect 435836 57836 435837 57900
rect 435771 57835 435837 57836
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436878 57629 436938 59470
rect 434667 57628 434733 57629
rect 434667 57564 434668 57628
rect 434732 57564 434733 57628
rect 434667 57563 434733 57564
rect 436875 57628 436941 57629
rect 436875 57564 436876 57628
rect 436940 57564 436941 57628
rect 436875 57563 436941 57564
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 56405 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 439086 57629 439146 59470
rect 439083 57628 439149 57629
rect 439083 57564 439084 57628
rect 439148 57564 439149 57628
rect 439083 57563 439149 57564
rect 440926 57221 440986 59470
rect 440923 57220 440989 57221
rect 440923 57156 440924 57220
rect 440988 57156 440989 57220
rect 440923 57155 440989 57156
rect 438347 56404 438413 56405
rect 438347 56340 438348 56404
rect 438412 56340 438413 56404
rect 438347 56339 438413 56340
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 57901 443562 59470
rect 443499 57900 443565 57901
rect 443499 57836 443500 57900
rect 443564 57836 443565 57900
rect 443499 57835 443565 57836
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57901 445954 59470
rect 448286 57901 448346 59470
rect 445891 57900 445957 57901
rect 445891 57836 445892 57900
rect 445956 57836 445957 57900
rect 445891 57835 445957 57836
rect 448283 57900 448349 57901
rect 448283 57836 448284 57900
rect 448348 57836 448349 57900
rect 448283 57835 448349 57836
rect 451046 57357 451106 59470
rect 453438 59470 453508 59530
rect 455896 59530 455956 60106
rect 458480 59530 458540 60106
rect 455896 59470 456442 59530
rect 453438 59397 453498 59470
rect 453435 59396 453501 59397
rect 453435 59332 453436 59396
rect 453500 59332 453501 59396
rect 453435 59331 453501 59332
rect 451794 57454 452414 58000
rect 451043 57356 451109 57357
rect 451043 57292 451044 57356
rect 451108 57292 451109 57356
rect 451043 57291 451109 57292
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 456382 57493 456442 59470
rect 458406 59470 458540 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 458406 58581 458466 59470
rect 458403 58580 458469 58581
rect 458403 58516 458404 58580
rect 458468 58516 458469 58580
rect 458403 58515 458469 58516
rect 456379 57492 456445 57493
rect 456379 57428 456380 57492
rect 456444 57428 456445 57492
rect 456379 57427 456445 57428
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 56677 461042 59470
rect 463558 58717 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59530 480980 60106
rect 473440 59470 473554 59530
rect 463555 58716 463621 58717
rect 463555 58652 463556 58716
rect 463620 58652 463621 58716
rect 463555 58651 463621 58652
rect 460979 56676 461045 56677
rect 460979 56612 460980 56676
rect 461044 56612 461045 56676
rect 460979 56611 461045 56612
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 465950 57901 466010 59470
rect 468526 58989 468586 59470
rect 468523 58988 468589 58989
rect 468523 58924 468524 58988
rect 468588 58924 468589 58988
rect 468523 58923 468589 58924
rect 465947 57900 466013 57901
rect 465947 57836 465948 57900
rect 466012 57836 466013 57900
rect 465947 57835 466013 57836
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 470918 57765 470978 59470
rect 473494 58853 473554 59470
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 480854 59470 480980 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59530 503284 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 475886 58989 475946 59470
rect 475883 58988 475949 58989
rect 475883 58924 475884 58988
rect 475948 58924 475949 58988
rect 475883 58923 475949 58924
rect 473491 58852 473557 58853
rect 473491 58788 473492 58852
rect 473556 58788 473557 58852
rect 473491 58787 473557 58788
rect 470915 57764 470981 57765
rect 470915 57700 470916 57764
rect 470980 57700 470981 57764
rect 470915 57699 470981 57700
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 478462 57901 478522 59470
rect 480854 59125 480914 59470
rect 483430 59261 483490 59470
rect 483427 59260 483493 59261
rect 483427 59196 483428 59260
rect 483492 59196 483493 59260
rect 483427 59195 483493 59196
rect 480851 59124 480917 59125
rect 480851 59060 480852 59124
rect 480916 59060 480917 59124
rect 480851 59059 480917 59060
rect 478459 57900 478525 57901
rect 478459 57836 478460 57900
rect 478524 57836 478525 57900
rect 478459 57835 478525 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 486006 57901 486066 59470
rect 503118 59470 503284 59530
rect 503360 59530 503420 60106
rect 503360 59470 503546 59530
rect 486003 57900 486069 57901
rect 486003 57836 486004 57900
rect 486068 57836 486069 57900
rect 486003 57835 486069 57836
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503118 57901 503178 59470
rect 503486 57901 503546 59470
rect 503115 57900 503181 57901
rect 503115 57836 503116 57900
rect 503180 57836 503181 57900
rect 503115 57835 503181 57836
rect 503483 57900 503549 57901
rect 503483 57836 503484 57900
rect 503548 57836 503549 57900
rect 503483 57835 503549 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 551598 63502 551834
rect 63586 551598 63822 551834
rect 63266 551278 63502 551514
rect 63586 551278 63822 551514
rect 66986 555318 67222 555554
rect 67306 555318 67542 555554
rect 66986 554998 67222 555234
rect 67306 554998 67542 555234
rect 73826 560278 74062 560514
rect 74146 560278 74382 560514
rect 73826 559958 74062 560194
rect 74146 559958 74382 560194
rect 77546 563998 77782 564234
rect 77866 563998 78102 564234
rect 77546 563678 77782 563914
rect 77866 563678 78102 563914
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 551598 99502 551834
rect 99586 551598 99822 551834
rect 99266 551278 99502 551514
rect 99586 551278 99822 551514
rect 102986 555318 103222 555554
rect 103306 555318 103542 555554
rect 102986 554998 103222 555234
rect 103306 554998 103542 555234
rect 109826 560278 110062 560514
rect 110146 560278 110382 560514
rect 109826 559958 110062 560194
rect 110146 559958 110382 560194
rect 113546 563998 113782 564234
rect 113866 563998 114102 564234
rect 113546 563678 113782 563914
rect 113866 563678 114102 563914
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 144250 615218 144486 615454
rect 144250 614898 144486 615134
rect 174970 615218 175206 615454
rect 174970 614898 175206 615134
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 159610 597218 159846 597454
rect 159610 596898 159846 597134
rect 190330 597218 190566 597454
rect 190330 596898 190566 597134
rect 144250 579218 144486 579454
rect 144250 578898 144486 579134
rect 174970 579218 175206 579454
rect 174970 578898 175206 579134
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 551598 135502 551834
rect 135586 551598 135822 551834
rect 135266 551278 135502 551514
rect 135586 551278 135822 551514
rect 138986 555318 139222 555554
rect 139306 555318 139542 555554
rect 138986 554998 139222 555234
rect 139306 554998 139542 555234
rect 145826 560278 146062 560514
rect 146146 560278 146382 560514
rect 145826 559958 146062 560194
rect 146146 559958 146382 560194
rect 149546 563998 149782 564234
rect 149866 563998 150102 564234
rect 149546 563678 149782 563914
rect 149866 563678 150102 563914
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 551598 171502 551834
rect 171586 551598 171822 551834
rect 171266 551278 171502 551514
rect 171586 551278 171822 551514
rect 174986 555318 175222 555554
rect 175306 555318 175542 555554
rect 174986 554998 175222 555234
rect 175306 554998 175542 555234
rect 181826 560278 182062 560514
rect 182146 560278 182382 560514
rect 181826 559958 182062 560194
rect 182146 559958 182382 560194
rect 185546 563998 185782 564234
rect 185866 563998 186102 564234
rect 185546 563678 185782 563914
rect 185866 563678 186102 563914
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 551598 207502 551834
rect 207586 551598 207822 551834
rect 207266 551278 207502 551514
rect 207586 551278 207822 551514
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 224250 615218 224486 615454
rect 224250 614898 224486 615134
rect 254970 615218 255206 615454
rect 254970 614898 255206 615134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 239610 597218 239846 597454
rect 239610 596898 239846 597134
rect 270330 597218 270566 597454
rect 270330 596898 270566 597134
rect 224250 579218 224486 579454
rect 224250 578898 224486 579134
rect 254970 579218 255206 579454
rect 254970 578898 255206 579134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 555318 211222 555554
rect 211306 555318 211542 555554
rect 210986 554998 211222 555234
rect 211306 554998 211542 555234
rect 217826 560278 218062 560514
rect 218146 560278 218382 560514
rect 217826 559958 218062 560194
rect 218146 559958 218382 560194
rect 221546 563998 221782 564234
rect 221866 563998 222102 564234
rect 221546 563678 221782 563914
rect 221866 563678 222102 563914
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 551598 243502 551834
rect 243586 551598 243822 551834
rect 243266 551278 243502 551514
rect 243586 551278 243822 551514
rect 246986 555318 247222 555554
rect 247306 555318 247542 555554
rect 246986 554998 247222 555234
rect 247306 554998 247542 555234
rect 253826 560278 254062 560514
rect 254146 560278 254382 560514
rect 253826 559958 254062 560194
rect 254146 559958 254382 560194
rect 257546 563998 257782 564234
rect 257866 563998 258102 564234
rect 257546 563678 257782 563914
rect 257866 563678 258102 563914
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 551598 279502 551834
rect 279586 551598 279822 551834
rect 279266 551278 279502 551514
rect 279586 551278 279822 551514
rect 282986 555318 283222 555554
rect 283306 555318 283542 555554
rect 282986 554998 283222 555234
rect 283306 554998 283542 555234
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 64250 543218 64486 543454
rect 64250 542898 64486 543134
rect 94970 543218 95206 543454
rect 94970 542898 95206 543134
rect 125690 543218 125926 543454
rect 125690 542898 125926 543134
rect 156410 543218 156646 543454
rect 156410 542898 156646 543134
rect 187130 543218 187366 543454
rect 187130 542898 187366 543134
rect 217850 543218 218086 543454
rect 217850 542898 218086 543134
rect 248570 543218 248806 543454
rect 248570 542898 248806 543134
rect 279290 543218 279526 543454
rect 279290 542898 279526 543134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 475878 59782 476114
rect 59866 475878 60102 476114
rect 59546 475558 59782 475794
rect 59866 475558 60102 475794
rect 63266 477718 63502 477954
rect 63586 477718 63822 477954
rect 63266 477398 63502 477634
rect 63586 477398 63822 477634
rect 66986 481438 67222 481674
rect 67306 481438 67542 481674
rect 66986 481118 67222 481354
rect 67306 481118 67542 481354
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 472158 92062 472394
rect 92146 472158 92382 472394
rect 91826 471838 92062 472074
rect 92146 471838 92382 472074
rect 95546 475878 95782 476114
rect 95866 475878 96102 476114
rect 95546 475558 95782 475794
rect 95866 475558 96102 475794
rect 99266 477718 99502 477954
rect 99586 477718 99822 477954
rect 99266 477398 99502 477634
rect 99586 477398 99822 477634
rect 102986 481438 103222 481674
rect 103306 481438 103542 481674
rect 102986 481118 103222 481354
rect 103306 481118 103542 481354
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 472158 128062 472394
rect 128146 472158 128382 472394
rect 127826 471838 128062 472074
rect 128146 471838 128382 472074
rect 131546 475878 131782 476114
rect 131866 475878 132102 476114
rect 131546 475558 131782 475794
rect 131866 475558 132102 475794
rect 135266 477718 135502 477954
rect 135586 477718 135822 477954
rect 135266 477398 135502 477634
rect 135586 477398 135822 477634
rect 138986 481438 139222 481674
rect 139306 481438 139542 481674
rect 138986 481118 139222 481354
rect 139306 481118 139542 481354
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 472158 164062 472394
rect 164146 472158 164382 472394
rect 163826 471838 164062 472074
rect 164146 471838 164382 472074
rect 167546 475878 167782 476114
rect 167866 475878 168102 476114
rect 167546 475558 167782 475794
rect 167866 475558 168102 475794
rect 171266 477718 171502 477954
rect 171586 477718 171822 477954
rect 171266 477398 171502 477634
rect 171586 477398 171822 477634
rect 174986 481438 175222 481674
rect 175306 481438 175542 481674
rect 174986 481118 175222 481354
rect 175306 481118 175542 481354
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 59546 367878 59782 368114
rect 59866 367878 60102 368114
rect 59546 367558 59782 367794
rect 59866 367558 60102 367794
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 373438 67222 373674
rect 67306 373438 67542 373674
rect 66986 373118 67222 373354
rect 67306 373118 67542 373354
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 367878 95782 368114
rect 95866 367878 96102 368114
rect 95546 367558 95782 367794
rect 95866 367558 96102 367794
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 373438 103222 373674
rect 103306 373438 103542 373674
rect 102986 373118 103222 373354
rect 103306 373118 103542 373354
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 367878 131782 368114
rect 131866 367878 132102 368114
rect 131546 367558 131782 367794
rect 131866 367558 132102 367794
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 373438 139222 373674
rect 139306 373438 139542 373674
rect 138986 373118 139222 373354
rect 139306 373118 139542 373354
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 367878 167782 368114
rect 167866 367878 168102 368114
rect 167546 367558 167782 367794
rect 167866 367558 168102 367794
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 373438 175222 373674
rect 175306 373438 175542 373674
rect 174986 373118 175222 373354
rect 175306 373118 175542 373354
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 155598 63502 155834
rect 63586 155598 63822 155834
rect 63266 155278 63502 155514
rect 63586 155278 63822 155514
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 155598 99502 155834
rect 99586 155598 99822 155834
rect 99266 155278 99502 155514
rect 99586 155278 99822 155514
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 155598 135502 155834
rect 135586 155598 135822 155834
rect 135266 155278 135502 155514
rect 135586 155278 135822 155514
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 155598 171502 155834
rect 171586 155598 171822 155834
rect 171266 155278 171502 155514
rect 171586 155278 171822 155514
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 199826 472158 200062 472394
rect 200146 472158 200382 472394
rect 199826 471838 200062 472074
rect 200146 471838 200382 472074
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 203546 475878 203782 476114
rect 203866 475878 204102 476114
rect 203546 475558 203782 475794
rect 203866 475558 204102 475794
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 367878 203782 368114
rect 203866 367878 204102 368114
rect 203546 367558 203782 367794
rect 203866 367558 204102 367794
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 207266 477718 207502 477954
rect 207586 477718 207822 477954
rect 207266 477398 207502 477634
rect 207586 477398 207822 477634
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 155598 207502 155834
rect 207586 155598 207822 155834
rect 207266 155278 207502 155514
rect 207586 155278 207822 155514
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 210986 481438 211222 481674
rect 211306 481438 211542 481674
rect 210986 481118 211222 481354
rect 211306 481118 211542 481354
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 373438 211222 373674
rect 211306 373438 211542 373674
rect 210986 373118 211222 373354
rect 211306 373118 211542 373354
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 472158 236062 472394
rect 236146 472158 236382 472394
rect 235826 471838 236062 472074
rect 236146 471838 236382 472074
rect 239546 475878 239782 476114
rect 239866 475878 240102 476114
rect 239546 475558 239782 475794
rect 239866 475558 240102 475794
rect 243266 477718 243502 477954
rect 243586 477718 243822 477954
rect 243266 477398 243502 477634
rect 243586 477398 243822 477634
rect 246986 481438 247222 481674
rect 247306 481438 247542 481674
rect 246986 481118 247222 481354
rect 247306 481118 247542 481354
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 472158 272062 472394
rect 272146 472158 272382 472394
rect 271826 471838 272062 472074
rect 272146 471838 272382 472074
rect 275546 475878 275782 476114
rect 275866 475878 276102 476114
rect 275546 475558 275782 475794
rect 275866 475558 276102 475794
rect 279266 477718 279502 477954
rect 279586 477718 279822 477954
rect 279266 477398 279502 477634
rect 279586 477398 279822 477634
rect 282986 481438 283222 481674
rect 283306 481438 283542 481674
rect 282986 481118 283222 481354
rect 283306 481118 283542 481354
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 339610 633218 339846 633454
rect 339610 632898 339846 633134
rect 370330 633218 370566 633454
rect 370330 632898 370566 633134
rect 401050 633218 401286 633454
rect 401050 632898 401286 633134
rect 324250 615218 324486 615454
rect 324250 614898 324486 615134
rect 354970 615218 355206 615454
rect 354970 614898 355206 615134
rect 385690 615218 385926 615454
rect 385690 614898 385926 615134
rect 416410 615218 416646 615454
rect 416410 614898 416646 615134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 339610 597218 339846 597454
rect 339610 596898 339846 597134
rect 370330 597218 370566 597454
rect 370330 596898 370566 597134
rect 401050 597218 401286 597454
rect 401050 596898 401286 597134
rect 324250 579218 324486 579454
rect 324250 578898 324486 579134
rect 354970 579218 355206 579454
rect 354970 578898 355206 579134
rect 385690 579218 385926 579454
rect 385690 578898 385926 579134
rect 416410 579218 416646 579454
rect 416410 578898 416646 579134
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 339610 561218 339846 561454
rect 339610 560898 339846 561134
rect 370330 561218 370566 561454
rect 370330 560898 370566 561134
rect 401050 561218 401286 561454
rect 401050 560898 401286 561134
rect 324250 543218 324486 543454
rect 324250 542898 324486 543134
rect 354970 543218 355206 543454
rect 354970 542898 355206 543134
rect 385690 543218 385926 543454
rect 385690 542898 385926 543134
rect 416410 543218 416646 543454
rect 416410 542898 416646 543134
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 367878 239782 368114
rect 239866 367878 240102 368114
rect 239546 367558 239782 367794
rect 239866 367558 240102 367794
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 373438 247222 373674
rect 247306 373438 247542 373674
rect 246986 373118 247222 373354
rect 247306 373118 247542 373354
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 367878 275782 368114
rect 275866 367878 276102 368114
rect 275546 367558 275782 367794
rect 275866 367558 276102 367794
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 373438 283222 373674
rect 283306 373438 283542 373674
rect 282986 373118 283222 373354
rect 283306 373118 283542 373354
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 367878 311782 368114
rect 311866 367878 312102 368114
rect 311546 367558 311782 367794
rect 311866 367558 312102 367794
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 373438 319222 373674
rect 319306 373438 319542 373674
rect 318986 373118 319222 373354
rect 319306 373118 319542 373354
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 367878 347782 368114
rect 347866 367878 348102 368114
rect 347546 367558 347782 367794
rect 347866 367558 348102 367794
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 373438 355222 373674
rect 355306 373438 355542 373674
rect 354986 373118 355222 373354
rect 355306 373118 355542 373354
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 155598 243502 155834
rect 243586 155598 243822 155834
rect 243266 155278 243502 155514
rect 243586 155278 243822 155514
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 155598 279502 155834
rect 279586 155598 279822 155834
rect 279266 155278 279502 155514
rect 279586 155278 279822 155514
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 155598 315502 155834
rect 315586 155598 315822 155834
rect 315266 155278 315502 155514
rect 315586 155278 315822 155514
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 155598 351502 155834
rect 351586 155598 351822 155834
rect 351266 155278 351502 155514
rect 351586 155278 351822 155514
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 367878 383782 368114
rect 383866 367878 384102 368114
rect 383546 367558 383782 367794
rect 383866 367558 384102 367794
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 373438 391222 373674
rect 391306 373438 391542 373674
rect 390986 373118 391222 373354
rect 391306 373118 391542 373354
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 367878 419782 368114
rect 419866 367878 420102 368114
rect 419546 367558 419782 367794
rect 419866 367558 420102 367794
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 373438 427222 373674
rect 427306 373438 427542 373674
rect 426986 373118 427222 373354
rect 427306 373118 427542 373354
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 367878 455782 368114
rect 455866 367878 456102 368114
rect 455546 367558 455782 367794
rect 455866 367558 456102 367794
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 373438 463222 373674
rect 463306 373438 463542 373674
rect 462986 373118 463222 373354
rect 463306 373118 463542 373354
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 367878 491782 368114
rect 491866 367878 492102 368114
rect 491546 367558 491782 367794
rect 491866 367558 492102 367794
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 373438 499222 373674
rect 499306 373438 499542 373674
rect 498986 373118 499222 373354
rect 499306 373118 499542 373354
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 155598 387502 155834
rect 387586 155598 387822 155834
rect 387266 155278 387502 155514
rect 387586 155278 387822 155514
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 155598 423502 155834
rect 423586 155598 423822 155834
rect 423266 155278 423502 155514
rect 423586 155278 423822 155514
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 459266 155598 459502 155834
rect 459586 155598 459822 155834
rect 459266 155278 459502 155514
rect 459586 155278 459822 155514
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 155598 495502 155834
rect 495586 155598 495822 155834
rect 495266 155278 495502 155514
rect 495586 155278 495822 155514
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 339610 633454
rect 339846 633218 370330 633454
rect 370566 633218 401050 633454
rect 401286 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 339610 633134
rect 339846 632898 370330 633134
rect 370566 632898 401050 633134
rect 401286 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 144250 615454
rect 144486 615218 174970 615454
rect 175206 615218 224250 615454
rect 224486 615218 254970 615454
rect 255206 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 324250 615454
rect 324486 615218 354970 615454
rect 355206 615218 385690 615454
rect 385926 615218 416410 615454
rect 416646 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 144250 615134
rect 144486 614898 174970 615134
rect 175206 614898 224250 615134
rect 224486 614898 254970 615134
rect 255206 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 324250 615134
rect 324486 614898 354970 615134
rect 355206 614898 385690 615134
rect 385926 614898 416410 615134
rect 416646 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 159610 597454
rect 159846 597218 190330 597454
rect 190566 597218 239610 597454
rect 239846 597218 270330 597454
rect 270566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 339610 597454
rect 339846 597218 370330 597454
rect 370566 597218 401050 597454
rect 401286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 159610 597134
rect 159846 596898 190330 597134
rect 190566 596898 239610 597134
rect 239846 596898 270330 597134
rect 270566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 339610 597134
rect 339846 596898 370330 597134
rect 370566 596898 401050 597134
rect 401286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 144250 579454
rect 144486 579218 174970 579454
rect 175206 579218 224250 579454
rect 224486 579218 254970 579454
rect 255206 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 324250 579454
rect 324486 579218 354970 579454
rect 355206 579218 385690 579454
rect 385926 579218 416410 579454
rect 416646 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 144250 579134
rect 144486 578898 174970 579134
rect 175206 578898 224250 579134
rect 224486 578898 254970 579134
rect 255206 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 324250 579134
rect 324486 578898 354970 579134
rect 355206 578898 385690 579134
rect 385926 578898 416410 579134
rect 416646 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect 77514 564234 258134 564266
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 258134 564234
rect 77514 563914 258134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 258134 563914
rect 77514 563646 258134 563678
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 339610 561454
rect 339846 561218 370330 561454
rect 370566 561218 401050 561454
rect 401286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 339610 561134
rect 339846 560898 370330 561134
rect 370566 560898 401050 561134
rect 401286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect 73794 560514 254414 560546
rect 73794 560278 73826 560514
rect 74062 560278 74146 560514
rect 74382 560278 109826 560514
rect 110062 560278 110146 560514
rect 110382 560278 145826 560514
rect 146062 560278 146146 560514
rect 146382 560278 181826 560514
rect 182062 560278 182146 560514
rect 182382 560278 217826 560514
rect 218062 560278 218146 560514
rect 218382 560278 253826 560514
rect 254062 560278 254146 560514
rect 254382 560278 254414 560514
rect 73794 560194 254414 560278
rect 73794 559958 73826 560194
rect 74062 559958 74146 560194
rect 74382 559958 109826 560194
rect 110062 559958 110146 560194
rect 110382 559958 145826 560194
rect 146062 559958 146146 560194
rect 146382 559958 181826 560194
rect 182062 559958 182146 560194
rect 182382 559958 217826 560194
rect 218062 559958 218146 560194
rect 218382 559958 253826 560194
rect 254062 559958 254146 560194
rect 254382 559958 254414 560194
rect 73794 559926 254414 559958
rect 66954 555554 283574 555586
rect 66954 555318 66986 555554
rect 67222 555318 67306 555554
rect 67542 555318 102986 555554
rect 103222 555318 103306 555554
rect 103542 555318 138986 555554
rect 139222 555318 139306 555554
rect 139542 555318 174986 555554
rect 175222 555318 175306 555554
rect 175542 555318 210986 555554
rect 211222 555318 211306 555554
rect 211542 555318 246986 555554
rect 247222 555318 247306 555554
rect 247542 555318 282986 555554
rect 283222 555318 283306 555554
rect 283542 555318 283574 555554
rect 66954 555234 283574 555318
rect 66954 554998 66986 555234
rect 67222 554998 67306 555234
rect 67542 554998 102986 555234
rect 103222 554998 103306 555234
rect 103542 554998 138986 555234
rect 139222 554998 139306 555234
rect 139542 554998 174986 555234
rect 175222 554998 175306 555234
rect 175542 554998 210986 555234
rect 211222 554998 211306 555234
rect 211542 554998 246986 555234
rect 247222 554998 247306 555234
rect 247542 554998 282986 555234
rect 283222 554998 283306 555234
rect 283542 554998 283574 555234
rect 66954 554966 283574 554998
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect 63234 551834 279854 551866
rect 63234 551598 63266 551834
rect 63502 551598 63586 551834
rect 63822 551598 99266 551834
rect 99502 551598 99586 551834
rect 99822 551598 135266 551834
rect 135502 551598 135586 551834
rect 135822 551598 171266 551834
rect 171502 551598 171586 551834
rect 171822 551598 207266 551834
rect 207502 551598 207586 551834
rect 207822 551598 243266 551834
rect 243502 551598 243586 551834
rect 243822 551598 279266 551834
rect 279502 551598 279586 551834
rect 279822 551598 279854 551834
rect 63234 551514 279854 551598
rect 63234 551278 63266 551514
rect 63502 551278 63586 551514
rect 63822 551278 99266 551514
rect 99502 551278 99586 551514
rect 99822 551278 135266 551514
rect 135502 551278 135586 551514
rect 135822 551278 171266 551514
rect 171502 551278 171586 551514
rect 171822 551278 207266 551514
rect 207502 551278 207586 551514
rect 207822 551278 243266 551514
rect 243502 551278 243586 551514
rect 243822 551278 279266 551514
rect 279502 551278 279586 551514
rect 279822 551278 279854 551514
rect 63234 551246 279854 551278
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64250 543454
rect 64486 543218 94970 543454
rect 95206 543218 125690 543454
rect 125926 543218 156410 543454
rect 156646 543218 187130 543454
rect 187366 543218 217850 543454
rect 218086 543218 248570 543454
rect 248806 543218 279290 543454
rect 279526 543218 324250 543454
rect 324486 543218 354970 543454
rect 355206 543218 385690 543454
rect 385926 543218 416410 543454
rect 416646 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64250 543134
rect 64486 542898 94970 543134
rect 95206 542898 125690 543134
rect 125926 542898 156410 543134
rect 156646 542898 187130 543134
rect 187366 542898 217850 543134
rect 218086 542898 248570 543134
rect 248806 542898 279290 543134
rect 279526 542898 324250 543134
rect 324486 542898 354970 543134
rect 355206 542898 385690 543134
rect 385926 542898 416410 543134
rect 416646 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect 66954 481674 283574 481706
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 66954 481354 283574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 66954 481086 283574 481118
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect 63234 477954 279854 477986
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 63234 477634 279854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 63234 477366 279854 477398
rect 59514 476114 276134 476146
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 59514 475794 276134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 59514 475526 276134 475558
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect 91794 472394 272414 472426
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 91794 472074 272414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 91794 471806 272414 471838
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect 66954 373674 499574 373706
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 66954 373354 499574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 66954 373086 499574 373118
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect 59514 368114 492134 368146
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 59514 367794 492134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 59514 367526 492134 367558
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect 63234 155834 495854 155866
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 63234 155514 495854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 63234 155246 495854 155278
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 381000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 568000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 220000 0 1 568000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 140000 0 1 568000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 488000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 320000 0 1 528000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 578000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s 73794 559926 254414 560546 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 252308 74414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 252308 110414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 252308 146414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 252308 182414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252308 218414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252308 254414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252308 290414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252308 326414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252308 398414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 252308 434414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 252308 470414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 252308 506414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 359308 74414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 359308 110414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 359308 146414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 359308 182414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 359308 218414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 359308 254414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 359308 290414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 359308 326414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 359308 398414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 359308 434414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 359308 470414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 359308 506414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 466308 74414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 466308 110414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 466308 146414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 466308 182414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 466308 218414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 466308 254414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 466308 290414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 466308 326414 526000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 526000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 466308 398414 526000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 550000 74414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 550000 110414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 550000 146414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 550000 182414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 550000 218414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 550000 254414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 466308 470414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 466308 506414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 633099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 633099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 633099 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 633099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 633099 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 633099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 550000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 641033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 641033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 641033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 466308 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 630000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 630000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s 77514 563646 258134 564266 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 252308 78134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 252308 114134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 252308 150134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 252308 186134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252308 222134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252308 258134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252308 294134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252308 330134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252308 402134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 252308 438134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 252308 474134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 252308 510134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 359308 78134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 359308 114134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 359308 150134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 359308 186134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 359308 222134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 359308 258134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 359308 294134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 359308 330134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 359308 402134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 359308 438134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 359308 474134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 359308 510134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 466308 78134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 466308 114134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 466308 150134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 466308 186134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 466308 222134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 466308 258134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 466308 294134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 466308 330134 526000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 526000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 466308 402134 526000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 550000 78134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 550000 114134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 550000 150134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 550000 186134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 550000 222134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 550000 258134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 466308 474134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 466308 510134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 633099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 633099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 633099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 633099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 633099 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 633099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 550000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 641033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 641033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 641033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 466308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 630000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 630000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 252308 81854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 252308 117854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 252308 153854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252308 189854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252308 225854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252308 261854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252308 297854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252308 333854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252308 405854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 252308 441854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 252308 477854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 252308 513854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 359308 81854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 359308 117854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 359308 153854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 359308 189854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 359308 225854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 359308 261854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 359308 297854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 359308 333854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 359308 405854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 359308 441854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 359308 477854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 359308 513854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 466308 81854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 466308 117854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 466308 153854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 466308 189854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 466308 225854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 466308 261854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 466308 297854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 466308 333854 526000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 526000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 466308 405854 526000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 550000 81854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 550000 117854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 550000 153854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 550000 189854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 550000 225854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 550000 261854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 466308 477854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 633099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 633099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 633099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 633099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 633099 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 633099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 550000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 641033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 641033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 641033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 466308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 630000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 466308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 252308 85574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 252308 121574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 252308 157574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252308 193574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252308 229574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252308 265574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252308 301574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252308 337574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252308 409574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 252308 445574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 252308 481574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 252308 517574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 359308 85574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 359308 121574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 359308 157574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 359308 193574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 359308 229574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 359308 265574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 359308 301574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 359308 337574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 359308 409574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 359308 445574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 359308 481574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 359308 517574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 466308 85574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 466308 121574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 466308 157574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 466308 193574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 466308 229574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 466308 265574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 466308 301574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 466308 337574 526000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 526000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 466308 409574 526000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 550000 85574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 550000 121574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 550000 157574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 550000 193574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 550000 229574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 550000 265574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 466308 481574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 633099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 633099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 633099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 633099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 633099 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 633099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 550000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 641033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 641033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 641033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 466308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 630000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 466308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 155246 495854 155866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 477366 279854 477986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 551246 279854 551866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 252308 63854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 252308 99854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 252308 135854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 252308 171854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252308 243854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252308 279854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252308 315854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252308 351854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252308 387854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 252308 423854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 252308 459854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 252308 495854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 359308 63854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 359308 99854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 359308 135854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 359308 171854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 359308 243854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 359308 279854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 359308 315854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 359308 351854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 359308 387854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 359308 423854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 359308 459854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 359308 495854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 466308 63854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 466308 99854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 466308 135854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 466308 171854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 466308 243854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 466308 279854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 466308 351854 526000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 466308 387854 526000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 466308 423854 526000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 550000 63854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 550000 99854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 550000 171854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 550000 243854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 550000 279854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 466308 459854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 466308 495854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 633099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 633099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 550000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 633099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 550000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 633099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 633099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 466308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 641033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 641033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 641033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 630000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 630000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 373086 499574 373706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 481086 283574 481706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 554966 283574 555586 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 252308 67574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 252308 103574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 252308 139574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 252308 175574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252308 247574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252308 283574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252308 319574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252308 355574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252308 391574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 252308 427574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 252308 463574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 252308 499574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 359308 67574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 359308 103574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 359308 139574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 359308 175574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 359308 247574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 359308 283574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 359308 319574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 359308 355574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 359308 391574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 359308 427574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 359308 463574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 359308 499574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 466308 67574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 466308 103574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 466308 139574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 466308 175574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 466308 247574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 466308 283574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 466308 319574 526000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 466308 355574 526000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 466308 391574 526000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 466308 427574 526000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 550000 67574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 550000 103574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 550000 139574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 550000 175574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 550000 247574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 550000 283574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 466308 463574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 466308 499574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 633099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 633099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 633099 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 633099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 550000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 633099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 633099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 641033 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 641033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 641033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 641033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 630000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 630000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 471806 272414 472426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 252308 92414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 252308 128414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 252308 164414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252308 236414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252308 272414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252308 308414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252308 344414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252308 380414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 252308 416414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 252308 452414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 252308 488414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 359308 92414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 359308 128414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 359308 164414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 359308 236414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 359308 272414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 359308 308414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 359308 344414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 359308 380414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 359308 416414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 359308 452414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 359308 488414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 466308 92414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 466308 128414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 466308 164414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 466308 236414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 466308 272414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 466308 344414 526000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 466308 380414 526000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 466308 416414 526000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 550000 92414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 550000 164414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 550000 200414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 550000 236414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 550000 272414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 466308 488414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 633099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 550000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 633099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 633099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 633099 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 633099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 466308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 641033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 641033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 641033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 466308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 630000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 367526 492134 368146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 252308 60134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 252308 96134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 252308 132134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 252308 168134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252308 240134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252308 276134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252308 312134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252308 348134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252308 384134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 252308 420134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 252308 456134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 252308 492134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 359308 60134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 359308 96134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 359308 132134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 359308 168134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 359308 240134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 359308 276134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 359308 312134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 359308 348134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 359308 384134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 359308 420134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 359308 456134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 359308 492134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 466308 60134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 466308 96134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 466308 132134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 466308 168134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 466308 240134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 466308 276134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 466308 348134 526000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 466308 384134 526000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 466308 420134 526000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 550000 60134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 550000 96134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 550000 168134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 550000 240134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 550000 276134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 466308 492134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 633099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 633099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 550000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 633099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 550000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 633099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 633099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 466308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 641033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 641033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 641033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 466308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 630000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
