magic
tech sky130A
magscale 1 2
timestamp 1655448201
<< metal1 >>
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 305638 700448 305644 700460
rect 235224 700420 305644 700448
rect 235224 700408 235230 700420
rect 305638 700408 305644 700420
rect 305696 700408 305702 700460
rect 429838 700408 429844 700460
rect 429896 700448 429902 700460
rect 434714 700448 434720 700460
rect 429896 700420 434720 700448
rect 429896 700408 429902 700420
rect 434714 700408 434720 700420
rect 434772 700408 434778 700460
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 434806 700380 434812 700392
rect 170364 700352 434812 700380
rect 170364 700340 170370 700352
rect 434806 700340 434812 700352
rect 434864 700340 434870 700392
rect 57698 700272 57704 700324
rect 57756 700312 57762 700324
rect 543458 700312 543464 700324
rect 57756 700284 543464 700312
rect 57756 700272 57762 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 147214 683136 147220 683188
rect 147272 683176 147278 683188
rect 580166 683176 580172 683188
rect 147272 683148 580172 683176
rect 147272 683136 147278 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 104894 647844 104900 647896
rect 104952 647884 104958 647896
rect 434898 647884 434904 647896
rect 104952 647856 434904 647884
rect 104952 647844 104958 647856
rect 434898 647844 434904 647856
rect 434956 647844 434962 647896
rect 299474 646484 299480 646536
rect 299532 646524 299538 646536
rect 405918 646524 405924 646536
rect 299532 646496 405924 646524
rect 299532 646484 299538 646496
rect 405918 646484 405924 646496
rect 405976 646484 405982 646536
rect 364334 645124 364340 645176
rect 364392 645164 364398 645176
rect 428366 645164 428372 645176
rect 364392 645136 428372 645164
rect 364392 645124 364398 645136
rect 428366 645124 428372 645136
rect 428424 645124 428430 645176
rect 322566 643084 322572 643136
rect 322624 643124 322630 643136
rect 436094 643124 436100 643136
rect 322624 643096 436100 643124
rect 322624 643084 322630 643096
rect 436094 643084 436100 643096
rect 436152 643084 436158 643136
rect 322474 642676 322480 642728
rect 322532 642716 322538 642728
rect 346578 642716 346584 642728
rect 322532 642688 346584 642716
rect 322532 642676 322538 642688
rect 346578 642676 346584 642688
rect 346636 642676 346642 642728
rect 323670 642608 323676 642660
rect 323728 642648 323734 642660
rect 401686 642648 401692 642660
rect 323728 642620 401692 642648
rect 323728 642608 323734 642620
rect 401686 642608 401692 642620
rect 401744 642608 401750 642660
rect 316770 642540 316776 642592
rect 316828 642580 316834 642592
rect 342254 642580 342260 642592
rect 316828 642552 342260 642580
rect 316828 642540 316834 642552
rect 342254 642540 342260 642552
rect 342312 642540 342318 642592
rect 309778 642472 309784 642524
rect 309836 642512 309842 642524
rect 373994 642512 374000 642524
rect 309836 642484 374000 642512
rect 309836 642472 309842 642484
rect 373994 642472 374000 642484
rect 374052 642472 374058 642524
rect 323762 642404 323768 642456
rect 323820 642444 323826 642456
rect 369118 642444 369124 642456
rect 323820 642416 369124 642444
rect 323820 642404 323826 642416
rect 369118 642404 369124 642416
rect 369176 642404 369182 642456
rect 318150 642336 318156 642388
rect 318208 642376 318214 642388
rect 364610 642376 364616 642388
rect 318208 642348 364616 642376
rect 318208 642336 318214 642348
rect 364610 642336 364616 642348
rect 364668 642336 364674 642388
rect 324866 642268 324872 642320
rect 324924 642308 324930 642320
rect 378134 642308 378140 642320
rect 324924 642280 378140 642308
rect 324924 642268 324930 642280
rect 378134 642268 378140 642280
rect 378192 642268 378198 642320
rect 322290 642200 322296 642252
rect 322348 642240 322354 642252
rect 355594 642240 355600 642252
rect 322348 642212 355600 642240
rect 322348 642200 322354 642212
rect 355594 642200 355600 642212
rect 355652 642200 355658 642252
rect 355686 642200 355692 642252
rect 355744 642240 355750 642252
rect 414842 642240 414848 642252
rect 355744 642212 414848 642240
rect 355744 642200 355750 642212
rect 414842 642200 414848 642212
rect 414900 642200 414906 642252
rect 307018 642132 307024 642184
rect 307076 642172 307082 642184
rect 337562 642172 337568 642184
rect 307076 642144 337568 642172
rect 307076 642132 307082 642144
rect 337562 642132 337568 642144
rect 337620 642132 337626 642184
rect 347590 642132 347596 642184
rect 347648 642172 347654 642184
rect 410334 642172 410340 642184
rect 347648 642144 410340 642172
rect 347648 642132 347654 642144
rect 410334 642132 410340 642144
rect 410392 642132 410398 642184
rect 323946 642064 323952 642116
rect 324004 642104 324010 642116
rect 387794 642104 387800 642116
rect 324004 642076 387800 642104
rect 324004 642064 324010 642076
rect 387794 642064 387800 642076
rect 387852 642064 387858 642116
rect 320910 641996 320916 642048
rect 320968 642036 320974 642048
rect 392302 642036 392308 642048
rect 320968 642008 392308 642036
rect 320968 641996 320974 642008
rect 392302 641996 392308 642008
rect 392360 641996 392366 642048
rect 311158 641928 311164 641980
rect 311216 641968 311222 641980
rect 383654 641968 383660 641980
rect 311216 641940 383660 641968
rect 311216 641928 311222 641940
rect 383654 641928 383660 641940
rect 383712 641928 383718 641980
rect 337102 641860 337108 641912
rect 337160 641900 337166 641912
rect 351086 641900 351092 641912
rect 337160 641872 351092 641900
rect 337160 641860 337166 641872
rect 351086 641860 351092 641872
rect 351144 641860 351150 641912
rect 322382 641792 322388 641844
rect 322440 641832 322446 641844
rect 432874 641832 432880 641844
rect 322440 641804 432880 641832
rect 322440 641792 322446 641804
rect 432874 641792 432880 641804
rect 432932 641792 432938 641844
rect 323854 641724 323860 641776
rect 323912 641764 323918 641776
rect 328546 641764 328552 641776
rect 323912 641736 328552 641764
rect 323912 641724 323918 641736
rect 328546 641724 328552 641736
rect 328604 641724 328610 641776
rect 365622 641724 365628 641776
rect 365680 641764 365686 641776
rect 419534 641764 419540 641776
rect 365680 641736 419540 641764
rect 365680 641724 365686 641736
rect 419534 641724 419540 641736
rect 419592 641764 419598 641776
rect 457438 641764 457444 641776
rect 419592 641736 457444 641764
rect 419592 641724 419598 641736
rect 457438 641724 457444 641736
rect 457496 641724 457502 641776
rect 319438 641180 319444 641232
rect 319496 641220 319502 641232
rect 436186 641220 436192 641232
rect 319496 641192 436192 641220
rect 319496 641180 319502 641192
rect 436186 641180 436192 641192
rect 436244 641180 436250 641232
rect 233234 641112 233240 641164
rect 233292 641152 233298 641164
rect 360194 641152 360200 641164
rect 233292 641124 360200 641152
rect 233292 641112 233298 641124
rect 360194 641112 360200 641124
rect 360252 641112 360258 641164
rect 147582 641044 147588 641096
rect 147640 641084 147646 641096
rect 164510 641084 164516 641096
rect 147640 641056 164516 641084
rect 147640 641044 147646 641056
rect 164510 641044 164516 641056
rect 164568 641044 164574 641096
rect 324222 641044 324228 641096
rect 324280 641084 324286 641096
rect 494054 641084 494060 641096
rect 324280 641056 494060 641084
rect 324280 641044 324286 641056
rect 494054 641044 494060 641056
rect 494112 641044 494118 641096
rect 131114 640976 131120 641028
rect 131172 641016 131178 641028
rect 161566 641016 161572 641028
rect 131172 640988 161572 641016
rect 131172 640976 131178 640988
rect 161566 640976 161572 640988
rect 161624 640976 161630 641028
rect 238018 640976 238024 641028
rect 238076 641016 238082 641028
rect 365622 641016 365628 641028
rect 238076 640988 365628 641016
rect 238076 640976 238082 640988
rect 365622 640976 365628 640988
rect 365680 640976 365686 641028
rect 145006 640908 145012 640960
rect 145064 640948 145070 640960
rect 207658 640948 207664 640960
rect 145064 640920 207664 640948
rect 145064 640908 145070 640920
rect 207658 640908 207664 640920
rect 207716 640908 207722 640960
rect 239490 640908 239496 640960
rect 239548 640948 239554 640960
rect 257430 640948 257436 640960
rect 239548 640920 257436 640948
rect 239548 640908 239554 640920
rect 257430 640908 257436 640920
rect 257488 640908 257494 640960
rect 323578 640908 323584 640960
rect 323636 640948 323642 640960
rect 457622 640948 457628 640960
rect 323636 640920 457628 640948
rect 323636 640908 323642 640920
rect 457622 640908 457628 640920
rect 457680 640908 457686 640960
rect 115382 640840 115388 640892
rect 115440 640880 115446 640892
rect 124674 640880 124680 640892
rect 115440 640852 124680 640880
rect 115440 640840 115446 640852
rect 124674 640840 124680 640852
rect 124732 640840 124738 640892
rect 148870 640840 148876 640892
rect 148928 640880 148934 640892
rect 172882 640880 172888 640892
rect 148928 640852 172888 640880
rect 148928 640840 148934 640852
rect 172882 640840 172888 640852
rect 172940 640840 172946 640892
rect 235258 640840 235264 640892
rect 235316 640880 235322 640892
rect 292206 640880 292212 640892
rect 235316 640852 292212 640880
rect 235316 640840 235322 640852
rect 292206 640840 292212 640852
rect 292264 640840 292270 640892
rect 322658 640840 322664 640892
rect 322716 640880 322722 640892
rect 457714 640880 457720 640892
rect 322716 640852 457720 640880
rect 322716 640840 322722 640852
rect 457714 640840 457720 640852
rect 457772 640840 457778 640892
rect 124398 640812 124404 640824
rect 103486 640784 124404 640812
rect 69014 640704 69020 640756
rect 69072 640744 69078 640756
rect 103486 640744 103514 640784
rect 124398 640772 124404 640784
rect 124456 640772 124462 640824
rect 140774 640772 140780 640824
rect 140832 640812 140838 640824
rect 167086 640812 167092 640824
rect 140832 640784 167092 640812
rect 140832 640772 140838 640784
rect 167086 640772 167092 640784
rect 167144 640772 167150 640824
rect 226334 640772 226340 640824
rect 226392 640812 226398 640824
rect 300578 640812 300584 640824
rect 226392 640784 300584 640812
rect 226392 640772 226398 640784
rect 300578 640772 300584 640784
rect 300636 640772 300642 640824
rect 314102 640772 314108 640824
rect 314160 640812 314166 640824
rect 457806 640812 457812 640824
rect 314160 640784 457812 640812
rect 314160 640772 314166 640784
rect 457806 640772 457812 640784
rect 457864 640772 457870 640824
rect 69072 640716 103514 640744
rect 69072 640704 69078 640716
rect 117958 640704 117964 640756
rect 118016 640744 118022 640756
rect 124490 640744 124496 640756
rect 118016 640716 124496 640744
rect 118016 640704 118022 640716
rect 124490 640704 124496 640716
rect 124548 640704 124554 640756
rect 148778 640704 148784 640756
rect 148836 640744 148842 640756
rect 176102 640744 176108 640756
rect 148836 640716 176108 640744
rect 148836 640704 148842 640716
rect 176102 640704 176108 640716
rect 176160 640704 176166 640756
rect 239582 640704 239588 640756
rect 239640 640744 239646 640756
rect 274818 640744 274824 640756
rect 239640 640716 274824 640744
rect 239640 640704 239646 640716
rect 274818 640704 274824 640716
rect 274876 640704 274882 640756
rect 316678 640704 316684 640756
rect 316736 640744 316742 640756
rect 471606 640744 471612 640756
rect 316736 640716 471612 640744
rect 316736 640704 316742 640716
rect 471606 640704 471612 640716
rect 471664 640704 471670 640756
rect 112162 640636 112168 640688
rect 112220 640676 112226 640688
rect 122834 640676 122840 640688
rect 112220 640648 122840 640676
rect 112220 640636 112226 640648
rect 122834 640636 122840 640648
rect 122892 640636 122898 640688
rect 149514 640636 149520 640688
rect 149572 640676 149578 640688
rect 190546 640676 190552 640688
rect 149572 640648 190552 640676
rect 149572 640636 149578 640648
rect 190546 640636 190552 640648
rect 190604 640636 190610 640688
rect 236638 640636 236644 640688
rect 236696 640676 236702 640688
rect 396810 640676 396816 640688
rect 236696 640648 396816 640676
rect 236696 640636 236702 640648
rect 396810 640636 396816 640648
rect 396868 640636 396874 640688
rect 60734 640568 60740 640620
rect 60792 640608 60798 640620
rect 97994 640608 98000 640620
rect 60792 640580 98000 640608
rect 60792 640568 60798 640580
rect 97994 640568 98000 640580
rect 98052 640568 98058 640620
rect 106366 640568 106372 640620
rect 106424 640608 106430 640620
rect 121454 640608 121460 640620
rect 106424 640580 121460 640608
rect 106424 640568 106430 640580
rect 121454 640568 121460 640580
rect 121512 640568 121518 640620
rect 142154 640568 142160 640620
rect 142212 640608 142218 640620
rect 184474 640608 184480 640620
rect 142212 640580 184480 640608
rect 142212 640568 142218 640580
rect 184474 640568 184480 640580
rect 184532 640568 184538 640620
rect 217410 640568 217416 640620
rect 217468 640608 217474 640620
rect 254854 640608 254860 640620
rect 217468 640580 254860 640608
rect 217468 640568 217474 640580
rect 254854 640568 254860 640580
rect 254912 640568 254918 640620
rect 314010 640568 314016 640620
rect 314068 640608 314074 640620
rect 483198 640608 483204 640620
rect 314068 640580 483204 640608
rect 314068 640568 314074 640580
rect 483198 640568 483204 640580
rect 483256 640568 483262 640620
rect 54846 640500 54852 640552
rect 54904 640540 54910 640552
rect 88978 640540 88984 640552
rect 54904 640512 88984 640540
rect 54904 640500 54910 640512
rect 88978 640500 88984 640512
rect 89036 640500 89042 640552
rect 103790 640500 103796 640552
rect 103848 640540 103854 640552
rect 121546 640540 121552 640552
rect 103848 640512 121552 640540
rect 103848 640500 103854 640512
rect 121546 640500 121552 640512
rect 121604 640500 121610 640552
rect 144914 640500 144920 640552
rect 144972 640540 144978 640552
rect 196066 640540 196072 640552
rect 144972 640512 196072 640540
rect 144972 640500 144978 640512
rect 196066 640500 196072 640512
rect 196124 640500 196130 640552
rect 231118 640500 231124 640552
rect 231176 640540 231182 640552
rect 243538 640540 243544 640552
rect 231176 640512 243544 640540
rect 231176 640500 231182 640512
rect 243538 640500 243544 640512
rect 243596 640500 243602 640552
rect 249702 640500 249708 640552
rect 249760 640540 249766 640552
rect 295426 640540 295432 640552
rect 249760 640512 295432 640540
rect 249760 640500 249766 640512
rect 295426 640500 295432 640512
rect 295484 640500 295490 640552
rect 319530 640500 319536 640552
rect 319588 640540 319594 640552
rect 494790 640540 494796 640552
rect 319588 640512 494796 640540
rect 319588 640500 319594 640512
rect 494790 640500 494796 640512
rect 494848 640500 494854 640552
rect 55122 640432 55128 640484
rect 55180 640472 55186 640484
rect 92198 640472 92204 640484
rect 55180 640444 92204 640472
rect 55180 640432 55186 640444
rect 92198 640432 92204 640444
rect 92256 640432 92262 640484
rect 94774 640432 94780 640484
rect 94832 640472 94838 640484
rect 120902 640472 120908 640484
rect 94832 640444 120908 640472
rect 94832 640432 94838 640444
rect 120902 640432 120908 640444
rect 120960 640432 120966 640484
rect 147306 640432 147312 640484
rect 147364 640472 147370 640484
rect 199286 640472 199292 640484
rect 147364 640444 199292 640472
rect 147364 640432 147370 640444
rect 199286 640432 199292 640444
rect 199344 640432 199350 640484
rect 237374 640432 237380 640484
rect 237432 640472 237438 640484
rect 289630 640472 289636 640484
rect 237432 640444 289636 640472
rect 237432 640432 237438 640444
rect 289630 640432 289636 640444
rect 289688 640432 289694 640484
rect 322198 640432 322204 640484
rect 322256 640472 322262 640484
rect 501230 640472 501236 640484
rect 322256 640444 501236 640472
rect 322256 640432 322262 640444
rect 501230 640432 501236 640444
rect 501288 640432 501294 640484
rect 55030 640364 55036 640416
rect 55088 640404 55094 640416
rect 65794 640404 65800 640416
rect 55088 640376 65800 640404
rect 55088 640364 55094 640376
rect 65794 640364 65800 640376
rect 65852 640364 65858 640416
rect 100570 640364 100576 640416
rect 100628 640404 100634 640416
rect 117958 640404 117964 640416
rect 100628 640376 117964 640404
rect 100628 640364 100634 640376
rect 117958 640364 117964 640376
rect 118016 640364 118022 640416
rect 120994 640404 121000 640416
rect 118068 640376 121000 640404
rect 56502 640296 56508 640348
rect 56560 640336 56566 640348
rect 77386 640336 77392 640348
rect 56560 640308 77392 640336
rect 56560 640296 56566 640308
rect 77386 640296 77392 640308
rect 77444 640296 77450 640348
rect 109586 640296 109592 640348
rect 109644 640336 109650 640348
rect 118068 640336 118096 640376
rect 120994 640364 121000 640376
rect 121052 640364 121058 640416
rect 149606 640364 149612 640416
rect 149664 640404 149670 640416
rect 201862 640404 201868 640416
rect 149664 640376 201868 640404
rect 149664 640364 149670 640376
rect 201862 640364 201868 640376
rect 201920 640364 201926 640416
rect 205542 640364 205548 640416
rect 205600 640404 205606 640416
rect 212626 640404 212632 640416
rect 205600 640376 212632 640404
rect 205600 640364 205606 640376
rect 212626 640364 212632 640376
rect 212684 640364 212690 640416
rect 238110 640364 238116 640416
rect 238168 640404 238174 640416
rect 251634 640404 251640 640416
rect 238168 640376 251640 640404
rect 238168 640364 238174 640376
rect 251634 640364 251640 640376
rect 251692 640364 251698 640416
rect 319622 640364 319628 640416
rect 319680 640404 319686 640416
rect 511994 640404 512000 640416
rect 319680 640376 512000 640404
rect 319680 640364 319686 640376
rect 511994 640364 512000 640376
rect 512052 640364 512058 640416
rect 109644 640308 118096 640336
rect 109644 640296 109650 640308
rect 118234 640296 118240 640348
rect 118292 640336 118298 640348
rect 124582 640336 124588 640348
rect 118292 640308 124588 640336
rect 118292 640296 118298 640308
rect 124582 640296 124588 640308
rect 124640 640296 124646 640348
rect 133874 640296 133880 640348
rect 133932 640336 133938 640348
rect 149974 640336 149980 640348
rect 133932 640308 149980 640336
rect 133932 640296 133938 640308
rect 149974 640296 149980 640308
rect 150032 640296 150038 640348
rect 243538 640296 243544 640348
rect 243596 640336 243602 640348
rect 249058 640336 249064 640348
rect 243596 640308 249064 640336
rect 243596 640296 243602 640308
rect 249058 640296 249064 640308
rect 249116 640296 249122 640348
rect 255314 640296 255320 640348
rect 255372 640336 255378 640348
rect 263226 640336 263232 640348
rect 255372 640308 263232 640336
rect 255372 640296 255378 640308
rect 263226 640296 263232 640308
rect 263284 640296 263290 640348
rect 316862 640296 316868 640348
rect 316920 640336 316926 640348
rect 512178 640336 512184 640348
rect 316920 640308 512184 640336
rect 316920 640296 316926 640308
rect 512178 640296 512184 640308
rect 512236 640296 512242 640348
rect 223574 639820 223580 639872
rect 223632 639860 223638 639872
rect 249702 639860 249708 639872
rect 223632 639832 249708 639860
rect 223632 639820 223638 639832
rect 249702 639820 249708 639832
rect 249760 639820 249766 639872
rect 222194 639752 222200 639804
rect 222252 639792 222258 639804
rect 255314 639792 255320 639804
rect 222252 639764 255320 639792
rect 222252 639752 222258 639764
rect 255314 639752 255320 639764
rect 255372 639752 255378 639804
rect 3418 639684 3424 639736
rect 3476 639724 3482 639736
rect 337102 639724 337108 639736
rect 3476 639696 337108 639724
rect 3476 639684 3482 639696
rect 337102 639684 337108 639696
rect 337160 639684 337166 639736
rect 3602 639616 3608 639668
rect 3660 639656 3666 639668
rect 347590 639656 347596 639668
rect 3660 639628 347596 639656
rect 3660 639616 3666 639628
rect 347590 639616 347596 639628
rect 347648 639616 347654 639668
rect 3694 639548 3700 639600
rect 3752 639588 3758 639600
rect 355502 639588 355508 639600
rect 3752 639560 355508 639588
rect 3752 639548 3758 639560
rect 355502 639548 355508 639560
rect 355560 639548 355566 639600
rect 238938 639208 238944 639260
rect 238996 639248 239002 639260
rect 580350 639248 580356 639260
rect 238996 639220 580356 639248
rect 238996 639208 239002 639220
rect 580350 639208 580356 639220
rect 580408 639208 580414 639260
rect 231210 639140 231216 639192
rect 231268 639180 231274 639192
rect 272242 639180 272248 639192
rect 231268 639152 272248 639180
rect 231268 639140 231274 639152
rect 272242 639140 272248 639152
rect 272300 639140 272306 639192
rect 316954 639140 316960 639192
rect 317012 639180 317018 639192
rect 457530 639180 457536 639192
rect 317012 639152 457536 639180
rect 317012 639140 317018 639152
rect 457530 639140 457536 639152
rect 457588 639140 457594 639192
rect 239030 639072 239036 639124
rect 239088 639112 239094 639124
rect 433334 639112 433340 639124
rect 239088 639084 433340 639112
rect 239088 639072 239094 639084
rect 433334 639072 433340 639084
rect 433392 639072 433398 639124
rect 149882 639004 149888 639056
rect 149940 639044 149946 639056
rect 170306 639044 170312 639056
rect 149940 639016 170312 639044
rect 149940 639004 149946 639016
rect 170306 639004 170312 639016
rect 170364 639004 170370 639056
rect 215938 639004 215944 639056
rect 215996 639044 216002 639056
rect 269022 639044 269028 639056
rect 215996 639016 269028 639044
rect 215996 639004 216002 639016
rect 269022 639004 269028 639016
rect 269080 639004 269086 639056
rect 317046 639004 317052 639056
rect 317104 639044 317110 639056
rect 512086 639044 512092 639056
rect 317104 639016 512092 639044
rect 317104 639004 317110 639016
rect 512086 639004 512092 639016
rect 512144 639004 512150 639056
rect 148318 638936 148324 638988
rect 148376 638976 148382 638988
rect 153194 638976 153200 638988
rect 148376 638948 153200 638976
rect 148376 638936 148382 638948
rect 153194 638936 153200 638948
rect 153252 638936 153258 638988
rect 3510 638188 3516 638240
rect 3568 638228 3574 638240
rect 321002 638228 321008 638240
rect 3568 638200 321008 638228
rect 3568 638188 3574 638200
rect 321002 638188 321008 638200
rect 321060 638188 321066 638240
rect 236730 638052 236736 638104
rect 236788 638092 236794 638104
rect 245654 638092 245660 638104
rect 236788 638064 245660 638092
rect 236788 638052 236794 638064
rect 245654 638052 245660 638064
rect 245712 638052 245718 638104
rect 126238 637984 126244 638036
rect 126296 638024 126302 638036
rect 187694 638024 187700 638036
rect 126296 637996 187700 638024
rect 126296 637984 126302 637996
rect 187694 637984 187700 637996
rect 187752 637984 187758 638036
rect 228358 637984 228364 638036
rect 228416 638024 228422 638036
rect 266262 638024 266268 638036
rect 228416 637996 266268 638024
rect 228416 637984 228422 637996
rect 266262 637984 266268 637996
rect 266320 637984 266326 638036
rect 59354 637916 59360 637968
rect 59412 637956 59418 637968
rect 60734 637956 60740 637968
rect 59412 637928 60740 637956
rect 59412 637916 59418 637928
rect 60734 637916 60740 637928
rect 60792 637916 60798 637968
rect 148962 637916 148968 637968
rect 149020 637956 149026 637968
rect 158714 637956 158720 637968
rect 149020 637928 158720 637956
rect 149020 637916 149026 637928
rect 158714 637916 158720 637928
rect 158772 637916 158778 637968
rect 216030 637916 216036 637968
rect 216088 637956 216094 637968
rect 260374 637956 260380 637968
rect 216088 637928 260380 637956
rect 216088 637916 216094 637928
rect 260374 637916 260380 637928
rect 260432 637916 260438 637968
rect 54938 637848 54944 637900
rect 54996 637888 55002 637900
rect 62942 637888 62948 637900
rect 54996 637860 62948 637888
rect 54996 637848 55002 637860
rect 62942 637848 62948 637860
rect 63000 637848 63006 637900
rect 136634 637848 136640 637900
rect 136692 637888 136698 637900
rect 178678 637888 178684 637900
rect 136692 637860 178684 637888
rect 136692 637848 136698 637860
rect 178678 637848 178684 637860
rect 178736 637848 178742 637900
rect 226978 637848 226984 637900
rect 227036 637888 227042 637900
rect 283558 637888 283564 637900
rect 227036 637860 283564 637888
rect 227036 637848 227042 637860
rect 283558 637848 283564 637860
rect 283616 637848 283622 637900
rect 56410 637780 56416 637832
rect 56468 637820 56474 637832
rect 71222 637820 71228 637832
rect 56468 637792 71228 637820
rect 56468 637780 56474 637792
rect 71222 637780 71228 637792
rect 71280 637780 71286 637832
rect 86770 637780 86776 637832
rect 86828 637820 86834 637832
rect 125778 637820 125784 637832
rect 86828 637792 125784 637820
rect 86828 637780 86834 637792
rect 125778 637780 125784 637792
rect 125836 637780 125842 637832
rect 140038 637780 140044 637832
rect 140096 637820 140102 637832
rect 193490 637820 193496 637832
rect 140096 637792 193496 637820
rect 140096 637780 140102 637792
rect 193490 637780 193496 637792
rect 193548 637780 193554 637832
rect 220078 637780 220084 637832
rect 220136 637820 220142 637832
rect 280246 637820 280252 637832
rect 220136 637792 280252 637820
rect 220136 637780 220142 637792
rect 280246 637780 280252 637792
rect 280304 637780 280310 637832
rect 56318 637712 56324 637764
rect 56376 637752 56382 637764
rect 74626 637752 74632 637764
rect 56376 637724 74632 637752
rect 56376 637712 56382 637724
rect 74626 637712 74632 637724
rect 74684 637712 74690 637764
rect 124214 637712 124220 637764
rect 124272 637752 124278 637764
rect 182082 637752 182088 637764
rect 124272 637724 182088 637752
rect 124272 637712 124278 637724
rect 182082 637712 182088 637724
rect 182140 637712 182146 637764
rect 214558 637712 214564 637764
rect 214616 637752 214622 637764
rect 286134 637752 286140 637764
rect 214616 637724 286140 637752
rect 214616 637712 214622 637724
rect 286134 637712 286140 637724
rect 286192 637712 286198 637764
rect 57790 637644 57796 637696
rect 57848 637684 57854 637696
rect 80238 637684 80244 637696
rect 57848 637656 80244 637684
rect 57848 637644 57854 637656
rect 80238 637644 80244 637656
rect 80296 637644 80302 637696
rect 83458 637644 83464 637696
rect 83516 637684 83522 637696
rect 124306 637684 124312 637696
rect 83516 637656 124312 637684
rect 83516 637644 83522 637656
rect 124306 637644 124312 637656
rect 124364 637644 124370 637696
rect 146110 637644 146116 637696
rect 146168 637684 146174 637696
rect 155494 637684 155500 637696
rect 146168 637656 155500 637684
rect 146168 637644 146174 637656
rect 155494 637644 155500 637656
rect 155552 637644 155558 637696
rect 217318 637644 217324 637696
rect 217376 637684 217382 637696
rect 297726 637684 297732 637696
rect 217376 637656 297732 637684
rect 217376 637644 217382 637656
rect 297726 637644 297732 637656
rect 297784 637644 297790 637696
rect 57882 637576 57888 637628
rect 57940 637616 57946 637628
rect 146202 637616 146208 637628
rect 57940 637588 146208 637616
rect 57940 637576 57946 637588
rect 146202 637576 146208 637588
rect 146260 637616 146266 637628
rect 238018 637616 238024 637628
rect 146260 637588 238024 637616
rect 146260 637576 146266 637588
rect 238018 637576 238024 637588
rect 238076 637576 238082 637628
rect 238202 637576 238208 637628
rect 238260 637616 238266 637628
rect 277670 637616 277676 637628
rect 238260 637588 277676 637616
rect 238260 637576 238266 637588
rect 277670 637576 277676 637588
rect 277728 637576 277734 637628
rect 239398 637508 239404 637560
rect 239456 637548 239462 637560
rect 242894 637548 242900 637560
rect 239456 637520 242900 637548
rect 239456 637508 239462 637520
rect 242894 637508 242900 637520
rect 242952 637508 242958 637560
rect 213914 636828 213920 636880
rect 213972 636868 213978 636880
rect 237374 636868 237380 636880
rect 213972 636840 237380 636868
rect 213972 636828 213978 636840
rect 237374 636828 237380 636840
rect 237432 636828 237438 636880
rect 144178 635196 144184 635248
rect 144236 635236 144242 635248
rect 147122 635236 147128 635248
rect 144236 635208 147128 635236
rect 144236 635196 144242 635208
rect 147122 635196 147128 635208
rect 147180 635196 147186 635248
rect 232498 635128 232504 635180
rect 232556 635168 232562 635180
rect 237374 635168 237380 635180
rect 232556 635140 237380 635168
rect 232556 635128 232562 635140
rect 237374 635128 237380 635140
rect 237432 635128 237438 635180
rect 465442 634856 465448 634908
rect 465500 634896 465506 634908
rect 465500 634868 470594 634896
rect 465500 634856 465506 634868
rect 470566 634828 470594 634868
rect 580258 634828 580264 634840
rect 470566 634800 580264 634828
rect 580258 634788 580264 634800
rect 580316 634788 580322 634840
rect 312538 633428 312544 633480
rect 312596 633468 312602 633480
rect 321554 633468 321560 633480
rect 312596 633440 321560 633468
rect 312596 633428 312602 633440
rect 321554 633428 321560 633440
rect 321612 633428 321618 633480
rect 238846 629960 238852 630012
rect 238904 630000 238910 630012
rect 239766 630000 239772 630012
rect 238904 629972 239772 630000
rect 238904 629960 238910 629972
rect 239766 629960 239772 629972
rect 239824 629960 239830 630012
rect 233326 629280 233332 629332
rect 233384 629320 233390 629332
rect 237374 629320 237380 629332
rect 233384 629292 237380 629320
rect 233384 629280 233390 629292
rect 237374 629280 237380 629292
rect 237432 629280 237438 629332
rect 313918 629280 313924 629332
rect 313976 629320 313982 629332
rect 321554 629320 321560 629332
rect 313976 629292 321560 629320
rect 313976 629280 313982 629292
rect 321554 629280 321560 629292
rect 321612 629280 321618 629332
rect 140866 626560 140872 626612
rect 140924 626600 140930 626612
rect 146294 626600 146300 626612
rect 140924 626572 146300 626600
rect 140924 626560 140930 626572
rect 146294 626560 146300 626572
rect 146352 626560 146358 626612
rect 216122 626560 216128 626612
rect 216180 626600 216186 626612
rect 237374 626600 237380 626612
rect 216180 626572 237380 626600
rect 216180 626560 216186 626572
rect 237374 626560 237380 626572
rect 237432 626560 237438 626612
rect 318058 623772 318064 623824
rect 318116 623812 318122 623824
rect 321554 623812 321560 623824
rect 318116 623784 321560 623812
rect 318116 623772 318122 623784
rect 321554 623772 321560 623784
rect 321612 623772 321618 623824
rect 132494 622412 132500 622464
rect 132552 622452 132558 622464
rect 146294 622452 146300 622464
rect 132552 622424 146300 622452
rect 132552 622412 132558 622424
rect 146294 622412 146300 622424
rect 146352 622412 146358 622464
rect 222838 622412 222844 622464
rect 222896 622452 222902 622464
rect 237374 622452 237380 622464
rect 222896 622424 237380 622452
rect 222896 622412 222902 622424
rect 237374 622412 237380 622424
rect 237432 622412 237438 622464
rect 223666 619624 223672 619676
rect 223724 619664 223730 619676
rect 237374 619664 237380 619676
rect 223724 619636 237380 619664
rect 223724 619624 223730 619636
rect 237374 619624 237380 619636
rect 237432 619624 237438 619676
rect 311250 619624 311256 619676
rect 311308 619664 311314 619676
rect 321554 619664 321560 619676
rect 311308 619636 321560 619664
rect 311308 619624 311314 619636
rect 321554 619624 321560 619636
rect 321612 619624 321618 619676
rect 218054 616836 218060 616888
rect 218112 616876 218118 616888
rect 237374 616876 237380 616888
rect 218112 616848 237380 616876
rect 218112 616836 218118 616848
rect 237374 616836 237380 616848
rect 237432 616836 237438 616888
rect 309870 614116 309876 614168
rect 309928 614156 309934 614168
rect 321554 614156 321560 614168
rect 309928 614128 321560 614156
rect 309928 614116 309934 614128
rect 321554 614116 321560 614128
rect 321612 614116 321618 614168
rect 314194 609968 314200 610020
rect 314252 610008 314258 610020
rect 321554 610008 321560 610020
rect 314252 609980 321560 610008
rect 314252 609968 314258 609980
rect 321554 609968 321560 609980
rect 321612 609968 321618 610020
rect 220170 607180 220176 607232
rect 220228 607220 220234 607232
rect 237374 607220 237380 607232
rect 220228 607192 237380 607220
rect 220228 607180 220234 607192
rect 237374 607180 237380 607192
rect 237432 607180 237438 607232
rect 311342 605820 311348 605872
rect 311400 605860 311406 605872
rect 321554 605860 321560 605872
rect 311400 605832 321560 605860
rect 311400 605820 311406 605832
rect 321554 605820 321560 605832
rect 321612 605820 321618 605872
rect 128998 604460 129004 604512
rect 129056 604500 129062 604512
rect 146294 604500 146300 604512
rect 129056 604472 146300 604500
rect 129056 604460 129062 604472
rect 146294 604460 146300 604472
rect 146352 604460 146358 604512
rect 235442 604460 235448 604512
rect 235500 604500 235506 604512
rect 237374 604500 237380 604512
rect 235500 604472 237380 604500
rect 235500 604460 235506 604472
rect 237374 604460 237380 604472
rect 237432 604460 237438 604512
rect 303154 603712 303160 603764
rect 303212 603752 303218 603764
rect 322658 603752 322664 603764
rect 303212 603724 322664 603752
rect 303212 603712 303218 603724
rect 322658 603712 322664 603724
rect 322716 603712 322722 603764
rect 124122 603100 124128 603152
rect 124180 603140 124186 603152
rect 145558 603140 145564 603152
rect 124180 603112 145564 603140
rect 124180 603100 124186 603112
rect 145558 603100 145564 603112
rect 145616 603100 145622 603152
rect 214650 601672 214656 601724
rect 214708 601712 214714 601724
rect 237374 601712 237380 601724
rect 214708 601684 237380 601712
rect 214708 601672 214714 601684
rect 237374 601672 237380 601684
rect 237432 601672 237438 601724
rect 123294 600992 123300 601044
rect 123352 601032 123358 601044
rect 123478 601032 123484 601044
rect 123352 601004 123484 601032
rect 123352 600992 123358 601004
rect 123478 600992 123484 601004
rect 123536 600992 123542 601044
rect 229738 597524 229744 597576
rect 229796 597564 229802 597576
rect 237374 597564 237380 597576
rect 229796 597536 237380 597564
rect 229796 597524 229802 597536
rect 237374 597524 237380 597536
rect 237432 597524 237438 597576
rect 304258 596164 304264 596216
rect 304316 596204 304322 596216
rect 321554 596204 321560 596216
rect 304316 596176 321560 596204
rect 304316 596164 304322 596176
rect 321554 596164 321560 596176
rect 321612 596164 321618 596216
rect 231854 594804 231860 594856
rect 231912 594844 231918 594856
rect 237374 594844 237380 594856
rect 231912 594816 237380 594844
rect 231912 594804 231918 594816
rect 237374 594804 237380 594816
rect 237432 594804 237438 594856
rect 125594 592016 125600 592068
rect 125652 592056 125658 592068
rect 146294 592056 146300 592068
rect 125652 592028 146300 592056
rect 125652 592016 125658 592028
rect 146294 592016 146300 592028
rect 146352 592016 146358 592068
rect 235350 592016 235356 592068
rect 235408 592056 235414 592068
rect 237374 592056 237380 592068
rect 235408 592028 237380 592056
rect 235408 592016 235414 592028
rect 237374 592016 237380 592028
rect 237432 592016 237438 592068
rect 307110 590656 307116 590708
rect 307168 590696 307174 590708
rect 321554 590696 321560 590708
rect 307168 590668 321560 590696
rect 307168 590656 307174 590668
rect 321554 590656 321560 590668
rect 321612 590656 321618 590708
rect 130378 589296 130384 589348
rect 130436 589336 130442 589348
rect 146294 589336 146300 589348
rect 130436 589308 146300 589336
rect 130436 589296 130442 589308
rect 146294 589296 146300 589308
rect 146352 589296 146358 589348
rect 233878 589296 233884 589348
rect 233936 589336 233942 589348
rect 237374 589336 237380 589348
rect 233936 589308 237380 589336
rect 233936 589296 233942 589308
rect 237374 589296 237380 589308
rect 237432 589296 237438 589348
rect 57698 589228 57704 589280
rect 57756 589268 57762 589280
rect 58618 589268 58624 589280
rect 57756 589240 58624 589268
rect 57756 589228 57762 589240
rect 58618 589228 58624 589240
rect 58676 589228 58682 589280
rect 139394 586508 139400 586560
rect 139452 586548 139458 586560
rect 146294 586548 146300 586560
rect 139452 586520 146300 586548
rect 139452 586508 139458 586520
rect 146294 586508 146300 586520
rect 146352 586508 146358 586560
rect 214742 586508 214748 586560
rect 214800 586548 214806 586560
rect 237374 586548 237380 586560
rect 214800 586520 237380 586548
rect 214800 586508 214806 586520
rect 237374 586508 237380 586520
rect 237432 586508 237438 586560
rect 309962 586508 309968 586560
rect 310020 586548 310026 586560
rect 321554 586548 321560 586560
rect 310020 586520 321560 586548
rect 310020 586508 310026 586520
rect 321554 586508 321560 586520
rect 321612 586508 321618 586560
rect 513282 586508 513288 586560
rect 513340 586548 513346 586560
rect 560938 586548 560944 586560
rect 513340 586520 560944 586548
rect 513340 586508 513346 586520
rect 560938 586508 560944 586520
rect 560996 586508 561002 586560
rect 226426 583720 226432 583772
rect 226484 583760 226490 583772
rect 237374 583760 237380 583772
rect 226484 583732 237380 583760
rect 226484 583720 226490 583732
rect 237374 583720 237380 583732
rect 237432 583720 237438 583772
rect 120718 581612 120724 581664
rect 120776 581652 120782 581664
rect 121178 581652 121184 581664
rect 120776 581624 121184 581652
rect 120776 581612 120782 581624
rect 121178 581612 121184 581624
rect 121236 581612 121242 581664
rect 305730 581000 305736 581052
rect 305788 581040 305794 581052
rect 321554 581040 321560 581052
rect 305788 581012 321560 581040
rect 305788 581000 305794 581012
rect 321554 581000 321560 581012
rect 321612 581000 321618 581052
rect 218146 579640 218152 579692
rect 218204 579680 218210 579692
rect 237374 579680 237380 579692
rect 218204 579652 237380 579680
rect 218204 579640 218210 579652
rect 237374 579640 237380 579652
rect 237432 579640 237438 579692
rect 216674 576852 216680 576904
rect 216732 576892 216738 576904
rect 237374 576892 237380 576904
rect 216732 576864 237380 576892
rect 216732 576852 216738 576864
rect 237374 576852 237380 576864
rect 237432 576852 237438 576904
rect 148410 576784 148416 576836
rect 148468 576824 148474 576836
rect 149422 576824 149428 576836
rect 148468 576796 149428 576824
rect 148468 576784 148474 576796
rect 149422 576784 149428 576796
rect 149480 576784 149486 576836
rect 57146 575696 57152 575748
rect 57204 575736 57210 575748
rect 59906 575736 59912 575748
rect 57204 575708 59912 575736
rect 57204 575696 57210 575708
rect 59906 575696 59912 575708
rect 59964 575696 59970 575748
rect 3786 575424 3792 575476
rect 3844 575464 3850 575476
rect 307110 575464 307116 575476
rect 3844 575436 307116 575464
rect 3844 575424 3850 575436
rect 307110 575424 307116 575436
rect 307168 575424 307174 575476
rect 145558 575356 145564 575408
rect 145616 575396 145622 575408
rect 214006 575396 214012 575408
rect 145616 575368 214012 575396
rect 145616 575356 145622 575368
rect 214006 575356 214012 575368
rect 214064 575396 214070 575408
rect 302878 575396 302884 575408
rect 214064 575368 302884 575396
rect 214064 575356 214070 575368
rect 302878 575356 302884 575368
rect 302936 575356 302942 575408
rect 57054 575288 57060 575340
rect 57112 575328 57118 575340
rect 62114 575328 62120 575340
rect 57112 575300 62120 575328
rect 57112 575288 57118 575300
rect 62114 575288 62120 575300
rect 62172 575288 62178 575340
rect 106274 575288 106280 575340
rect 106332 575328 106338 575340
rect 124674 575328 124680 575340
rect 106332 575300 124680 575328
rect 106332 575288 106338 575300
rect 124674 575288 124680 575300
rect 124732 575288 124738 575340
rect 149330 575288 149336 575340
rect 149388 575328 149394 575340
rect 151814 575328 151820 575340
rect 149388 575300 151820 575328
rect 149388 575288 149394 575300
rect 151814 575288 151820 575300
rect 151872 575288 151878 575340
rect 289814 575288 289820 575340
rect 289872 575328 289878 575340
rect 314010 575328 314016 575340
rect 289872 575300 314016 575328
rect 289872 575288 289878 575300
rect 314010 575288 314016 575300
rect 314068 575288 314074 575340
rect 99558 575220 99564 575272
rect 99616 575260 99622 575272
rect 122282 575260 122288 575272
rect 99616 575232 122288 575260
rect 99616 575220 99622 575232
rect 122282 575220 122288 575232
rect 122340 575220 122346 575272
rect 149698 575220 149704 575272
rect 149756 575260 149762 575272
rect 154758 575260 154764 575272
rect 149756 575232 154764 575260
rect 149756 575220 149762 575232
rect 154758 575220 154764 575232
rect 154816 575220 154822 575272
rect 293954 575220 293960 575272
rect 294012 575260 294018 575272
rect 319622 575260 319628 575272
rect 294012 575232 319628 575260
rect 294012 575220 294018 575232
rect 319622 575220 319628 575232
rect 319680 575220 319686 575272
rect 98086 575152 98092 575204
rect 98144 575192 98150 575204
rect 120994 575192 121000 575204
rect 98144 575164 121000 575192
rect 98144 575152 98150 575164
rect 120994 575152 121000 575164
rect 121052 575152 121058 575204
rect 148594 575152 148600 575204
rect 148652 575192 148658 575204
rect 150526 575192 150532 575204
rect 148652 575164 150532 575192
rect 148652 575152 148658 575164
rect 150526 575152 150532 575164
rect 150584 575152 150590 575204
rect 288526 575152 288532 575204
rect 288584 575192 288590 575204
rect 316954 575192 316960 575204
rect 288584 575164 316960 575192
rect 288584 575152 288590 575164
rect 316954 575152 316960 575164
rect 317012 575152 317018 575204
rect 96798 575084 96804 575136
rect 96856 575124 96862 575136
rect 122834 575124 122840 575136
rect 96856 575096 122840 575124
rect 96856 575084 96862 575096
rect 122834 575084 122840 575096
rect 122892 575084 122898 575136
rect 288434 575084 288440 575136
rect 288492 575124 288498 575136
rect 316862 575124 316868 575136
rect 288492 575096 316868 575124
rect 288492 575084 288498 575096
rect 316862 575084 316868 575096
rect 316920 575084 316926 575136
rect 93854 575016 93860 575068
rect 93912 575056 93918 575068
rect 124490 575056 124496 575068
rect 93912 575028 124496 575056
rect 93912 575016 93918 575028
rect 124490 575016 124496 575028
rect 124548 575016 124554 575068
rect 147306 575016 147312 575068
rect 147364 575056 147370 575068
rect 156046 575056 156052 575068
rect 147364 575028 156052 575056
rect 147364 575016 147370 575028
rect 156046 575016 156052 575028
rect 156104 575016 156110 575068
rect 195238 575016 195244 575068
rect 195296 575056 195302 575068
rect 212810 575056 212816 575068
rect 195296 575028 212816 575056
rect 195296 575016 195302 575028
rect 212810 575016 212816 575028
rect 212868 575016 212874 575068
rect 287054 575016 287060 575068
rect 287112 575056 287118 575068
rect 317046 575056 317052 575068
rect 287112 575028 317052 575056
rect 287112 575016 287118 575028
rect 317046 575016 317052 575028
rect 317104 575016 317110 575068
rect 58894 574948 58900 575000
rect 58952 574988 58958 575000
rect 74534 574988 74540 575000
rect 58952 574960 74540 574988
rect 58952 574948 58958 574960
rect 74534 574948 74540 574960
rect 74592 574948 74598 575000
rect 86954 574948 86960 575000
rect 87012 574988 87018 575000
rect 121454 574988 121460 575000
rect 87012 574960 121460 574988
rect 87012 574948 87018 574960
rect 121454 574948 121460 574960
rect 121512 574948 121518 575000
rect 149790 574948 149796 575000
rect 149848 574988 149854 575000
rect 160278 574988 160284 575000
rect 149848 574960 160284 574988
rect 149848 574948 149854 574960
rect 160278 574948 160284 574960
rect 160336 574948 160342 575000
rect 164326 574948 164332 575000
rect 164384 574988 164390 575000
rect 212626 574988 212632 575000
rect 164384 574960 212632 574988
rect 164384 574948 164390 574960
rect 212626 574948 212632 574960
rect 212684 574948 212690 575000
rect 260834 574948 260840 575000
rect 260892 574988 260898 575000
rect 319438 574988 319444 575000
rect 260892 574960 319444 574988
rect 260892 574948 260898 574960
rect 319438 574948 319444 574960
rect 319496 574948 319502 575000
rect 54846 574880 54852 574932
rect 54904 574920 54910 574932
rect 78674 574920 78680 574932
rect 54904 574892 78680 574920
rect 54904 574880 54910 574892
rect 78674 574880 78680 574892
rect 78732 574880 78738 574932
rect 87046 574880 87052 574932
rect 87104 574920 87110 574932
rect 124582 574920 124588 574932
rect 87104 574892 124588 574920
rect 87104 574880 87110 574892
rect 124582 574880 124588 574892
rect 124640 574880 124646 574932
rect 126974 574880 126980 574932
rect 127032 574920 127038 574932
rect 211798 574920 211804 574932
rect 127032 574892 211804 574920
rect 127032 574880 127038 574892
rect 211798 574880 211804 574892
rect 211856 574880 211862 574932
rect 227714 574880 227720 574932
rect 227772 574920 227778 574932
rect 300946 574920 300952 574932
rect 227772 574892 300952 574920
rect 227772 574880 227778 574892
rect 300946 574880 300952 574892
rect 301004 574880 301010 574932
rect 58710 574812 58716 574864
rect 58768 574852 58774 574864
rect 67634 574852 67640 574864
rect 58768 574824 67640 574852
rect 58768 574812 58774 574824
rect 67634 574812 67640 574824
rect 67692 574812 67698 574864
rect 69014 574812 69020 574864
rect 69072 574852 69078 574864
rect 122190 574852 122196 574864
rect 69072 574824 122196 574852
rect 69072 574812 69078 574824
rect 122190 574812 122196 574824
rect 122248 574812 122254 574864
rect 148778 574812 148784 574864
rect 148836 574852 148842 574864
rect 161474 574852 161480 574864
rect 148836 574824 161480 574852
rect 148836 574812 148842 574824
rect 161474 574812 161480 574824
rect 161532 574812 161538 574864
rect 183646 574812 183652 574864
rect 183704 574852 183710 574864
rect 301038 574852 301044 574864
rect 183704 574824 301044 574852
rect 183704 574812 183710 574824
rect 301038 574812 301044 574824
rect 301096 574812 301102 574864
rect 63494 574744 63500 574796
rect 63552 574784 63558 574796
rect 123570 574784 123576 574796
rect 63552 574756 123576 574784
rect 63552 574744 63558 574756
rect 123570 574744 123576 574756
rect 123628 574744 123634 574796
rect 148870 574744 148876 574796
rect 148928 574784 148934 574796
rect 164234 574784 164240 574796
rect 148928 574756 164240 574784
rect 148928 574744 148934 574756
rect 164234 574744 164240 574756
rect 164292 574744 164298 574796
rect 179414 574744 179420 574796
rect 179472 574784 179478 574796
rect 300854 574784 300860 574796
rect 179472 574756 300860 574784
rect 179472 574744 179478 574756
rect 300854 574744 300860 574756
rect 300912 574744 300918 574796
rect 291194 574676 291200 574728
rect 291252 574716 291258 574728
rect 314102 574716 314108 574728
rect 291252 574688 314108 574716
rect 291252 574676 291258 574688
rect 314102 574676 314108 574688
rect 314160 574676 314166 574728
rect 119338 574608 119344 574660
rect 119396 574648 119402 574660
rect 123386 574648 123392 574660
rect 119396 574620 123392 574648
rect 119396 574608 119402 574620
rect 123386 574608 123392 574620
rect 123444 574608 123450 574660
rect 296898 574608 296904 574660
rect 296956 574648 296962 574660
rect 319530 574648 319536 574660
rect 296956 574620 319536 574648
rect 296956 574608 296962 574620
rect 319530 574608 319536 574620
rect 319588 574608 319594 574660
rect 57422 574268 57428 574320
rect 57480 574308 57486 574320
rect 60734 574308 60740 574320
rect 57480 574280 60740 574308
rect 57480 574268 57486 574280
rect 60734 574268 60740 574280
rect 60792 574268 60798 574320
rect 302878 574064 302884 574116
rect 302936 574104 302942 574116
rect 303338 574104 303344 574116
rect 302936 574076 303344 574104
rect 302936 574064 302942 574076
rect 303338 574064 303344 574076
rect 303396 574064 303402 574116
rect 111886 573588 111892 573640
rect 111944 573628 111950 573640
rect 123018 573628 123024 573640
rect 111944 573600 123024 573628
rect 111944 573588 111950 573600
rect 123018 573588 123024 573600
rect 123076 573588 123082 573640
rect 229094 573588 229100 573640
rect 229152 573628 229158 573640
rect 303062 573628 303068 573640
rect 229152 573600 303068 573628
rect 229152 573588 229158 573600
rect 303062 573588 303068 573600
rect 303120 573588 303126 573640
rect 59078 573520 59084 573572
rect 59136 573560 59142 573572
rect 92566 573560 92572 573572
rect 59136 573532 92572 573560
rect 59136 573520 59142 573532
rect 92566 573520 92572 573532
rect 92624 573520 92630 573572
rect 122834 573520 122840 573572
rect 122892 573560 122898 573572
rect 211430 573560 211436 573572
rect 122892 573532 211436 573560
rect 122892 573520 122898 573532
rect 211430 573520 211436 573532
rect 211488 573520 211494 573572
rect 245654 573520 245660 573572
rect 245712 573560 245718 573572
rect 322566 573560 322572 573572
rect 245712 573532 322572 573560
rect 245712 573520 245718 573532
rect 322566 573520 322572 573532
rect 322624 573520 322630 573572
rect 57514 573452 57520 573504
rect 57572 573492 57578 573504
rect 82906 573492 82912 573504
rect 57572 573464 82912 573492
rect 57572 573452 57578 573464
rect 82906 573452 82912 573464
rect 82964 573452 82970 573504
rect 84194 573452 84200 573504
rect 84252 573492 84258 573504
rect 122098 573492 122104 573504
rect 84252 573464 122104 573492
rect 84252 573452 84258 573464
rect 122098 573452 122104 573464
rect 122156 573452 122162 573504
rect 201678 573452 201684 573504
rect 201736 573492 201742 573504
rect 302234 573492 302240 573504
rect 201736 573464 302240 573492
rect 201736 573452 201742 573464
rect 302234 573452 302240 573464
rect 302292 573452 302298 573504
rect 65058 573384 65064 573436
rect 65116 573424 65122 573436
rect 122006 573424 122012 573436
rect 65116 573396 122012 573424
rect 65116 573384 65122 573396
rect 122006 573384 122012 573396
rect 122064 573384 122070 573436
rect 149606 573384 149612 573436
rect 149664 573424 149670 573436
rect 158714 573424 158720 573436
rect 149664 573396 158720 573424
rect 149664 573384 149670 573396
rect 158714 573384 158720 573396
rect 158772 573384 158778 573436
rect 179506 573384 179512 573436
rect 179564 573424 179570 573436
rect 301590 573424 301596 573436
rect 179564 573396 301596 573424
rect 179564 573384 179570 573396
rect 301590 573384 301596 573396
rect 301648 573384 301654 573436
rect 3510 573316 3516 573368
rect 3568 573356 3574 573368
rect 324038 573356 324044 573368
rect 3568 573328 324044 573356
rect 3568 573316 3574 573328
rect 324038 573316 324044 573328
rect 324096 573316 324102 573368
rect 147122 572704 147128 572756
rect 147180 572744 147186 572756
rect 151078 572744 151084 572756
rect 147180 572716 151084 572744
rect 147180 572704 147186 572716
rect 151078 572704 151084 572716
rect 151136 572704 151142 572756
rect 62758 572500 62764 572552
rect 62816 572540 62822 572552
rect 65150 572540 65156 572552
rect 62816 572512 65156 572540
rect 62816 572500 62822 572512
rect 65150 572500 65156 572512
rect 65208 572500 65214 572552
rect 161566 572432 161572 572484
rect 161624 572472 161630 572484
rect 178034 572472 178040 572484
rect 161624 572444 178040 572472
rect 161624 572432 161630 572444
rect 178034 572432 178040 572444
rect 178092 572432 178098 572484
rect 163038 572364 163044 572416
rect 163096 572404 163102 572416
rect 183830 572404 183836 572416
rect 163096 572376 183836 572404
rect 163096 572364 163102 572376
rect 183830 572364 183836 572376
rect 183888 572364 183894 572416
rect 235534 572364 235540 572416
rect 235592 572404 235598 572416
rect 248414 572404 248420 572416
rect 235592 572376 248420 572404
rect 235592 572364 235598 572376
rect 248414 572364 248420 572376
rect 248472 572364 248478 572416
rect 143534 572296 143540 572348
rect 143592 572336 143598 572348
rect 166442 572336 166448 572348
rect 143592 572308 166448 572336
rect 143592 572296 143598 572308
rect 166442 572296 166448 572308
rect 166500 572296 166506 572348
rect 169846 572296 169852 572348
rect 169904 572336 169910 572348
rect 175458 572336 175464 572348
rect 169904 572308 175464 572336
rect 169904 572296 169910 572308
rect 175458 572296 175464 572308
rect 175516 572296 175522 572348
rect 197998 572296 198004 572348
rect 198056 572336 198062 572348
rect 201494 572336 201500 572348
rect 198056 572308 201500 572336
rect 198056 572296 198062 572308
rect 201494 572296 201500 572308
rect 201552 572296 201558 572348
rect 220814 572296 220820 572348
rect 220872 572336 220878 572348
rect 240042 572336 240048 572348
rect 220872 572308 240048 572336
rect 220872 572296 220878 572308
rect 240042 572296 240048 572308
rect 240100 572296 240106 572348
rect 249058 572296 249064 572348
rect 249116 572336 249122 572348
rect 271598 572336 271604 572348
rect 249116 572308 271604 572336
rect 249116 572296 249122 572308
rect 271598 572296 271604 572308
rect 271656 572296 271662 572348
rect 154666 572228 154672 572280
rect 154724 572268 154730 572280
rect 181254 572268 181260 572280
rect 154724 572240 181260 572268
rect 154724 572228 154730 572240
rect 181254 572228 181260 572240
rect 181312 572228 181318 572280
rect 230474 572228 230480 572280
rect 230532 572268 230538 572280
rect 260006 572268 260012 572280
rect 230532 572240 260012 572268
rect 230532 572228 230538 572240
rect 260006 572228 260012 572240
rect 260064 572228 260070 572280
rect 70946 572160 70952 572212
rect 71004 572200 71010 572212
rect 86218 572200 86224 572212
rect 71004 572172 86224 572200
rect 71004 572160 71010 572172
rect 86218 572160 86224 572172
rect 86276 572160 86282 572212
rect 94130 572160 94136 572212
rect 94188 572200 94194 572212
rect 104894 572200 104900 572212
rect 94188 572172 104900 572200
rect 94188 572160 94194 572172
rect 104894 572160 104900 572172
rect 104952 572160 104958 572212
rect 158806 572160 158812 572212
rect 158864 572200 158870 572212
rect 192846 572200 192852 572212
rect 158864 572172 192852 572200
rect 158864 572160 158870 572172
rect 192846 572160 192852 572172
rect 192904 572160 192910 572212
rect 227806 572160 227812 572212
rect 227864 572200 227870 572212
rect 265802 572200 265808 572212
rect 227864 572172 265808 572200
rect 227864 572160 227870 572172
rect 265802 572160 265808 572172
rect 265860 572160 265866 572212
rect 273898 572160 273904 572212
rect 273956 572200 273962 572212
rect 283190 572200 283196 572212
rect 273956 572172 283196 572200
rect 273956 572160 273962 572172
rect 283190 572160 283196 572172
rect 283248 572160 283254 572212
rect 287698 572160 287704 572212
rect 287756 572200 287762 572212
rect 300578 572200 300584 572212
rect 287756 572172 300584 572200
rect 287756 572160 287762 572172
rect 300578 572160 300584 572172
rect 300636 572160 300642 572212
rect 74626 572092 74632 572144
rect 74684 572132 74690 572144
rect 97350 572132 97356 572144
rect 74684 572104 97356 572132
rect 74684 572092 74690 572104
rect 97350 572092 97356 572104
rect 97408 572092 97414 572144
rect 99926 572092 99932 572144
rect 99984 572132 99990 572144
rect 115198 572132 115204 572144
rect 99984 572104 115204 572132
rect 99984 572092 99990 572104
rect 115198 572092 115204 572104
rect 115256 572092 115262 572144
rect 129734 572092 129740 572144
rect 129792 572132 129798 572144
rect 163866 572132 163872 572144
rect 129792 572104 163872 572132
rect 129792 572092 129798 572104
rect 163866 572092 163872 572104
rect 163924 572092 163930 572144
rect 173894 572092 173900 572144
rect 173952 572132 173958 572144
rect 189626 572132 189632 572144
rect 173952 572104 189632 572132
rect 173952 572092 173958 572104
rect 189626 572092 189632 572104
rect 189684 572092 189690 572144
rect 193858 572092 193864 572144
rect 193916 572132 193922 572144
rect 210234 572132 210240 572144
rect 193916 572104 210240 572132
rect 193916 572092 193922 572104
rect 210234 572092 210240 572104
rect 210292 572092 210298 572144
rect 231946 572092 231952 572144
rect 232004 572132 232010 572144
rect 279970 572132 279976 572144
rect 232004 572104 279976 572132
rect 232004 572092 232010 572104
rect 279970 572092 279976 572104
rect 280028 572092 280034 572144
rect 280798 572092 280804 572144
rect 280856 572132 280862 572144
rect 297358 572132 297364 572144
rect 280856 572104 297364 572132
rect 280856 572092 280862 572104
rect 297358 572092 297364 572104
rect 297416 572092 297422 572144
rect 57330 572024 57336 572076
rect 57388 572064 57394 572076
rect 79318 572064 79324 572076
rect 57388 572036 79324 572064
rect 57388 572024 57394 572036
rect 79318 572024 79324 572036
rect 79376 572024 79382 572076
rect 85758 572024 85764 572076
rect 85816 572064 85822 572076
rect 108298 572064 108304 572076
rect 85816 572036 108304 572064
rect 85816 572024 85822 572036
rect 108298 572024 108304 572036
rect 108356 572024 108362 572076
rect 110414 572024 110420 572076
rect 110472 572064 110478 572076
rect 121178 572064 121184 572076
rect 110472 572036 121184 572064
rect 110472 572024 110478 572036
rect 121178 572024 121184 572036
rect 121236 572024 121242 572076
rect 132586 572024 132592 572076
rect 132644 572064 132650 572076
rect 187050 572064 187056 572076
rect 132644 572036 187056 572064
rect 132644 572024 132650 572036
rect 187050 572024 187056 572036
rect 187108 572024 187114 572076
rect 192478 572024 192484 572076
rect 192536 572064 192542 572076
rect 213270 572064 213276 572076
rect 192536 572036 213276 572064
rect 192536 572024 192542 572036
rect 213270 572024 213276 572036
rect 213328 572024 213334 572076
rect 219434 572024 219440 572076
rect 219492 572064 219498 572076
rect 268378 572064 268384 572076
rect 219492 572036 268384 572064
rect 219492 572024 219498 572036
rect 268378 572024 268384 572036
rect 268436 572024 268442 572076
rect 269114 572024 269120 572076
rect 269172 572064 269178 572076
rect 309962 572064 309968 572076
rect 269172 572036 309968 572064
rect 269172 572024 269178 572036
rect 309962 572024 309968 572036
rect 310020 572024 310026 572076
rect 59998 571956 60004 572008
rect 60056 571996 60062 572008
rect 71038 571996 71044 572008
rect 60056 571968 71044 571996
rect 60056 571956 60062 571968
rect 71038 571956 71044 571968
rect 71096 571956 71102 572008
rect 79962 571956 79968 572008
rect 80020 571996 80026 572008
rect 114738 571996 114744 572008
rect 80020 571968 114744 571996
rect 80020 571956 80026 571968
rect 114738 571956 114744 571968
rect 114796 571956 114802 572008
rect 133966 571956 133972 572008
rect 134024 571996 134030 572008
rect 207014 571996 207020 572008
rect 134024 571968 207020 571996
rect 134024 571956 134030 571968
rect 207014 571956 207020 571968
rect 207072 571956 207078 572008
rect 222286 571956 222292 572008
rect 222344 571996 222350 572008
rect 274174 571996 274180 572008
rect 222344 571968 274180 571996
rect 222344 571956 222350 571968
rect 274174 571956 274180 571968
rect 274232 571956 274238 572008
rect 280154 571956 280160 572008
rect 280212 571996 280218 572008
rect 322474 571996 322480 572008
rect 280212 571968 322480 571996
rect 280212 571956 280218 571968
rect 322474 571956 322480 571968
rect 322532 571956 322538 572008
rect 246298 571480 246304 571532
rect 246356 571520 246362 571532
rect 250990 571520 250996 571532
rect 246356 571492 250996 571520
rect 246356 571480 246362 571492
rect 250990 571480 250996 571492
rect 251048 571480 251054 571532
rect 116670 571412 116676 571464
rect 116728 571452 116734 571464
rect 120534 571452 120540 571464
rect 116728 571424 120540 571452
rect 116728 571412 116734 571424
rect 120534 571412 120540 571424
rect 120592 571412 120598 571464
rect 71774 571344 71780 571396
rect 71832 571384 71838 571396
rect 74166 571384 74172 571396
rect 71832 571356 74172 571384
rect 71832 571344 71838 571356
rect 74166 571344 74172 571356
rect 74224 571344 74230 571396
rect 116578 571344 116584 571396
rect 116636 571384 116642 571396
rect 117314 571384 117320 571396
rect 116636 571356 117320 571384
rect 116636 571344 116642 571356
rect 117314 571344 117320 571356
rect 117372 571344 117378 571396
rect 150342 571344 150348 571396
rect 150400 571384 150406 571396
rect 151170 571384 151176 571396
rect 150400 571356 151176 571384
rect 150400 571344 150406 571356
rect 151170 571344 151176 571356
rect 151228 571344 151234 571396
rect 191098 571344 191104 571396
rect 191156 571384 191162 571396
rect 195422 571384 195428 571396
rect 191156 571356 195428 571384
rect 191156 571344 191162 571356
rect 195422 571344 195428 571356
rect 195480 571344 195486 571396
rect 200114 570800 200120 570852
rect 200172 570840 200178 570852
rect 239582 570840 239588 570852
rect 200172 570812 239588 570840
rect 200172 570800 200178 570812
rect 239582 570800 239588 570812
rect 239640 570800 239646 570852
rect 58802 570732 58808 570784
rect 58860 570772 58866 570784
rect 91094 570772 91100 570784
rect 58860 570744 91100 570772
rect 58860 570732 58866 570744
rect 91094 570732 91100 570744
rect 91152 570732 91158 570784
rect 91554 570732 91560 570784
rect 91612 570772 91618 570784
rect 96706 570772 96712 570784
rect 91612 570744 96712 570772
rect 91612 570732 91618 570744
rect 96706 570732 96712 570744
rect 96764 570732 96770 570784
rect 121454 570732 121460 570784
rect 121512 570772 121518 570784
rect 211154 570772 211160 570784
rect 121512 570744 211160 570772
rect 121512 570732 121518 570744
rect 211154 570732 211160 570744
rect 211212 570732 211218 570784
rect 215294 570732 215300 570784
rect 215352 570772 215358 570784
rect 301498 570772 301504 570784
rect 215352 570744 301504 570772
rect 215352 570732 215358 570744
rect 301498 570732 301504 570744
rect 301556 570732 301562 570784
rect 66346 570664 66352 570716
rect 66404 570704 66410 570716
rect 120718 570704 120724 570716
rect 66404 570676 120724 570704
rect 66404 570664 66410 570676
rect 120718 570664 120724 570676
rect 120776 570664 120782 570716
rect 180794 570664 180800 570716
rect 180852 570704 180858 570716
rect 301130 570704 301136 570716
rect 180852 570676 301136 570704
rect 180852 570664 180858 570676
rect 301130 570664 301136 570676
rect 301188 570664 301194 570716
rect 10318 570596 10324 570648
rect 10376 570636 10382 570648
rect 321554 570636 321560 570648
rect 10376 570608 321560 570636
rect 10376 570596 10382 570608
rect 321554 570596 321560 570608
rect 321612 570596 321618 570648
rect 118694 569372 118700 569424
rect 118752 569412 118758 569424
rect 154850 569412 154856 569424
rect 118752 569384 154856 569412
rect 118752 569372 118758 569384
rect 154850 569372 154856 569384
rect 154908 569372 154914 569424
rect 191834 569372 191840 569424
rect 191892 569412 191898 569424
rect 238846 569412 238852 569424
rect 191892 569384 238852 569412
rect 191892 569372 191898 569384
rect 238846 569372 238852 569384
rect 238904 569372 238910 569424
rect 80054 569304 80060 569356
rect 80112 569344 80118 569356
rect 120810 569344 120816 569356
rect 80112 569316 120816 569344
rect 80112 569304 80118 569316
rect 120810 569304 120816 569316
rect 120868 569304 120874 569356
rect 157426 569304 157432 569356
rect 157484 569344 157490 569356
rect 213178 569344 213184 569356
rect 157484 569316 213184 569344
rect 157484 569304 157490 569316
rect 213178 569304 213184 569316
rect 213236 569304 213242 569356
rect 255314 569304 255320 569356
rect 255372 569344 255378 569356
rect 324774 569344 324780 569356
rect 255372 569316 324780 569344
rect 255372 569304 255378 569316
rect 324774 569304 324780 569316
rect 324832 569304 324838 569356
rect 58526 569236 58532 569288
rect 58584 569276 58590 569288
rect 110506 569276 110512 569288
rect 58584 569248 110512 569276
rect 58584 569236 58590 569248
rect 110506 569236 110512 569248
rect 110564 569236 110570 569288
rect 142798 569236 142804 569288
rect 142856 569276 142862 569288
rect 213086 569276 213092 569288
rect 142856 569248 213092 569276
rect 142856 569236 142862 569248
rect 213086 569236 213092 569248
rect 213144 569236 213150 569288
rect 240134 569236 240140 569288
rect 240192 569276 240198 569288
rect 309778 569276 309784 569288
rect 240192 569248 309784 569276
rect 240192 569236 240198 569248
rect 309778 569236 309784 569248
rect 309836 569236 309842 569288
rect 67726 569168 67732 569220
rect 67784 569208 67790 569220
rect 123110 569208 123116 569220
rect 67784 569180 123116 569208
rect 67784 569168 67790 569180
rect 123110 569168 123116 569180
rect 123168 569168 123174 569220
rect 147398 569168 147404 569220
rect 147456 569208 147462 569220
rect 165614 569208 165620 569220
rect 147456 569180 165620 569208
rect 147456 569168 147462 569180
rect 165614 569168 165620 569180
rect 165672 569168 165678 569220
rect 186314 569168 186320 569220
rect 186372 569208 186378 569220
rect 301406 569208 301412 569220
rect 186372 569180 301412 569208
rect 186372 569168 186378 569180
rect 301406 569168 301412 569180
rect 301464 569168 301470 569220
rect 176654 568012 176660 568064
rect 176712 568052 176718 568064
rect 235442 568052 235448 568064
rect 176712 568024 235448 568052
rect 176712 568012 176718 568024
rect 235442 568012 235448 568024
rect 235500 568012 235506 568064
rect 59446 567944 59452 567996
rect 59504 567984 59510 567996
rect 75914 567984 75920 567996
rect 59504 567956 75920 567984
rect 59504 567944 59510 567956
rect 75914 567944 75920 567956
rect 75972 567944 75978 567996
rect 128354 567944 128360 567996
rect 128412 567984 128418 567996
rect 211338 567984 211344 567996
rect 128412 567956 211344 567984
rect 128412 567944 128418 567956
rect 211338 567944 211344 567956
rect 211396 567944 211402 567996
rect 69106 567876 69112 567928
rect 69164 567916 69170 567928
rect 114554 567916 114560 567928
rect 69164 567888 114560 567916
rect 69164 567876 69170 567888
rect 114554 567876 114560 567888
rect 114612 567876 114618 567928
rect 125686 567876 125692 567928
rect 125744 567916 125750 567928
rect 211246 567916 211252 567928
rect 125744 567888 211252 567916
rect 125744 567876 125750 567888
rect 211246 567876 211252 567888
rect 211304 567876 211310 567928
rect 244458 567876 244464 567928
rect 244516 567916 244522 567928
rect 318150 567916 318156 567928
rect 244516 567888 318156 567916
rect 244516 567876 244522 567888
rect 318150 567876 318156 567888
rect 318208 567876 318214 567928
rect 70394 567808 70400 567860
rect 70452 567848 70458 567860
rect 121822 567848 121828 567860
rect 70452 567820 121828 567848
rect 70452 567808 70458 567820
rect 121822 567808 121828 567820
rect 121880 567808 121886 567860
rect 194594 567808 194600 567860
rect 194652 567848 194658 567860
rect 302970 567848 302976 567860
rect 194652 567820 302976 567848
rect 194652 567808 194658 567820
rect 302970 567808 302976 567820
rect 303028 567808 303034 567860
rect 267734 567196 267740 567248
rect 267792 567236 267798 567248
rect 321554 567236 321560 567248
rect 267792 567208 321560 567236
rect 267792 567196 267798 567208
rect 321554 567196 321560 567208
rect 321612 567196 321618 567248
rect 198734 566652 198740 566704
rect 198792 566692 198798 566704
rect 239490 566692 239496 566704
rect 198792 566664 239496 566692
rect 198792 566652 198798 566664
rect 239490 566652 239496 566664
rect 239548 566652 239554 566704
rect 269206 566652 269212 566704
rect 269264 566692 269270 566704
rect 311342 566692 311348 566704
rect 269264 566664 311348 566692
rect 269264 566652 269270 566664
rect 311342 566652 311348 566664
rect 311400 566652 311406 566704
rect 57238 566584 57244 566636
rect 57296 566624 57302 566636
rect 89714 566624 89720 566636
rect 57296 566596 89720 566624
rect 57296 566584 57302 566596
rect 89714 566584 89720 566596
rect 89772 566584 89778 566636
rect 123018 566584 123024 566636
rect 123076 566624 123082 566636
rect 211706 566624 211712 566636
rect 123076 566596 211712 566624
rect 123076 566584 123082 566596
rect 211706 566584 211712 566596
rect 211764 566584 211770 566636
rect 247034 566584 247040 566636
rect 247092 566624 247098 566636
rect 324866 566624 324872 566636
rect 247092 566596 324872 566624
rect 247092 566584 247098 566596
rect 324866 566584 324872 566596
rect 324924 566584 324930 566636
rect 85574 566516 85580 566568
rect 85632 566556 85638 566568
rect 121730 566556 121736 566568
rect 85632 566528 121736 566556
rect 85632 566516 85638 566528
rect 121730 566516 121736 566528
rect 121788 566516 121794 566568
rect 184934 566516 184940 566568
rect 184992 566556 184998 566568
rect 294046 566556 294052 566568
rect 184992 566528 294052 566556
rect 184992 566516 184998 566528
rect 294046 566516 294052 566528
rect 294104 566516 294110 566568
rect 63586 566448 63592 566500
rect 63644 566488 63650 566500
rect 122926 566488 122932 566500
rect 63644 566460 122932 566488
rect 63644 566448 63650 566460
rect 122926 566448 122932 566460
rect 122984 566448 122990 566500
rect 147030 566448 147036 566500
rect 147088 566488 147094 566500
rect 168374 566488 168380 566500
rect 147088 566460 168380 566488
rect 147088 566448 147094 566460
rect 168374 566448 168380 566460
rect 168432 566448 168438 566500
rect 187694 566448 187700 566500
rect 187752 566488 187758 566500
rect 302326 566488 302332 566500
rect 187752 566460 302332 566488
rect 187752 566448 187758 566460
rect 302326 566448 302332 566460
rect 302384 566448 302390 566500
rect 176746 565292 176752 565344
rect 176804 565332 176810 565344
rect 244274 565332 244280 565344
rect 176804 565304 244280 565332
rect 176804 565292 176810 565304
rect 244274 565292 244280 565304
rect 244332 565292 244338 565344
rect 129826 565224 129832 565276
rect 129884 565264 129890 565276
rect 212718 565264 212724 565276
rect 129884 565236 212724 565264
rect 129884 565224 129890 565236
rect 212718 565224 212724 565236
rect 212776 565224 212782 565276
rect 274634 565224 274640 565276
rect 274692 565264 274698 565276
rect 316770 565264 316776 565276
rect 274692 565236 316776 565264
rect 274692 565224 274698 565236
rect 316770 565224 316776 565236
rect 316828 565224 316834 565276
rect 88518 565156 88524 565208
rect 88576 565196 88582 565208
rect 104986 565196 104992 565208
rect 88576 565168 104992 565196
rect 88576 565156 88582 565168
rect 104986 565156 104992 565168
rect 105044 565156 105050 565208
rect 168466 565156 168472 565208
rect 168524 565196 168530 565208
rect 210694 565196 210700 565208
rect 168524 565168 210700 565196
rect 168524 565156 168530 565168
rect 210694 565156 210700 565168
rect 210752 565156 210758 565208
rect 211154 565156 211160 565208
rect 211212 565196 211218 565208
rect 301314 565196 301320 565208
rect 211212 565168 301320 565196
rect 211212 565156 211218 565168
rect 301314 565156 301320 565168
rect 301372 565156 301378 565208
rect 64966 565088 64972 565140
rect 65024 565128 65030 565140
rect 123202 565128 123208 565140
rect 65024 565100 123208 565128
rect 65024 565088 65030 565100
rect 123202 565088 123208 565100
rect 123260 565088 123266 565140
rect 195974 565088 195980 565140
rect 196032 565128 196038 565140
rect 302510 565128 302516 565140
rect 196032 565100 302516 565128
rect 196032 565088 196038 565100
rect 302510 565088 302516 565100
rect 302568 565088 302574 565140
rect 136726 563864 136732 563916
rect 136784 563904 136790 563916
rect 210786 563904 210792 563916
rect 136784 563876 210792 563904
rect 136784 563864 136790 563876
rect 210786 563864 210792 563876
rect 210844 563864 210850 563916
rect 263594 563864 263600 563916
rect 263652 563904 263658 563916
rect 307018 563904 307024 563916
rect 263652 563876 307024 563904
rect 263652 563864 263658 563876
rect 307018 563864 307024 563876
rect 307076 563864 307082 563916
rect 81434 563796 81440 563848
rect 81492 563836 81498 563848
rect 89806 563836 89812 563848
rect 81492 563808 89812 563836
rect 81492 563796 81498 563808
rect 89806 563796 89812 563808
rect 89864 563796 89870 563848
rect 151998 563796 152004 563848
rect 152056 563836 152062 563848
rect 212994 563836 213000 563848
rect 152056 563808 213000 563836
rect 152056 563796 152062 563808
rect 212994 563796 213000 563808
rect 213052 563796 213058 563848
rect 273254 563796 273260 563848
rect 273312 563836 273318 563848
rect 322382 563836 322388 563848
rect 273312 563808 322388 563836
rect 273312 563796 273318 563808
rect 322382 563796 322388 563808
rect 322440 563796 322446 563848
rect 59538 563728 59544 563780
rect 59596 563768 59602 563780
rect 100754 563768 100760 563780
rect 59596 563740 100760 563768
rect 59596 563728 59602 563740
rect 100754 563728 100760 563740
rect 100812 563728 100818 563780
rect 210050 563728 210056 563780
rect 210108 563768 210114 563780
rect 302694 563768 302700 563780
rect 210108 563740 302700 563768
rect 210108 563728 210114 563740
rect 302694 563728 302700 563740
rect 302752 563728 302758 563780
rect 78766 563660 78772 563712
rect 78824 563700 78830 563712
rect 123478 563700 123484 563712
rect 78824 563672 123484 563700
rect 78824 563660 78830 563672
rect 123478 563660 123484 563672
rect 123536 563660 123542 563712
rect 186406 563660 186412 563712
rect 186464 563700 186470 563712
rect 302418 563700 302424 563712
rect 186464 563672 302424 563700
rect 186464 563660 186470 563672
rect 302418 563660 302424 563672
rect 302476 563660 302482 563712
rect 204346 562436 204352 562488
rect 204404 562476 204410 562488
rect 239398 562476 239404 562488
rect 204404 562448 239404 562476
rect 204404 562436 204410 562448
rect 239398 562436 239404 562448
rect 239456 562436 239462 562488
rect 146938 562368 146944 562420
rect 146996 562408 147002 562420
rect 212534 562408 212540 562420
rect 146996 562380 212540 562408
rect 146996 562368 147002 562380
rect 212534 562368 212540 562380
rect 212592 562368 212598 562420
rect 58986 562300 58992 562352
rect 59044 562340 59050 562352
rect 102226 562340 102232 562352
rect 59044 562312 102232 562340
rect 59044 562300 59050 562312
rect 102226 562300 102232 562312
rect 102284 562300 102290 562352
rect 189074 562300 189080 562352
rect 189132 562340 189138 562352
rect 288618 562340 288624 562352
rect 189132 562312 288624 562340
rect 189132 562300 189138 562312
rect 288618 562300 288624 562312
rect 288676 562300 288682 562352
rect 4798 561688 4804 561740
rect 4856 561728 4862 561740
rect 321554 561728 321560 561740
rect 4856 561700 321560 561728
rect 4856 561688 4862 561700
rect 321554 561688 321560 561700
rect 321612 561688 321618 561740
rect 178034 561144 178040 561196
rect 178092 561184 178098 561196
rect 233878 561184 233884 561196
rect 178092 561156 233884 561184
rect 178092 561144 178098 561156
rect 233878 561144 233884 561156
rect 233936 561144 233942 561196
rect 73246 561076 73252 561128
rect 73304 561116 73310 561128
rect 107654 561116 107660 561128
rect 73304 561088 107660 561116
rect 73304 561076 73310 561088
rect 107654 561076 107660 561088
rect 107712 561076 107718 561128
rect 187786 561076 187792 561128
rect 187844 561116 187850 561128
rect 253934 561116 253940 561128
rect 187844 561088 253940 561116
rect 187844 561076 187850 561088
rect 253934 561076 253940 561088
rect 253992 561076 253998 561128
rect 256786 561076 256792 561128
rect 256844 561116 256850 561128
rect 323946 561116 323952 561128
rect 256844 561088 323952 561116
rect 256844 561076 256850 561088
rect 323946 561076 323952 561088
rect 324004 561076 324010 561128
rect 80146 561008 80152 561060
rect 80204 561048 80210 561060
rect 121086 561048 121092 561060
rect 80204 561020 121092 561048
rect 80204 561008 80210 561020
rect 121086 561008 121092 561020
rect 121144 561008 121150 561060
rect 138014 561008 138020 561060
rect 138072 561048 138078 561060
rect 211614 561048 211620 561060
rect 138072 561020 211620 561048
rect 138072 561008 138078 561020
rect 211614 561008 211620 561020
rect 211672 561008 211678 561060
rect 249794 561008 249800 561060
rect 249852 561048 249858 561060
rect 323854 561048 323860 561060
rect 249852 561020 323860 561048
rect 249852 561008 249858 561020
rect 323854 561008 323860 561020
rect 323912 561008 323918 561060
rect 59262 560940 59268 560992
rect 59320 560980 59326 560992
rect 117314 560980 117320 560992
rect 59320 560952 117320 560980
rect 59320 560940 59326 560952
rect 117314 560940 117320 560952
rect 117372 560940 117378 560992
rect 147214 560940 147220 560992
rect 147272 560980 147278 560992
rect 173986 560980 173992 560992
rect 147272 560952 173992 560980
rect 147272 560940 147278 560952
rect 173986 560940 173992 560952
rect 174044 560940 174050 560992
rect 200206 560940 200212 560992
rect 200264 560980 200270 560992
rect 302786 560980 302792 560992
rect 200264 560952 302792 560980
rect 200264 560940 200270 560952
rect 302786 560940 302792 560952
rect 302844 560940 302850 560992
rect 207014 559716 207020 559768
rect 207072 559756 207078 559768
rect 220170 559756 220176 559768
rect 207072 559728 220176 559756
rect 207072 559716 207078 559728
rect 220170 559716 220176 559728
rect 220228 559716 220234 559768
rect 197354 559648 197360 559700
rect 197412 559688 197418 559700
rect 214742 559688 214748 559700
rect 197412 559660 214748 559688
rect 197412 559648 197418 559660
rect 214742 559648 214748 559660
rect 214800 559648 214806 559700
rect 259454 559648 259460 559700
rect 259512 559688 259518 559700
rect 305730 559688 305736 559700
rect 259512 559660 305736 559688
rect 259512 559648 259518 559660
rect 305730 559648 305736 559660
rect 305788 559648 305794 559700
rect 88426 559580 88432 559632
rect 88484 559620 88490 559632
rect 103514 559620 103520 559632
rect 88484 559592 103520 559620
rect 88484 559580 88490 559592
rect 103514 559580 103520 559592
rect 103572 559580 103578 559632
rect 127066 559580 127072 559632
rect 127124 559620 127130 559632
rect 204254 559620 204260 559632
rect 127124 559592 204260 559620
rect 127124 559580 127130 559592
rect 204254 559580 204260 559592
rect 204312 559580 204318 559632
rect 216766 559580 216772 559632
rect 216824 559620 216830 559632
rect 273898 559620 273904 559632
rect 216824 559592 273904 559620
rect 216824 559580 216830 559592
rect 273898 559580 273904 559592
rect 273956 559580 273962 559632
rect 59170 559512 59176 559564
rect 59228 559552 59234 559564
rect 107654 559552 107660 559564
rect 59228 559524 107660 559552
rect 59228 559512 59234 559524
rect 107654 559512 107660 559524
rect 107712 559512 107718 559564
rect 182174 559512 182180 559564
rect 182232 559552 182238 559564
rect 300670 559552 300676 559564
rect 182232 559524 300676 559552
rect 182232 559512 182238 559524
rect 300670 559512 300676 559524
rect 300728 559512 300734 559564
rect 40034 558832 40040 558884
rect 40092 558872 40098 558884
rect 321554 558872 321560 558884
rect 40092 558844 321560 558872
rect 40092 558832 40098 558844
rect 321554 558832 321560 558844
rect 321612 558832 321618 558884
rect 281534 558288 281540 558340
rect 281592 558328 281598 558340
rect 304258 558328 304264 558340
rect 281592 558300 304264 558328
rect 281592 558288 281598 558300
rect 304258 558288 304264 558300
rect 304316 558288 304322 558340
rect 190454 558220 190460 558272
rect 190512 558260 190518 558272
rect 222838 558260 222844 558272
rect 190512 558232 222844 558260
rect 190512 558220 190518 558232
rect 222838 558220 222844 558232
rect 222896 558220 222902 558272
rect 242894 558220 242900 558272
rect 242952 558260 242958 558272
rect 320910 558260 320916 558272
rect 242952 558232 320916 558260
rect 242952 558220 242958 558232
rect 320910 558220 320916 558232
rect 320968 558220 320974 558272
rect 67818 558152 67824 558204
rect 67876 558192 67882 558204
rect 107746 558192 107752 558204
rect 67876 558164 107752 558192
rect 67876 558152 67882 558164
rect 107746 558152 107752 558164
rect 107804 558152 107810 558204
rect 133138 558152 133144 558204
rect 133196 558192 133202 558204
rect 198826 558192 198832 558204
rect 133196 558164 198832 558192
rect 133196 558152 133202 558164
rect 198826 558152 198832 558164
rect 198884 558152 198890 558204
rect 205634 558152 205640 558204
rect 205692 558192 205698 558204
rect 285674 558192 285680 558204
rect 205692 558164 285680 558192
rect 205692 558152 205698 558164
rect 285674 558152 285680 558164
rect 285732 558152 285738 558204
rect 199194 556996 199200 557048
rect 199252 557036 199258 557048
rect 216122 557036 216128 557048
rect 199252 557008 216128 557036
rect 199252 556996 199258 557008
rect 216122 556996 216128 557008
rect 216180 556996 216186 557048
rect 76006 556928 76012 556980
rect 76064 556968 76070 556980
rect 86770 556968 86776 556980
rect 76064 556940 86776 556968
rect 76064 556928 76070 556940
rect 86770 556928 86776 556940
rect 86828 556928 86834 556980
rect 206370 556928 206376 556980
rect 206428 556968 206434 556980
rect 262214 556968 262220 556980
rect 206428 556940 262220 556968
rect 206428 556928 206434 556940
rect 262214 556928 262220 556940
rect 262272 556928 262278 556980
rect 266538 556928 266544 556980
rect 266596 556968 266602 556980
rect 322290 556968 322296 556980
rect 266596 556940 322296 556968
rect 266596 556928 266602 556940
rect 322290 556928 322296 556940
rect 322348 556928 322354 556980
rect 62206 556860 62212 556912
rect 62264 556900 62270 556912
rect 109678 556900 109684 556912
rect 62264 556872 109684 556900
rect 62264 556860 62270 556872
rect 109678 556860 109684 556872
rect 109736 556860 109742 556912
rect 124674 556860 124680 556912
rect 124732 556900 124738 556912
rect 210970 556900 210976 556912
rect 124732 556872 210976 556900
rect 124732 556860 124738 556872
rect 210970 556860 210976 556872
rect 211028 556860 211034 556912
rect 250070 556860 250076 556912
rect 250128 556900 250134 556912
rect 314194 556900 314200 556912
rect 250128 556872 314200 556900
rect 250128 556860 250134 556872
rect 314194 556860 314200 556872
rect 314252 556860 314258 556912
rect 71682 556792 71688 556844
rect 71740 556832 71746 556844
rect 121638 556832 121644 556844
rect 71740 556804 121644 556832
rect 71740 556792 71746 556804
rect 121638 556792 121644 556804
rect 121696 556792 121702 556844
rect 179138 556792 179144 556844
rect 179196 556832 179202 556844
rect 291286 556832 291292 556844
rect 179196 556804 291292 556832
rect 179196 556792 179202 556804
rect 291286 556792 291292 556804
rect 291344 556792 291350 556844
rect 215754 556180 215760 556232
rect 215812 556220 215818 556232
rect 217410 556220 217416 556232
rect 215812 556192 217416 556220
rect 215812 556180 215818 556192
rect 217410 556180 217416 556192
rect 217468 556180 217474 556232
rect 125594 556044 125600 556096
rect 125652 556084 125658 556096
rect 126882 556084 126888 556096
rect 125652 556056 126888 556084
rect 125652 556044 125658 556056
rect 126882 556044 126888 556056
rect 126940 556044 126946 556096
rect 193490 555704 193496 555756
rect 193548 555744 193554 555756
rect 232498 555744 232504 555756
rect 193548 555716 232504 555744
rect 193548 555704 193554 555716
rect 232498 555704 232504 555716
rect 232556 555704 232562 555756
rect 154114 555636 154120 555688
rect 154172 555676 154178 555688
rect 212902 555676 212908 555688
rect 154172 555648 212908 555676
rect 154172 555636 154178 555648
rect 212902 555636 212908 555648
rect 212960 555636 212966 555688
rect 121086 555568 121092 555620
rect 121144 555608 121150 555620
rect 197998 555608 198004 555620
rect 121144 555580 198004 555608
rect 121144 555568 121150 555580
rect 197998 555568 198004 555580
rect 198056 555568 198062 555620
rect 251542 555568 251548 555620
rect 251600 555608 251606 555620
rect 323762 555608 323768 555620
rect 251600 555580 323768 555608
rect 251600 555568 251606 555580
rect 323762 555568 323768 555580
rect 323820 555568 323826 555620
rect 71038 555500 71044 555552
rect 71096 555540 71102 555552
rect 105354 555540 105360 555552
rect 71096 555512 105360 555540
rect 71096 555500 71102 555512
rect 105354 555500 105360 555512
rect 105412 555500 105418 555552
rect 191374 555500 191380 555552
rect 191432 555540 191438 555552
rect 277394 555540 277400 555552
rect 191432 555512 277400 555540
rect 191432 555500 191438 555512
rect 277394 555500 277400 555512
rect 277452 555500 277458 555552
rect 279510 555500 279516 555552
rect 279568 555540 279574 555552
rect 313918 555540 313924 555552
rect 279568 555512 313924 555540
rect 279568 555500 279574 555512
rect 313918 555500 313924 555512
rect 313976 555500 313982 555552
rect 57606 555432 57612 555484
rect 57664 555472 57670 555484
rect 77202 555472 77208 555484
rect 57664 555444 77208 555472
rect 57664 555432 57670 555444
rect 77202 555432 77208 555444
rect 77260 555432 77266 555484
rect 82446 555432 82452 555484
rect 82504 555472 82510 555484
rect 116670 555472 116676 555484
rect 82504 555444 116676 555472
rect 82504 555432 82510 555444
rect 116670 555432 116676 555444
rect 116728 555432 116734 555484
rect 148686 555432 148692 555484
rect 148744 555472 148750 555484
rect 160554 555472 160560 555484
rect 148744 555444 160560 555472
rect 148744 555432 148750 555444
rect 160554 555432 160560 555444
rect 160612 555432 160618 555484
rect 198550 555432 198556 555484
rect 198608 555472 198614 555484
rect 287698 555472 287704 555484
rect 198608 555444 287704 555472
rect 198608 555432 198614 555444
rect 287698 555432 287704 555444
rect 287756 555432 287762 555484
rect 259454 554208 259460 554260
rect 259512 554248 259518 554260
rect 320818 554248 320824 554260
rect 259512 554220 320824 554248
rect 259512 554208 259518 554220
rect 320818 554208 320824 554220
rect 320876 554208 320882 554260
rect 184934 554140 184940 554192
rect 184992 554180 184998 554192
rect 235350 554180 235356 554192
rect 184992 554152 235356 554180
rect 184992 554140 184998 554152
rect 235350 554140 235356 554152
rect 235408 554140 235414 554192
rect 253658 554140 253664 554192
rect 253716 554180 253722 554192
rect 323670 554180 323676 554192
rect 253716 554152 323676 554180
rect 253716 554140 253722 554152
rect 323670 554140 323676 554152
rect 323728 554140 323734 554192
rect 76742 554072 76748 554124
rect 76800 554112 76806 554124
rect 116578 554112 116584 554124
rect 76800 554084 116584 554112
rect 76800 554072 76806 554084
rect 116578 554072 116584 554084
rect 116636 554072 116642 554124
rect 148410 554072 148416 554124
rect 148468 554112 148474 554124
rect 172514 554112 172520 554124
rect 148468 554084 172520 554112
rect 148468 554072 148474 554084
rect 172514 554072 172520 554084
rect 172572 554072 172578 554124
rect 192754 554072 192760 554124
rect 192812 554112 192818 554124
rect 280798 554112 280804 554124
rect 192812 554084 280804 554112
rect 192812 554072 192818 554084
rect 280798 554072 280804 554084
rect 280856 554072 280862 554124
rect 63126 554004 63132 554056
rect 63184 554044 63190 554056
rect 110598 554044 110604 554056
rect 63184 554016 110604 554044
rect 63184 554004 63190 554016
rect 110598 554004 110604 554016
rect 110656 554004 110662 554056
rect 140498 554004 140504 554056
rect 140556 554044 140562 554056
rect 193858 554044 193864 554056
rect 140556 554016 193864 554044
rect 140556 554004 140562 554016
rect 193858 554004 193864 554016
rect 193916 554004 193922 554056
rect 197078 554004 197084 554056
rect 197136 554044 197142 554056
rect 302602 554044 302608 554056
rect 197136 554016 302608 554044
rect 197136 554004 197142 554016
rect 302602 554004 302608 554016
rect 302660 554004 302666 554056
rect 290918 552916 290924 552968
rect 290976 552956 290982 552968
rect 295334 552956 295340 552968
rect 290976 552928 295340 552956
rect 290976 552916 290982 552928
rect 295334 552916 295340 552928
rect 295392 552916 295398 552968
rect 145006 552848 145012 552900
rect 145064 552888 145070 552900
rect 146202 552888 146208 552900
rect 145064 552860 146208 552888
rect 145064 552848 145070 552860
rect 146202 552848 146208 552860
rect 146260 552848 146266 552900
rect 235258 552888 235264 552900
rect 219406 552860 235264 552888
rect 107746 552780 107752 552832
rect 107804 552820 107810 552832
rect 108942 552820 108948 552832
rect 107804 552792 108948 552820
rect 107804 552780 107810 552792
rect 108942 552780 108948 552792
rect 109000 552780 109006 552832
rect 123294 552820 123300 552832
rect 122806 552792 123300 552820
rect 64966 552712 64972 552764
rect 65024 552752 65030 552764
rect 65978 552752 65984 552764
rect 65024 552724 65984 552752
rect 65024 552712 65030 552724
rect 65978 552712 65984 552724
rect 66036 552712 66042 552764
rect 67634 552712 67640 552764
rect 67692 552752 67698 552764
rect 68830 552752 68836 552764
rect 67692 552724 68836 552752
rect 67692 552712 67698 552724
rect 68830 552712 68836 552724
rect 68888 552712 68894 552764
rect 69014 552712 69020 552764
rect 69072 552752 69078 552764
rect 70302 552752 70308 552764
rect 69072 552724 70308 552752
rect 69072 552712 69078 552724
rect 70302 552712 70308 552724
rect 70360 552712 70366 552764
rect 78674 552712 78680 552764
rect 78732 552752 78738 552764
rect 79594 552752 79600 552764
rect 78732 552724 79600 552752
rect 78732 552712 78738 552724
rect 79594 552712 79600 552724
rect 79652 552712 79658 552764
rect 89714 552712 89720 552764
rect 89772 552752 89778 552764
rect 91002 552752 91008 552764
rect 89772 552724 91008 552752
rect 89772 552712 89778 552724
rect 91002 552712 91008 552724
rect 91060 552712 91066 552764
rect 94590 552712 94596 552764
rect 94648 552752 94654 552764
rect 122806 552752 122834 552792
rect 123294 552780 123300 552792
rect 123352 552780 123358 552832
rect 171318 552780 171324 552832
rect 171376 552820 171382 552832
rect 210878 552820 210884 552832
rect 171376 552792 210884 552820
rect 171376 552780 171382 552792
rect 210878 552780 210884 552792
rect 210936 552780 210942 552832
rect 211154 552780 211160 552832
rect 211212 552820 211218 552832
rect 212166 552820 212172 552832
rect 211212 552792 212172 552820
rect 211212 552780 211218 552792
rect 212166 552780 212172 552792
rect 212224 552780 212230 552832
rect 213546 552780 213552 552832
rect 213604 552820 213610 552832
rect 219406 552820 219434 552860
rect 235258 552848 235264 552860
rect 235316 552848 235322 552900
rect 283742 552848 283748 552900
rect 283800 552888 283806 552900
rect 309870 552888 309876 552900
rect 283800 552860 309876 552888
rect 283800 552848 283806 552860
rect 309870 552848 309876 552860
rect 309928 552848 309934 552900
rect 213604 552792 219434 552820
rect 213604 552780 213610 552792
rect 222194 552780 222200 552832
rect 222252 552820 222258 552832
rect 222838 552820 222844 552832
rect 222252 552792 222844 552820
rect 222252 552780 222258 552792
rect 222838 552780 222844 552792
rect 222896 552780 222902 552832
rect 227714 552780 227720 552832
rect 227772 552820 227778 552832
rect 228634 552820 228640 552832
rect 227772 552792 228640 552820
rect 227772 552780 227778 552792
rect 228634 552780 228640 552792
rect 228692 552780 228698 552832
rect 238294 552820 238300 552832
rect 230952 552792 238300 552820
rect 94648 552724 122834 552752
rect 94648 552712 94654 552724
rect 124214 552712 124220 552764
rect 124272 552752 124278 552764
rect 125410 552752 125416 552764
rect 124272 552724 125416 552752
rect 124272 552712 124278 552724
rect 125410 552712 125416 552724
rect 125468 552712 125474 552764
rect 126974 552712 126980 552764
rect 127032 552752 127038 552764
rect 128262 552752 128268 552764
rect 127032 552724 128268 552752
rect 127032 552712 127038 552724
rect 128262 552712 128268 552724
rect 128320 552712 128326 552764
rect 129734 552712 129740 552764
rect 129792 552752 129798 552764
rect 130470 552752 130476 552764
rect 129792 552724 130476 552752
rect 129792 552712 129798 552724
rect 130470 552712 130476 552724
rect 130528 552712 130534 552764
rect 136634 552712 136640 552764
rect 136692 552752 136698 552764
rect 137646 552752 137652 552764
rect 136692 552724 137652 552752
rect 136692 552712 136698 552724
rect 137646 552712 137652 552724
rect 137704 552712 137710 552764
rect 140774 552712 140780 552764
rect 140832 552752 140838 552764
rect 141878 552752 141884 552764
rect 140832 552724 141884 552752
rect 140832 552712 140838 552724
rect 141878 552712 141884 552724
rect 141936 552712 141942 552764
rect 142154 552712 142160 552764
rect 142212 552752 142218 552764
rect 143350 552752 143356 552764
rect 142212 552724 143356 552752
rect 142212 552712 142218 552724
rect 143350 552712 143356 552724
rect 143408 552712 143414 552764
rect 143534 552712 143540 552764
rect 143592 552752 143598 552764
rect 144730 552752 144736 552764
rect 143592 552724 144736 552752
rect 143592 552712 143598 552724
rect 144730 552712 144736 552724
rect 144788 552712 144794 552764
rect 147674 552712 147680 552764
rect 147732 552752 147738 552764
rect 191098 552752 191104 552764
rect 147732 552724 191104 552752
rect 147732 552712 147738 552724
rect 191098 552712 191104 552724
rect 191156 552712 191162 552764
rect 198734 552712 198740 552764
rect 198792 552752 198798 552764
rect 199930 552752 199936 552764
rect 198792 552724 199936 552752
rect 198792 552712 198798 552724
rect 199930 552712 199936 552724
rect 199988 552712 199994 552764
rect 200114 552712 200120 552764
rect 200172 552752 200178 552764
rect 201402 552752 201408 552764
rect 200172 552724 201408 552752
rect 200172 552712 200178 552724
rect 201402 552712 201408 552724
rect 201460 552712 201466 552764
rect 208578 552712 208584 552764
rect 208636 552752 208642 552764
rect 230952 552752 230980 552792
rect 238294 552780 238300 552792
rect 238352 552780 238358 552832
rect 255314 552780 255320 552832
rect 255372 552820 255378 552832
rect 256510 552820 256516 552832
rect 255372 552792 256516 552820
rect 255372 552780 255378 552792
rect 256510 552780 256516 552792
rect 256568 552780 256574 552832
rect 256786 552780 256792 552832
rect 256844 552820 256850 552832
rect 257982 552820 257988 552832
rect 256844 552792 257988 552820
rect 256844 552780 256850 552792
rect 257982 552780 257988 552792
rect 258040 552780 258046 552832
rect 267274 552780 267280 552832
rect 267332 552820 267338 552832
rect 311158 552820 311164 552832
rect 267332 552792 311164 552820
rect 267332 552780 267338 552792
rect 311158 552780 311164 552792
rect 311216 552780 311222 552832
rect 208636 552724 230980 552752
rect 208636 552712 208642 552724
rect 231854 552712 231860 552764
rect 231912 552752 231918 552764
rect 232866 552752 232872 552764
rect 231912 552724 232872 552752
rect 231912 552712 231918 552724
rect 232866 552712 232872 552724
rect 232924 552712 232930 552764
rect 233234 552712 233240 552764
rect 233292 552752 233298 552764
rect 234338 552752 234344 552764
rect 233292 552724 234344 552752
rect 233292 552712 233298 552724
rect 234338 552712 234344 552724
rect 234396 552712 234402 552764
rect 246482 552712 246488 552764
rect 246540 552752 246546 552764
rect 311250 552752 311256 552764
rect 246540 552724 311256 552752
rect 246540 552712 246546 552724
rect 311250 552712 311256 552724
rect 311308 552712 311314 552764
rect 57698 552644 57704 552696
rect 57756 552684 57762 552696
rect 103238 552684 103244 552696
rect 57756 552656 103244 552684
rect 57756 552644 57762 552656
rect 103238 552644 103244 552656
rect 103296 552644 103302 552696
rect 104894 552644 104900 552696
rect 104952 552684 104958 552696
rect 106090 552684 106096 552696
rect 104952 552656 106096 552684
rect 104952 552644 104958 552656
rect 106090 552644 106096 552656
rect 106148 552644 106154 552696
rect 106274 552644 106280 552696
rect 106332 552684 106338 552696
rect 107562 552684 107568 552696
rect 106332 552656 107568 552684
rect 106332 552644 106338 552656
rect 107562 552644 107568 552656
rect 107620 552644 107626 552696
rect 121454 552644 121460 552696
rect 121512 552684 121518 552696
rect 122558 552684 122564 552696
rect 121512 552656 122564 552684
rect 121512 552644 121518 552656
rect 122558 552644 122564 552656
rect 122616 552644 122622 552696
rect 122834 552644 122840 552696
rect 122892 552684 122898 552696
rect 124030 552684 124036 552696
rect 122892 552656 124036 552684
rect 122892 552644 122898 552656
rect 124030 552644 124036 552656
rect 124088 552644 124094 552696
rect 151170 552644 151176 552696
rect 151228 552684 151234 552696
rect 163406 552684 163412 552696
rect 151228 552656 163412 552684
rect 151228 552644 151234 552656
rect 163406 552644 163412 552656
rect 163464 552644 163470 552696
rect 168374 552644 168380 552696
rect 168432 552684 168438 552696
rect 169110 552684 169116 552696
rect 168432 552656 169116 552684
rect 168432 552644 168438 552656
rect 169110 552644 169116 552656
rect 169168 552644 169174 552696
rect 179414 552644 179420 552696
rect 179472 552684 179478 552696
rect 180610 552684 180616 552696
rect 179472 552656 180616 552684
rect 179472 552644 179478 552656
rect 180610 552644 180616 552656
rect 180668 552644 180674 552696
rect 180794 552644 180800 552696
rect 180852 552684 180858 552696
rect 181990 552684 181996 552696
rect 180852 552656 181996 552684
rect 180852 552644 180858 552656
rect 181990 552644 181996 552656
rect 182048 552644 182054 552696
rect 301222 552684 301228 552696
rect 190426 552656 301228 552684
rect 181346 552576 181352 552628
rect 181404 552616 181410 552628
rect 190426 552616 190454 552656
rect 301222 552644 301228 552656
rect 301280 552644 301286 552696
rect 181404 552588 190454 552616
rect 181404 552576 181410 552588
rect 219434 552576 219440 552628
rect 219492 552616 219498 552628
rect 220722 552616 220728 552628
rect 219492 552588 220728 552616
rect 219492 552576 219498 552588
rect 220722 552576 220728 552588
rect 220780 552576 220786 552628
rect 273254 552576 273260 552628
rect 273312 552616 273318 552628
rect 274450 552616 274456 552628
rect 273312 552588 274456 552616
rect 273312 552576 273318 552588
rect 274450 552576 274456 552588
rect 274508 552576 274514 552628
rect 291194 552576 291200 552628
rect 291252 552616 291258 552628
rect 292390 552616 292396 552628
rect 291252 552588 292396 552616
rect 291252 552576 291258 552588
rect 292390 552576 292396 552588
rect 292448 552576 292454 552628
rect 293954 552576 293960 552628
rect 294012 552616 294018 552628
rect 295242 552616 295248 552628
rect 294012 552588 295248 552616
rect 294012 552576 294018 552588
rect 295242 552576 295248 552588
rect 295300 552576 295306 552628
rect 295334 552576 295340 552628
rect 295392 552616 295398 552628
rect 322474 552616 322480 552628
rect 295392 552588 322480 552616
rect 295392 552576 295398 552588
rect 322474 552576 322480 552588
rect 322532 552576 322538 552628
rect 286686 552508 286692 552560
rect 286744 552548 286750 552560
rect 319530 552548 319536 552560
rect 286744 552520 319536 552548
rect 286744 552508 286750 552520
rect 319530 552508 319536 552520
rect 319588 552508 319594 552560
rect 285674 552440 285680 552492
rect 285732 552480 285738 552492
rect 321002 552480 321008 552492
rect 285732 552452 321008 552480
rect 285732 552440 285738 552452
rect 321002 552440 321008 552452
rect 321060 552440 321066 552492
rect 285950 552372 285956 552424
rect 286008 552412 286014 552424
rect 322658 552412 322664 552424
rect 286008 552384 322664 552412
rect 286008 552372 286014 552384
rect 322658 552372 322664 552384
rect 322716 552372 322722 552424
rect 285214 552304 285220 552356
rect 285272 552344 285278 552356
rect 322290 552344 322296 552356
rect 285272 552316 322296 552344
rect 285272 552304 285278 552316
rect 322290 552304 322296 552316
rect 322348 552304 322354 552356
rect 258718 552236 258724 552288
rect 258776 552276 258782 552288
rect 321094 552276 321100 552288
rect 258776 552248 321100 552276
rect 258776 552236 258782 552248
rect 321094 552236 321100 552248
rect 321152 552236 321158 552288
rect 252278 552168 252284 552220
rect 252336 552208 252342 552220
rect 321554 552208 321560 552220
rect 252336 552180 321560 552208
rect 252336 552168 252342 552180
rect 321554 552168 321560 552180
rect 321612 552168 321618 552220
rect 241606 552100 241612 552152
rect 241664 552140 241670 552152
rect 320910 552140 320916 552152
rect 241664 552112 320916 552140
rect 241664 552100 241670 552112
rect 320910 552100 320916 552112
rect 320968 552100 320974 552152
rect 237926 552032 237932 552084
rect 237984 552072 237990 552084
rect 320818 552072 320824 552084
rect 237984 552044 320824 552072
rect 237984 552032 237990 552044
rect 320818 552032 320824 552044
rect 320876 552032 320882 552084
rect 113266 551964 113272 552016
rect 113324 552004 113330 552016
rect 121914 552004 121920 552016
rect 113324 551976 121920 552004
rect 113324 551964 113330 551976
rect 121914 551964 121920 551976
rect 121972 551964 121978 552016
rect 148502 551964 148508 552016
rect 148560 552004 148566 552016
rect 149054 552004 149060 552016
rect 148560 551976 149060 552004
rect 148560 551964 148566 551976
rect 149054 551964 149060 551976
rect 149112 551964 149118 552016
rect 211430 551964 211436 552016
rect 211488 552004 211494 552016
rect 214650 552004 214656 552016
rect 211488 551976 214656 552004
rect 211488 551964 211494 551976
rect 214650 551964 214656 551976
rect 214708 551964 214714 552016
rect 207106 551488 207112 551540
rect 207164 551528 207170 551540
rect 229738 551528 229744 551540
rect 207164 551500 229744 551528
rect 207164 551488 207170 551500
rect 229738 551488 229744 551500
rect 229796 551488 229802 551540
rect 244366 551488 244372 551540
rect 244424 551528 244430 551540
rect 304258 551528 304264 551540
rect 244424 551500 304264 551528
rect 244424 551488 244430 551500
rect 304258 551488 304264 551500
rect 304316 551488 304322 551540
rect 189902 551420 189908 551472
rect 189960 551460 189966 551472
rect 238110 551460 238116 551472
rect 189960 551432 238116 551460
rect 189960 551420 189966 551432
rect 238110 551420 238116 551432
rect 238168 551420 238174 551472
rect 249426 551420 249432 551472
rect 249484 551460 249490 551472
rect 321186 551460 321192 551472
rect 249484 551432 321192 551460
rect 249484 551420 249490 551432
rect 321186 551420 321192 551432
rect 321244 551420 321250 551472
rect 147490 551352 147496 551404
rect 147548 551392 147554 551404
rect 166994 551392 167000 551404
rect 147548 551364 167000 551392
rect 147548 551352 147554 551364
rect 166994 551352 167000 551364
rect 167052 551352 167058 551404
rect 202782 551352 202788 551404
rect 202840 551392 202846 551404
rect 256694 551392 256700 551404
rect 202840 551364 256700 551392
rect 202840 551352 202846 551364
rect 256694 551352 256700 551364
rect 256752 551352 256758 551404
rect 86218 551284 86224 551336
rect 86276 551324 86282 551336
rect 114646 551324 114652 551336
rect 86276 551296 114652 551324
rect 86276 551284 86282 551296
rect 114646 551284 114652 551296
rect 114704 551284 114710 551336
rect 120442 551284 120448 551336
rect 120500 551324 120506 551336
rect 130378 551324 130384 551336
rect 120500 551296 130384 551324
rect 120500 551284 120506 551296
rect 130378 551284 130384 551296
rect 130436 551284 130442 551336
rect 142614 551284 142620 551336
rect 142672 551324 142678 551336
rect 211522 551324 211528 551336
rect 142672 551296 211528 551324
rect 142672 551284 142678 551296
rect 211522 551284 211528 551296
rect 211580 551284 211586 551336
rect 271598 551284 271604 551336
rect 271656 551324 271662 551336
rect 312538 551324 312544 551336
rect 271656 551296 312544 551324
rect 271656 551284 271662 551296
rect 312538 551284 312544 551296
rect 312596 551284 312602 551336
rect 262306 551216 262312 551268
rect 262364 551256 262370 551268
rect 300118 551256 300124 551268
rect 262364 551228 300124 551256
rect 262364 551216 262370 551228
rect 300118 551216 300124 551228
rect 300176 551216 300182 551268
rect 264422 551148 264428 551200
rect 264480 551188 264486 551200
rect 302878 551188 302884 551200
rect 264480 551160 302884 551188
rect 264480 551148 264486 551160
rect 302878 551148 302884 551160
rect 302936 551148 302942 551200
rect 254394 551080 254400 551132
rect 254452 551120 254458 551132
rect 302970 551120 302976 551132
rect 254452 551092 302976 551120
rect 254452 551080 254458 551092
rect 302970 551080 302976 551092
rect 303028 551080 303034 551132
rect 273714 551012 273720 551064
rect 273772 551052 273778 551064
rect 322566 551052 322572 551064
rect 273772 551024 322572 551052
rect 273772 551012 273778 551024
rect 322566 551012 322572 551024
rect 322624 551012 322630 551064
rect 272334 550944 272340 550996
rect 272392 550984 272398 550996
rect 323670 550984 323676 550996
rect 272392 550956 323676 550984
rect 272392 550944 272398 550956
rect 323670 550944 323676 550956
rect 323728 550944 323734 550996
rect 273070 550876 273076 550928
rect 273128 550916 273134 550928
rect 324774 550916 324780 550928
rect 273128 550888 324780 550916
rect 273128 550876 273134 550888
rect 324774 550876 324780 550888
rect 324832 550876 324838 550928
rect 265894 550808 265900 550860
rect 265952 550848 265958 550860
rect 324682 550848 324688 550860
rect 265952 550820 324688 550848
rect 265952 550808 265958 550820
rect 324682 550808 324688 550820
rect 324740 550808 324746 550860
rect 135438 550740 135444 550792
rect 135496 550780 135502 550792
rect 144178 550780 144184 550792
rect 135496 550752 144184 550780
rect 135496 550740 135502 550752
rect 144178 550740 144184 550752
rect 144236 550740 144242 550792
rect 287330 550740 287336 550792
rect 287388 550780 287394 550792
rect 322382 550780 322388 550792
rect 287388 550752 322388 550780
rect 287388 550740 287394 550752
rect 322382 550740 322388 550752
rect 322440 550740 322446 550792
rect 164326 550672 164332 550724
rect 164384 550712 164390 550724
rect 165522 550712 165528 550724
rect 164384 550684 165528 550712
rect 164384 550672 164390 550684
rect 165522 550672 165528 550684
rect 165580 550672 165586 550724
rect 255866 550672 255872 550724
rect 255924 550712 255930 550724
rect 324866 550712 324872 550724
rect 255924 550684 324872 550712
rect 255924 550672 255930 550684
rect 324866 550672 324872 550684
rect 324924 550672 324930 550724
rect 291654 550604 291660 550656
rect 291712 550644 291718 550656
rect 319438 550644 319444 550656
rect 291712 550616 319444 550644
rect 291712 550604 291718 550616
rect 319438 550604 319444 550616
rect 319496 550604 319502 550656
rect 61654 550536 61660 550588
rect 61712 550576 61718 550588
rect 62758 550576 62764 550588
rect 61712 550548 62764 550576
rect 61712 550536 61718 550548
rect 62758 550536 62764 550548
rect 62816 550536 62822 550588
rect 79318 550536 79324 550588
rect 79376 550576 79382 550588
rect 81710 550576 81716 550588
rect 79376 550548 81716 550576
rect 79376 550536 79382 550548
rect 81710 550536 81716 550548
rect 81768 550536 81774 550588
rect 108298 550536 108304 550588
rect 108356 550576 108362 550588
rect 111794 550576 111800 550588
rect 108356 550548 111800 550576
rect 108356 550536 108362 550548
rect 111794 550536 111800 550548
rect 111852 550536 111858 550588
rect 115474 550536 115480 550588
rect 115532 550576 115538 550588
rect 116118 550576 116124 550588
rect 115532 550548 116124 550576
rect 115532 550536 115538 550548
rect 116118 550536 116124 550548
rect 116176 550536 116182 550588
rect 136174 550536 136180 550588
rect 136232 550576 136238 550588
rect 140038 550576 140044 550588
rect 136232 550548 140044 550576
rect 136232 550536 136238 550548
rect 140038 550536 140044 550548
rect 140096 550536 140102 550588
rect 144086 550536 144092 550588
rect 144144 550576 144150 550588
rect 146846 550576 146852 550588
rect 144144 550548 146852 550576
rect 144144 550536 144150 550548
rect 146846 550536 146852 550548
rect 146904 550536 146910 550588
rect 146938 550536 146944 550588
rect 146996 550576 147002 550588
rect 148318 550576 148324 550588
rect 146996 550548 148324 550576
rect 146996 550536 147002 550548
rect 148318 550536 148324 550548
rect 148376 550536 148382 550588
rect 149882 550536 149888 550588
rect 149940 550576 149946 550588
rect 151262 550576 151268 550588
rect 149940 550548 151268 550576
rect 149940 550536 149946 550548
rect 151262 550536 151268 550548
rect 151320 550536 151326 550588
rect 219986 550536 219992 550588
rect 220044 550576 220050 550588
rect 228358 550576 228364 550588
rect 220044 550548 228364 550576
rect 220044 550536 220050 550548
rect 228358 550536 228364 550548
rect 228416 550536 228422 550588
rect 230014 550536 230020 550588
rect 230072 550576 230078 550588
rect 231118 550576 231124 550588
rect 230072 550548 231124 550576
rect 230072 550536 230078 550548
rect 231118 550536 231124 550548
rect 231176 550536 231182 550588
rect 235074 550536 235080 550588
rect 235132 550576 235138 550588
rect 236638 550576 236644 550588
rect 235132 550548 236644 550576
rect 235132 550536 235138 550548
rect 236638 550536 236644 550548
rect 236696 550536 236702 550588
rect 55122 550468 55128 550520
rect 55180 550508 55186 550520
rect 67358 550508 67364 550520
rect 55180 550480 67364 550508
rect 55180 550468 55186 550480
rect 67358 550468 67364 550480
rect 67416 550468 67422 550520
rect 209222 550468 209228 550520
rect 209280 550508 209286 550520
rect 216030 550508 216036 550520
rect 209280 550480 216036 550508
rect 209280 550468 209286 550480
rect 216030 550468 216036 550480
rect 216088 550468 216094 550520
rect 118234 550400 118240 550452
rect 118292 550440 118298 550452
rect 126238 550440 126244 550452
rect 118292 550412 126244 550440
rect 118292 550400 118298 550412
rect 126238 550400 126244 550412
rect 126296 550400 126302 550452
rect 209958 550400 209964 550452
rect 210016 550440 210022 550452
rect 220078 550440 220084 550452
rect 210016 550412 220084 550440
rect 210016 550400 210022 550412
rect 220078 550400 220084 550412
rect 220136 550400 220142 550452
rect 54938 550332 54944 550384
rect 54996 550372 55002 550384
rect 88886 550372 88892 550384
rect 54996 550344 88892 550372
rect 54996 550332 55002 550344
rect 88886 550332 88892 550344
rect 88944 550332 88950 550384
rect 118970 550332 118976 550384
rect 119028 550372 119034 550384
rect 129090 550372 129096 550384
rect 119028 550344 129096 550372
rect 119028 550332 119034 550344
rect 129090 550332 129096 550344
rect 129148 550332 129154 550384
rect 203518 550332 203524 550384
rect 203576 550372 203582 550384
rect 214558 550372 214564 550384
rect 203576 550344 214564 550372
rect 203576 550332 203582 550344
rect 214558 550332 214564 550344
rect 214616 550332 214622 550384
rect 225046 550332 225052 550384
rect 225104 550372 225110 550384
rect 235534 550372 235540 550384
rect 225104 550344 235540 550372
rect 225104 550332 225110 550344
rect 235534 550332 235540 550344
rect 235592 550332 235598 550384
rect 57790 550264 57796 550316
rect 57848 550304 57854 550316
rect 93210 550304 93216 550316
rect 57848 550276 93216 550304
rect 57848 550264 57854 550276
rect 93210 550264 93216 550276
rect 93268 550264 93274 550316
rect 114002 550264 114008 550316
rect 114060 550304 114066 550316
rect 124398 550304 124404 550316
rect 114060 550276 124404 550304
rect 114060 550264 114066 550276
rect 124398 550264 124404 550276
rect 124456 550264 124462 550316
rect 151078 550264 151084 550316
rect 151136 550304 151142 550316
rect 153378 550304 153384 550316
rect 151136 550276 153384 550304
rect 151136 550264 151142 550276
rect 153378 550264 153384 550276
rect 153436 550264 153442 550316
rect 157334 550264 157340 550316
rect 157392 550304 157398 550316
rect 167086 550304 167092 550316
rect 157392 550276 167092 550304
rect 157392 550264 157398 550276
rect 167086 550264 167092 550276
rect 167144 550264 167150 550316
rect 204254 550264 204260 550316
rect 204312 550304 204318 550316
rect 217318 550304 217324 550316
rect 204312 550276 217324 550304
rect 204312 550264 204318 550276
rect 217318 550264 217324 550276
rect 217376 550264 217382 550316
rect 230750 550264 230756 550316
rect 230808 550304 230814 550316
rect 246298 550304 246304 550316
rect 230808 550276 246304 550304
rect 230808 550264 230814 550276
rect 246298 550264 246304 550276
rect 246356 550264 246362 550316
rect 56502 550196 56508 550248
rect 56560 550236 56566 550248
rect 83918 550236 83924 550248
rect 56560 550208 83924 550236
rect 56560 550196 56566 550208
rect 83918 550196 83924 550208
rect 83976 550196 83982 550248
rect 85298 550196 85304 550248
rect 85356 550236 85362 550248
rect 120902 550236 120908 550248
rect 85356 550208 120908 550236
rect 85356 550196 85362 550208
rect 120902 550196 120908 550208
rect 120960 550196 120966 550248
rect 195606 550196 195612 550248
rect 195664 550236 195670 550248
rect 215938 550236 215944 550248
rect 195664 550208 215944 550236
rect 195664 550196 195670 550208
rect 215938 550196 215944 550208
rect 215996 550196 216002 550248
rect 225782 550196 225788 550248
rect 225840 550236 225846 550248
rect 241514 550236 241520 550248
rect 225840 550208 241520 550236
rect 225840 550196 225846 550208
rect 241514 550196 241520 550208
rect 241572 550196 241578 550248
rect 295978 550196 295984 550248
rect 296036 550236 296042 550248
rect 300670 550236 300676 550248
rect 296036 550208 300676 550236
rect 296036 550196 296042 550208
rect 300670 550196 300676 550208
rect 300728 550196 300734 550248
rect 58618 550128 58624 550180
rect 58676 550168 58682 550180
rect 95326 550168 95332 550180
rect 58676 550140 95332 550168
rect 58676 550128 58682 550140
rect 95326 550128 95332 550140
rect 95384 550128 95390 550180
rect 96062 550128 96068 550180
rect 96120 550168 96126 550180
rect 119338 550168 119344 550180
rect 96120 550140 119344 550168
rect 96120 550128 96126 550140
rect 119338 550128 119344 550140
rect 119396 550128 119402 550180
rect 147582 550128 147588 550180
rect 147640 550168 147646 550180
rect 157702 550168 157708 550180
rect 147640 550140 157708 550168
rect 147640 550128 147646 550140
rect 157702 550128 157708 550140
rect 157760 550128 157766 550180
rect 160186 550128 160192 550180
rect 160244 550168 160250 550180
rect 172698 550168 172704 550180
rect 160244 550140 172704 550168
rect 160244 550128 160250 550140
rect 172698 550128 172704 550140
rect 172756 550128 172762 550180
rect 215018 550128 215024 550180
rect 215076 550168 215082 550180
rect 236730 550168 236736 550180
rect 215076 550140 236736 550168
rect 215076 550128 215082 550140
rect 236730 550128 236736 550140
rect 236788 550128 236794 550180
rect 242250 550128 242256 550180
rect 242308 550168 242314 550180
rect 303154 550168 303160 550180
rect 242308 550140 303160 550168
rect 242308 550128 242314 550140
rect 303154 550128 303160 550140
rect 303212 550128 303218 550180
rect 55030 550060 55036 550112
rect 55088 550100 55094 550112
rect 98914 550100 98920 550112
rect 55088 550072 98920 550100
rect 55088 550060 55094 550072
rect 98914 550060 98920 550072
rect 98972 550060 98978 550112
rect 106826 550060 106832 550112
rect 106884 550100 106890 550112
rect 124306 550100 124312 550112
rect 106884 550072 124312 550100
rect 106884 550060 106890 550072
rect 124306 550060 124312 550072
rect 124364 550060 124370 550112
rect 146110 550060 146116 550112
rect 146168 550100 146174 550112
rect 156966 550100 156972 550112
rect 146168 550072 156972 550100
rect 146168 550060 146174 550072
rect 156966 550060 156972 550072
rect 157024 550060 157030 550112
rect 170582 550060 170588 550112
rect 170640 550100 170646 550112
rect 195238 550100 195244 550112
rect 170640 550072 195244 550100
rect 170640 550060 170646 550072
rect 195238 550060 195244 550072
rect 195296 550060 195302 550112
rect 212810 550060 212816 550112
rect 212868 550100 212874 550112
rect 249058 550100 249064 550112
rect 212868 550072 249064 550100
rect 212868 550060 212874 550072
rect 249058 550060 249064 550072
rect 249116 550060 249122 550112
rect 270862 550060 270868 550112
rect 270920 550100 270926 550112
rect 322750 550100 322756 550112
rect 270920 550072 322756 550100
rect 270920 550060 270926 550072
rect 322750 550060 322756 550072
rect 322808 550060 322814 550112
rect 56410 549992 56416 550044
rect 56468 550032 56474 550044
rect 73798 550032 73804 550044
rect 56468 550004 73804 550032
rect 56468 549992 56474 550004
rect 73798 549992 73804 550004
rect 73856 549992 73862 550044
rect 78122 549992 78128 550044
rect 78180 550032 78186 550044
rect 121546 550032 121552 550044
rect 78180 550004 121552 550032
rect 78180 549992 78186 550004
rect 121546 549992 121552 550004
rect 121604 549992 121610 550044
rect 151998 549992 152004 550044
rect 152056 550032 152062 550044
rect 152056 550004 161704 550032
rect 152056 549992 152062 550004
rect 56318 549924 56324 549976
rect 56376 549964 56382 549976
rect 99650 549964 99656 549976
rect 56376 549936 99656 549964
rect 56376 549924 56382 549936
rect 99650 549924 99656 549936
rect 99708 549924 99714 549976
rect 103974 549924 103980 549976
rect 104032 549964 104038 549976
rect 125778 549964 125784 549976
rect 104032 549936 125784 549964
rect 104032 549924 104038 549936
rect 125778 549924 125784 549936
rect 125836 549924 125842 549976
rect 148962 549924 148968 549976
rect 149020 549964 149026 549976
rect 161676 549964 161704 550004
rect 166994 549992 167000 550044
rect 167052 550032 167058 550044
rect 175550 550032 175556 550044
rect 167052 550004 175556 550032
rect 167052 549992 167058 550004
rect 175550 549992 175556 550004
rect 175608 549992 175614 550044
rect 183462 549992 183468 550044
rect 183520 550032 183526 550044
rect 231210 550032 231216 550044
rect 183520 550004 231216 550032
rect 183520 549992 183526 550004
rect 231210 549992 231216 550004
rect 231268 549992 231274 550044
rect 252922 549992 252928 550044
rect 252980 550032 252986 550044
rect 321278 550032 321284 550044
rect 252980 550004 321284 550032
rect 252980 549992 252986 550004
rect 321278 549992 321284 550004
rect 321336 549992 321342 550044
rect 167730 549964 167736 549976
rect 149020 549936 161520 549964
rect 161676 549936 167736 549964
rect 149020 549924 149026 549936
rect 60366 549856 60372 549908
rect 60424 549896 60430 549908
rect 116854 549896 116860 549908
rect 60424 549868 116860 549896
rect 60424 549856 60430 549868
rect 116854 549856 116860 549868
rect 116912 549856 116918 549908
rect 121822 549856 121828 549908
rect 121880 549896 121886 549908
rect 121880 549868 157334 549896
rect 121880 549856 121886 549868
rect 157306 549760 157334 549868
rect 161492 549828 161520 549936
rect 167730 549924 167736 549936
rect 167788 549924 167794 549976
rect 176286 549924 176292 549976
rect 176344 549964 176350 549976
rect 238202 549964 238208 549976
rect 176344 549936 238208 549964
rect 176344 549924 176350 549936
rect 238202 549924 238208 549936
rect 238260 549924 238266 549976
rect 299566 549924 299572 549976
rect 299624 549964 299630 549976
rect 316678 549964 316684 549976
rect 299624 549936 316684 549964
rect 299624 549924 299630 549936
rect 316678 549924 316684 549936
rect 316736 549924 316742 549976
rect 171962 549896 171968 549908
rect 164206 549868 171968 549896
rect 164206 549828 164234 549868
rect 171962 549856 171968 549868
rect 172020 549856 172026 549908
rect 192478 549896 192484 549908
rect 173866 549868 192484 549896
rect 161492 549800 164234 549828
rect 157306 549732 164234 549760
rect 164206 549692 164234 549732
rect 169754 549720 169760 549772
rect 169812 549760 169818 549772
rect 173434 549760 173440 549772
rect 169812 549732 173440 549760
rect 169812 549720 169818 549732
rect 173434 549720 173440 549732
rect 173492 549720 173498 549772
rect 173866 549692 173894 549868
rect 192478 549856 192484 549868
rect 192536 549856 192542 549908
rect 194226 549856 194232 549908
rect 194284 549896 194290 549908
rect 226978 549896 226984 549908
rect 194284 549868 226984 549896
rect 194284 549856 194290 549868
rect 226978 549856 226984 549868
rect 227036 549856 227042 549908
rect 237190 549856 237196 549908
rect 237248 549896 237254 549908
rect 285674 549896 285680 549908
rect 237248 549868 285680 549896
rect 237248 549856 237254 549868
rect 285674 549856 285680 549868
rect 285732 549856 285738 549908
rect 298830 549856 298836 549908
rect 298888 549896 298894 549908
rect 323578 549896 323584 549908
rect 298888 549868 323584 549896
rect 298888 549856 298894 549868
rect 323578 549856 323584 549868
rect 323636 549856 323642 549908
rect 283098 549788 283104 549840
rect 283156 549828 283162 549840
rect 301866 549828 301872 549840
rect 283156 549800 301872 549828
rect 283156 549788 283162 549800
rect 301866 549788 301872 549800
rect 301924 549788 301930 549840
rect 280154 549720 280160 549772
rect 280212 549760 280218 549772
rect 300302 549760 300308 549772
rect 280212 549732 300308 549760
rect 280212 549720 280218 549732
rect 300302 549720 300308 549732
rect 300360 549720 300366 549772
rect 164206 549664 173894 549692
rect 275922 549652 275928 549704
rect 275980 549692 275986 549704
rect 300210 549692 300216 549704
rect 275980 549664 300216 549692
rect 275980 549652 275986 549664
rect 300210 549652 300216 549664
rect 300268 549652 300274 549704
rect 277302 549584 277308 549636
rect 277360 549624 277366 549636
rect 305730 549624 305736 549636
rect 277360 549596 305736 549624
rect 277360 549584 277366 549596
rect 305730 549584 305736 549596
rect 305788 549584 305794 549636
rect 257246 549516 257252 549568
rect 257304 549556 257310 549568
rect 301590 549556 301596 549568
rect 257304 549528 301596 549556
rect 257304 549516 257310 549528
rect 301590 549516 301596 549528
rect 301648 549516 301654 549568
rect 240042 549448 240048 549500
rect 240100 549488 240106 549500
rect 273254 549488 273260 549500
rect 240100 549460 273260 549488
rect 240100 549448 240106 549460
rect 273254 549448 273260 549460
rect 273312 549448 273318 549500
rect 278038 549448 278044 549500
rect 278096 549488 278102 549500
rect 324130 549488 324136 549500
rect 278096 549460 324136 549488
rect 278096 549448 278102 549460
rect 324130 549448 324136 549460
rect 324188 549448 324194 549500
rect 138290 549380 138296 549432
rect 138348 549420 138354 549432
rect 142798 549420 142804 549432
rect 138348 549392 142804 549420
rect 138348 549380 138354 549392
rect 142798 549380 142804 549392
rect 142856 549380 142862 549432
rect 284478 549380 284484 549432
rect 284536 549420 284542 549432
rect 300486 549420 300492 549432
rect 284536 549392 300492 549420
rect 284536 549380 284542 549392
rect 300486 549380 300492 549392
rect 300544 549380 300550 549432
rect 296714 549312 296720 549364
rect 296772 549352 296778 549364
rect 323762 549352 323768 549364
rect 296772 549324 323768 549352
rect 296772 549312 296778 549324
rect 323762 549312 323768 549324
rect 323820 549312 323826 549364
rect 131206 549244 131212 549296
rect 131264 549284 131270 549296
rect 133138 549284 133144 549296
rect 131264 549256 133144 549284
rect 131264 549244 131270 549256
rect 133138 549244 133144 549256
rect 133196 549244 133202 549296
rect 281626 549244 281632 549296
rect 281684 549284 281690 549296
rect 300578 549284 300584 549296
rect 281684 549256 300584 549284
rect 281684 549244 281690 549256
rect 300578 549244 300584 549256
rect 300636 549244 300642 549296
rect 293770 548768 293776 548820
rect 293828 548808 293834 548820
rect 322842 548808 322848 548820
rect 293828 548780 322848 548808
rect 293828 548768 293834 548780
rect 322842 548768 322848 548780
rect 322900 548768 322906 548820
rect 268746 548700 268752 548752
rect 268804 548740 268810 548752
rect 303062 548740 303068 548752
rect 268804 548712 303068 548740
rect 268804 548700 268810 548712
rect 303062 548700 303068 548712
rect 303120 548700 303126 548752
rect 265158 548632 265164 548684
rect 265216 548672 265222 548684
rect 307018 548672 307024 548684
rect 265216 548644 307024 548672
rect 265216 548632 265222 548644
rect 307018 548632 307024 548644
rect 307076 548632 307082 548684
rect 278774 548564 278780 548616
rect 278832 548604 278838 548616
rect 321554 548604 321560 548616
rect 278832 548576 321560 548604
rect 278832 548564 278838 548576
rect 321554 548564 321560 548576
rect 321612 548564 321618 548616
rect 273254 548496 273260 548548
rect 273312 548536 273318 548548
rect 322106 548536 322112 548548
rect 273312 548508 322112 548536
rect 273312 548496 273318 548508
rect 322106 548496 322112 548508
rect 322164 548496 322170 548548
rect 276566 548428 276572 548480
rect 276624 548468 276630 548480
rect 324590 548468 324596 548480
rect 276624 548440 324596 548468
rect 276624 548428 276630 548440
rect 324590 548428 324596 548440
rect 324648 548428 324654 548480
rect 247218 548360 247224 548412
rect 247276 548400 247282 548412
rect 301774 548400 301780 548412
rect 247276 548372 301780 548400
rect 247276 548360 247282 548372
rect 301774 548360 301780 548372
rect 301832 548360 301838 548412
rect 243630 548292 243636 548344
rect 243688 548332 243694 548344
rect 301958 548332 301964 548344
rect 243688 548304 301964 548332
rect 243688 548292 243694 548304
rect 301958 548292 301964 548304
rect 302016 548292 302022 548344
rect 263042 548224 263048 548276
rect 263100 548264 263106 548276
rect 324498 548264 324504 548276
rect 263100 548236 324504 548264
rect 263100 548224 263106 548236
rect 324498 548224 324504 548236
rect 324556 548224 324562 548276
rect 260834 548156 260840 548208
rect 260892 548196 260898 548208
rect 323854 548196 323860 548208
rect 260892 548168 323860 548196
rect 260892 548156 260898 548168
rect 323854 548156 323860 548168
rect 323912 548156 323918 548208
rect 235810 548088 235816 548140
rect 235868 548088 235874 548140
rect 236454 548088 236460 548140
rect 236512 548128 236518 548140
rect 301038 548128 301044 548140
rect 236512 548100 301044 548128
rect 236512 548088 236518 548100
rect 301038 548088 301044 548100
rect 301096 548088 301102 548140
rect 235828 548060 235856 548088
rect 323578 548060 323584 548072
rect 235828 548032 323584 548060
rect 323578 548020 323584 548032
rect 323636 548020 323642 548072
rect 301038 543668 301044 543720
rect 301096 543708 301102 543720
rect 321554 543708 321560 543720
rect 301096 543680 321560 543708
rect 301096 543668 301102 543680
rect 321554 543668 321560 543680
rect 321612 543668 321618 543720
rect 302786 539588 302792 539640
rect 302844 539628 302850 539640
rect 311158 539628 311164 539640
rect 302844 539600 311164 539628
rect 302844 539588 302850 539600
rect 311158 539588 311164 539600
rect 311216 539588 311222 539640
rect 301958 539520 301964 539572
rect 302016 539560 302022 539572
rect 321554 539560 321560 539572
rect 302016 539532 321560 539560
rect 302016 539520 302022 539532
rect 321554 539520 321560 539532
rect 321612 539520 321618 539572
rect 324682 533400 324688 533452
rect 324740 533440 324746 533452
rect 324740 533412 324820 533440
rect 324740 533400 324746 533412
rect 324792 533248 324820 533412
rect 324774 533196 324780 533248
rect 324832 533196 324838 533248
rect 300670 529864 300676 529916
rect 300728 529904 300734 529916
rect 457438 529904 457444 529916
rect 300728 529876 457444 529904
rect 300728 529864 300734 529876
rect 457438 529864 457444 529876
rect 457496 529864 457502 529916
rect 300578 529796 300584 529848
rect 300636 529836 300642 529848
rect 436462 529836 436468 529848
rect 300636 529808 436468 529836
rect 300636 529796 300642 529808
rect 436462 529796 436468 529808
rect 436520 529796 436526 529848
rect 300486 529728 300492 529780
rect 300544 529768 300550 529780
rect 436186 529768 436192 529780
rect 300544 529740 436192 529768
rect 300544 529728 300550 529740
rect 436186 529728 436192 529740
rect 436244 529728 436250 529780
rect 301866 529660 301872 529712
rect 301924 529700 301930 529712
rect 436094 529700 436100 529712
rect 301924 529672 436100 529700
rect 301924 529660 301930 529672
rect 436094 529660 436100 529672
rect 436152 529660 436158 529712
rect 303154 529592 303160 529644
rect 303212 529632 303218 529644
rect 436554 529632 436560 529644
rect 303212 529604 436560 529632
rect 303212 529592 303218 529604
rect 436554 529592 436560 529604
rect 436612 529592 436618 529644
rect 305730 529524 305736 529576
rect 305788 529564 305794 529576
rect 436370 529564 436376 529576
rect 305788 529536 436376 529564
rect 305788 529524 305794 529536
rect 436370 529524 436376 529536
rect 436428 529524 436434 529576
rect 322750 529456 322756 529508
rect 322808 529496 322814 529508
rect 436278 529496 436284 529508
rect 322808 529468 436284 529496
rect 322808 529456 322814 529468
rect 436278 529456 436284 529468
rect 436336 529456 436342 529508
rect 319530 528504 319536 528556
rect 319588 528544 319594 528556
rect 512178 528544 512184 528556
rect 319588 528516 512184 528544
rect 319588 528504 319594 528516
rect 512178 528504 512184 528516
rect 512236 528504 512242 528556
rect 322658 528436 322664 528488
rect 322716 528476 322722 528488
rect 495434 528476 495440 528488
rect 322716 528448 495440 528476
rect 322716 528436 322722 528448
rect 495434 528436 495440 528448
rect 495492 528436 495498 528488
rect 322474 528368 322480 528420
rect 322532 528408 322538 528420
rect 488534 528408 488540 528420
rect 322532 528380 488540 528408
rect 322532 528368 322538 528380
rect 488534 528368 488540 528380
rect 488592 528368 488598 528420
rect 322842 528300 322848 528352
rect 322900 528340 322906 528352
rect 465074 528340 465080 528352
rect 322900 528312 465080 528340
rect 322900 528300 322906 528312
rect 465074 528300 465080 528312
rect 465132 528300 465138 528352
rect 323762 528232 323768 528284
rect 323820 528272 323826 528284
rect 459554 528272 459560 528284
rect 323820 528244 459560 528272
rect 323820 528232 323826 528244
rect 459554 528232 459560 528244
rect 459612 528232 459618 528284
rect 300302 528164 300308 528216
rect 300360 528204 300366 528216
rect 436922 528204 436928 528216
rect 300360 528176 436928 528204
rect 300360 528164 300366 528176
rect 436922 528164 436928 528176
rect 436980 528164 436986 528216
rect 301590 528096 301596 528148
rect 301648 528136 301654 528148
rect 436830 528136 436836 528148
rect 301648 528108 436836 528136
rect 301648 528096 301654 528108
rect 436830 528096 436836 528108
rect 436888 528096 436894 528148
rect 321278 528028 321284 528080
rect 321336 528068 321342 528080
rect 436646 528068 436652 528080
rect 321336 528040 436652 528068
rect 321336 528028 321342 528040
rect 436646 528028 436652 528040
rect 436704 528028 436710 528080
rect 324130 527960 324136 528012
rect 324188 528000 324194 528012
rect 436738 528000 436744 528012
rect 324188 527972 436744 528000
rect 324188 527960 324194 527972
rect 436738 527960 436744 527972
rect 436796 527960 436802 528012
rect 305638 527892 305644 527944
rect 305696 527932 305702 527944
rect 374270 527932 374276 527944
rect 305696 527904 374276 527932
rect 305696 527892 305702 527904
rect 374270 527892 374276 527904
rect 374328 527892 374334 527944
rect 300210 527824 300216 527876
rect 300268 527864 300274 527876
rect 356238 527864 356244 527876
rect 300268 527836 356244 527864
rect 300268 527824 300274 527836
rect 356238 527824 356244 527836
rect 356296 527824 356302 527876
rect 324958 527184 324964 527196
rect 324516 527156 324964 527184
rect 307018 527076 307024 527128
rect 307076 527116 307082 527128
rect 324516 527116 324544 527156
rect 324958 527144 324964 527156
rect 325016 527144 325022 527196
rect 307076 527088 324544 527116
rect 307076 527076 307082 527088
rect 324590 527076 324596 527128
rect 324648 527116 324654 527128
rect 419994 527116 420000 527128
rect 324648 527088 420000 527116
rect 324648 527076 324654 527088
rect 419994 527076 420000 527088
rect 420052 527076 420058 527128
rect 323854 527008 323860 527060
rect 323912 527048 323918 527060
rect 347222 527048 347228 527060
rect 323912 527020 347228 527048
rect 323912 527008 323918 527020
rect 347222 527008 347228 527020
rect 347280 527008 347286 527060
rect 323578 526940 323584 526992
rect 323636 526980 323642 526992
rect 338206 526980 338212 526992
rect 323636 526952 338212 526980
rect 323636 526940 323642 526952
rect 338206 526940 338212 526952
rect 338264 526940 338270 526992
rect 324866 526872 324872 526924
rect 324924 526912 324930 526924
rect 411254 526912 411260 526924
rect 324924 526884 411260 526912
rect 324924 526872 324930 526884
rect 411254 526872 411260 526884
rect 411312 526872 411318 526924
rect 324498 526804 324504 526856
rect 324556 526844 324562 526856
rect 406470 526844 406476 526856
rect 324556 526816 406476 526844
rect 324556 526804 324562 526816
rect 406470 526804 406476 526816
rect 406528 526804 406534 526856
rect 322566 526736 322572 526788
rect 322624 526776 322630 526788
rect 401962 526776 401968 526788
rect 322624 526748 401968 526776
rect 322624 526736 322630 526748
rect 401962 526736 401968 526748
rect 402020 526736 402026 526788
rect 302878 526668 302884 526720
rect 302936 526708 302942 526720
rect 379514 526708 379520 526720
rect 302936 526680 379520 526708
rect 302936 526668 302942 526680
rect 379514 526668 379520 526680
rect 379572 526668 379578 526720
rect 324774 526600 324780 526652
rect 324832 526640 324838 526652
rect 388438 526640 388444 526652
rect 324832 526612 388444 526640
rect 324832 526600 324838 526612
rect 388438 526600 388444 526612
rect 388496 526600 388502 526652
rect 301774 526532 301780 526584
rect 301832 526572 301838 526584
rect 365254 526572 365260 526584
rect 301832 526544 365260 526572
rect 301832 526532 301838 526544
rect 365254 526532 365260 526544
rect 365312 526532 365318 526584
rect 302970 526464 302976 526516
rect 303028 526504 303034 526516
rect 351914 526504 351920 526516
rect 303028 526476 351920 526504
rect 303028 526464 303034 526476
rect 351914 526464 351920 526476
rect 351972 526464 351978 526516
rect 324682 526396 324688 526448
rect 324740 526436 324746 526448
rect 369854 526436 369860 526448
rect 324740 526408 369860 526436
rect 324740 526396 324746 526408
rect 369854 526396 369860 526408
rect 369912 526396 369918 526448
rect 323670 526328 323676 526380
rect 323728 526368 323734 526380
rect 415578 526368 415584 526380
rect 323728 526340 415584 526368
rect 323728 526328 323734 526340
rect 415578 526328 415584 526340
rect 415636 526328 415642 526380
rect 303062 526260 303068 526312
rect 303120 526300 303126 526312
rect 393314 526300 393320 526312
rect 303120 526272 393320 526300
rect 303120 526260 303126 526272
rect 393314 526260 393320 526272
rect 393372 526260 393378 526312
rect 300118 526192 300124 526244
rect 300176 526232 300182 526244
rect 333974 526232 333980 526244
rect 300176 526204 333980 526232
rect 300176 526192 300182 526204
rect 333974 526192 333980 526204
rect 334032 526192 334038 526244
rect 301498 525716 301504 525768
rect 301556 525756 301562 525768
rect 512270 525756 512276 525768
rect 301556 525728 512276 525756
rect 301556 525716 301562 525728
rect 512270 525716 512276 525728
rect 512328 525716 512334 525768
rect 322382 525648 322388 525700
rect 322440 525688 322446 525700
rect 476114 525688 476120 525700
rect 322440 525660 476120 525688
rect 322440 525648 322446 525660
rect 476114 525648 476120 525660
rect 476172 525648 476178 525700
rect 322290 525580 322296 525632
rect 322348 525620 322354 525632
rect 470594 525620 470600 525632
rect 322348 525592 470600 525620
rect 322348 525580 322354 525592
rect 470594 525580 470600 525592
rect 470652 525580 470658 525632
rect 321094 525512 321100 525564
rect 321152 525552 321158 525564
rect 433334 525552 433340 525564
rect 321152 525524 433340 525552
rect 321152 525512 321158 525524
rect 433334 525512 433340 525524
rect 433392 525512 433398 525564
rect 302878 524424 302884 524476
rect 302936 524464 302942 524476
rect 519538 524464 519544 524476
rect 302936 524436 519544 524464
rect 302936 524424 302942 524436
rect 519538 524424 519544 524436
rect 519596 524424 519602 524476
rect 319438 524356 319444 524408
rect 319496 524396 319502 524408
rect 457622 524396 457628 524408
rect 319496 524368 457628 524396
rect 319496 524356 319502 524368
rect 457622 524356 457628 524368
rect 457680 524356 457686 524408
rect 321002 524288 321008 524340
rect 321060 524328 321066 524340
rect 434622 524328 434628 524340
rect 321060 524300 434628 524328
rect 321060 524288 321066 524300
rect 434622 524288 434628 524300
rect 434680 524288 434686 524340
rect 320818 524220 320824 524272
rect 320876 524260 320882 524272
rect 433518 524260 433524 524272
rect 320876 524232 433524 524260
rect 320876 524220 320882 524232
rect 433518 524220 433524 524232
rect 433576 524220 433582 524272
rect 320910 524152 320916 524204
rect 320968 524192 320974 524204
rect 433426 524192 433432 524204
rect 320968 524164 433432 524192
rect 320968 524152 320974 524164
rect 433426 524152 433432 524164
rect 433484 524152 433490 524204
rect 329742 524084 329748 524136
rect 329800 524124 329806 524136
rect 434714 524124 434720 524136
rect 329800 524096 434720 524124
rect 329800 524084 329806 524096
rect 434714 524084 434720 524096
rect 434772 524084 434778 524136
rect 53742 517488 53748 517540
rect 53800 517528 53806 517540
rect 57882 517528 57888 517540
rect 53800 517500 57888 517528
rect 53800 517488 53806 517500
rect 57882 517488 57888 517500
rect 57940 517488 57946 517540
rect 311158 515380 311164 515432
rect 311216 515420 311222 515432
rect 580258 515420 580264 515432
rect 311216 515392 580264 515420
rect 311216 515380 311222 515392
rect 580258 515380 580264 515392
rect 580316 515380 580322 515432
rect 560938 511912 560944 511964
rect 560996 511952 561002 511964
rect 580166 511952 580172 511964
rect 560996 511924 580172 511952
rect 560996 511912 561002 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 302234 495456 302240 495508
rect 302292 495496 302298 495508
rect 520918 495496 520924 495508
rect 302292 495468 520924 495496
rect 302292 495456 302298 495468
rect 520918 495456 520924 495468
rect 520976 495456 520982 495508
rect 274650 487772 274656 487824
rect 274708 487812 274714 487824
rect 274818 487812 274824 487824
rect 274708 487784 274824 487812
rect 274708 487772 274714 487784
rect 274818 487772 274824 487784
rect 274876 487772 274882 487824
rect 64874 487024 64880 487076
rect 64932 487064 64938 487076
rect 65150 487064 65156 487076
rect 64932 487036 65156 487064
rect 64932 487024 64938 487036
rect 65150 487024 65156 487036
rect 65208 487024 65214 487076
rect 128354 487024 128360 487076
rect 128412 487064 128418 487076
rect 128630 487064 128636 487076
rect 128412 487036 128636 487064
rect 128412 487024 128418 487036
rect 128630 487024 128636 487036
rect 128688 487024 128694 487076
rect 207106 487024 207112 487076
rect 207164 487064 207170 487076
rect 207382 487064 207388 487076
rect 207164 487036 207388 487064
rect 207164 487024 207170 487036
rect 207382 487024 207388 487036
rect 207440 487024 207446 487076
rect 140866 486684 140872 486736
rect 140924 486724 140930 486736
rect 199102 486724 199108 486736
rect 140924 486696 199108 486724
rect 140924 486684 140930 486696
rect 199102 486684 199108 486696
rect 199160 486684 199166 486736
rect 121178 486616 121184 486668
rect 121236 486656 121242 486668
rect 197906 486656 197912 486668
rect 121236 486628 197912 486656
rect 121236 486616 121242 486628
rect 197906 486616 197912 486628
rect 197964 486616 197970 486668
rect 109402 486548 109408 486600
rect 109460 486588 109466 486600
rect 198366 486588 198372 486600
rect 109460 486560 198372 486588
rect 109460 486548 109466 486560
rect 198366 486548 198372 486560
rect 198424 486548 198430 486600
rect 109494 486480 109500 486532
rect 109552 486520 109558 486532
rect 204806 486520 204812 486532
rect 109552 486492 204812 486520
rect 109552 486480 109558 486492
rect 204806 486480 204812 486492
rect 204864 486480 204870 486532
rect 15838 486412 15844 486464
rect 15896 486452 15902 486464
rect 383654 486452 383660 486464
rect 15896 486424 383660 486452
rect 15896 486412 15902 486424
rect 383654 486412 383660 486424
rect 383712 486412 383718 486464
rect 73982 485732 73988 485784
rect 74040 485772 74046 485784
rect 105078 485772 105084 485784
rect 74040 485744 105084 485772
rect 74040 485732 74046 485744
rect 105078 485732 105084 485744
rect 105136 485732 105142 485784
rect 107838 485732 107844 485784
rect 107896 485772 107902 485784
rect 108022 485772 108028 485784
rect 107896 485744 108028 485772
rect 107896 485732 107902 485744
rect 108022 485732 108028 485744
rect 108080 485732 108086 485784
rect 151262 485732 151268 485784
rect 151320 485772 151326 485784
rect 204898 485772 204904 485784
rect 151320 485744 204904 485772
rect 151320 485732 151326 485744
rect 204898 485732 204904 485744
rect 204956 485732 204962 485784
rect 212074 485772 212080 485784
rect 209746 485744 212080 485772
rect 59998 485664 60004 485716
rect 60056 485704 60062 485716
rect 91830 485704 91836 485716
rect 60056 485676 91836 485704
rect 60056 485664 60062 485676
rect 91830 485664 91836 485676
rect 91888 485664 91894 485716
rect 149514 485664 149520 485716
rect 149572 485704 149578 485716
rect 201310 485704 201316 485716
rect 149572 485676 201316 485704
rect 149572 485664 149578 485676
rect 201310 485664 201316 485676
rect 201368 485664 201374 485716
rect 201402 485664 201408 485716
rect 201460 485704 201466 485716
rect 209746 485704 209774 485744
rect 212074 485732 212080 485744
rect 212132 485732 212138 485784
rect 262398 485732 262404 485784
rect 262456 485772 262462 485784
rect 262582 485772 262588 485784
rect 262456 485744 262588 485772
rect 262456 485732 262462 485744
rect 262582 485732 262588 485744
rect 262640 485732 262646 485784
rect 285766 485732 285772 485784
rect 285824 485772 285830 485784
rect 285950 485772 285956 485784
rect 285824 485744 285956 485772
rect 285824 485732 285830 485744
rect 285950 485732 285956 485744
rect 286008 485732 286014 485784
rect 201460 485676 209774 485704
rect 201460 485664 201466 485676
rect 234522 485664 234528 485716
rect 234580 485704 234586 485716
rect 234580 485676 238754 485704
rect 234580 485664 234586 485676
rect 56502 485596 56508 485648
rect 56560 485636 56566 485648
rect 89622 485636 89628 485648
rect 56560 485608 89628 485636
rect 56560 485596 56566 485608
rect 89622 485596 89628 485608
rect 89680 485596 89686 485648
rect 154298 485596 154304 485648
rect 154356 485636 154362 485648
rect 212534 485636 212540 485648
rect 154356 485608 212540 485636
rect 154356 485596 154362 485608
rect 212534 485596 212540 485608
rect 212592 485596 212598 485648
rect 59078 485528 59084 485580
rect 59136 485568 59142 485580
rect 92290 485568 92296 485580
rect 59136 485540 92296 485568
rect 59136 485528 59142 485540
rect 92290 485528 92296 485540
rect 92348 485528 92354 485580
rect 162118 485528 162124 485580
rect 162176 485568 162182 485580
rect 238726 485568 238754 485676
rect 244550 485664 244556 485716
rect 244608 485704 244614 485716
rect 356790 485704 356796 485716
rect 244608 485676 356796 485704
rect 244608 485664 244614 485676
rect 356790 485664 356796 485676
rect 356848 485664 356854 485716
rect 239674 485596 239680 485648
rect 239732 485636 239738 485648
rect 358262 485636 358268 485648
rect 239732 485608 358268 485636
rect 239732 485596 239738 485608
rect 358262 485596 358268 485608
rect 358320 485596 358326 485648
rect 364978 485568 364984 485580
rect 162176 485540 209774 485568
rect 238726 485540 364984 485568
rect 162176 485528 162182 485540
rect 64138 485460 64144 485512
rect 64196 485500 64202 485512
rect 72418 485500 72424 485512
rect 64196 485472 72424 485500
rect 64196 485460 64202 485472
rect 72418 485460 72424 485472
rect 72476 485460 72482 485512
rect 79318 485460 79324 485512
rect 79376 485500 79382 485512
rect 106366 485500 106372 485512
rect 79376 485472 106372 485500
rect 79376 485460 79382 485472
rect 106366 485460 106372 485472
rect 106424 485460 106430 485512
rect 152182 485460 152188 485512
rect 152240 485500 152246 485512
rect 204254 485500 204260 485512
rect 152240 485472 204260 485500
rect 152240 485460 152246 485472
rect 204254 485460 204260 485472
rect 204312 485460 204318 485512
rect 55122 485392 55128 485444
rect 55180 485432 55186 485444
rect 88334 485432 88340 485444
rect 55180 485404 88340 485432
rect 55180 485392 55186 485404
rect 88334 485392 88340 485404
rect 88392 485392 88398 485444
rect 149422 485392 149428 485444
rect 149480 485432 149486 485444
rect 200482 485432 200488 485444
rect 149480 485404 200488 485432
rect 149480 485392 149486 485404
rect 200482 485392 200488 485404
rect 200540 485392 200546 485444
rect 201310 485392 201316 485444
rect 201368 485432 201374 485444
rect 208486 485432 208492 485444
rect 201368 485404 208492 485432
rect 201368 485392 201374 485404
rect 208486 485392 208492 485404
rect 208544 485392 208550 485444
rect 209746 485432 209774 485540
rect 364978 485528 364984 485540
rect 365036 485528 365042 485580
rect 211062 485460 211068 485512
rect 211120 485500 211126 485512
rect 217410 485500 217416 485512
rect 211120 485472 217416 485500
rect 211120 485460 211126 485472
rect 217410 485460 217416 485472
rect 217468 485460 217474 485512
rect 226058 485460 226064 485512
rect 226116 485500 226122 485512
rect 356698 485500 356704 485512
rect 226116 485472 356704 485500
rect 226116 485460 226122 485472
rect 356698 485460 356704 485472
rect 356756 485460 356762 485512
rect 211154 485432 211160 485444
rect 209746 485404 211160 485432
rect 211154 485392 211160 485404
rect 211212 485392 211218 485444
rect 230842 485392 230848 485444
rect 230900 485432 230906 485444
rect 362218 485432 362224 485444
rect 230900 485404 362224 485432
rect 230900 485392 230906 485404
rect 362218 485392 362224 485404
rect 362276 485392 362282 485444
rect 56410 485324 56416 485376
rect 56468 485364 56474 485376
rect 90542 485364 90548 485376
rect 56468 485336 90548 485364
rect 56468 485324 56474 485336
rect 90542 485324 90548 485336
rect 90600 485324 90606 485376
rect 148226 485324 148232 485376
rect 148284 485364 148290 485376
rect 197446 485364 197452 485376
rect 148284 485336 197452 485364
rect 148284 485324 148290 485336
rect 197446 485324 197452 485336
rect 197504 485324 197510 485376
rect 209682 485324 209688 485376
rect 209740 485364 209746 485376
rect 221734 485364 221740 485376
rect 209740 485336 221740 485364
rect 209740 485324 209746 485336
rect 221734 485324 221740 485336
rect 221792 485324 221798 485376
rect 225598 485324 225604 485376
rect 225656 485364 225662 485376
rect 358170 485364 358176 485376
rect 225656 485336 358176 485364
rect 225656 485324 225662 485336
rect 358170 485324 358176 485336
rect 358228 485324 358234 485376
rect 50982 485256 50988 485308
rect 51040 485296 51046 485308
rect 93578 485296 93584 485308
rect 51040 485268 93584 485296
rect 51040 485256 51046 485268
rect 93578 485256 93584 485268
rect 93636 485256 93642 485308
rect 156690 485256 156696 485308
rect 156748 485296 156754 485308
rect 162118 485296 162124 485308
rect 156748 485268 162124 485296
rect 156748 485256 156754 485268
rect 162118 485256 162124 485268
rect 162176 485256 162182 485308
rect 162210 485256 162216 485308
rect 162268 485296 162274 485308
rect 205634 485296 205640 485308
rect 162268 485268 205640 485296
rect 162268 485256 162274 485268
rect 205634 485256 205640 485268
rect 205692 485256 205698 485308
rect 240042 485256 240048 485308
rect 240100 485296 240106 485308
rect 373258 485296 373264 485308
rect 240100 485268 373264 485296
rect 240100 485256 240106 485268
rect 373258 485256 373264 485268
rect 373316 485256 373322 485308
rect 51810 485188 51816 485240
rect 51868 485228 51874 485240
rect 99374 485228 99380 485240
rect 51868 485200 99380 485228
rect 51868 485188 51874 485200
rect 99374 485188 99380 485200
rect 99432 485188 99438 485240
rect 150434 485188 150440 485240
rect 150492 485228 150498 485240
rect 201494 485228 201500 485240
rect 150492 485200 190516 485228
rect 150492 485188 150498 485200
rect 42426 485120 42432 485172
rect 42484 485160 42490 485172
rect 102870 485160 102876 485172
rect 42484 485132 102876 485160
rect 42484 485120 42490 485132
rect 102870 485120 102876 485132
rect 102928 485120 102934 485172
rect 161474 485120 161480 485172
rect 161532 485160 161538 485172
rect 190488 485160 190516 485200
rect 197464 485200 201500 485228
rect 197354 485160 197360 485172
rect 161532 485132 176654 485160
rect 190488 485132 197360 485160
rect 161532 485120 161538 485132
rect 43622 485052 43628 485104
rect 43680 485092 43686 485104
rect 104618 485092 104624 485104
rect 43680 485064 104624 485092
rect 43680 485052 43686 485064
rect 104618 485052 104624 485064
rect 104676 485052 104682 485104
rect 110322 485052 110328 485104
rect 110380 485092 110386 485104
rect 170398 485092 170404 485104
rect 110380 485064 170404 485092
rect 110380 485052 110386 485064
rect 170398 485052 170404 485064
rect 170456 485052 170462 485104
rect 176626 485092 176654 485132
rect 197354 485120 197360 485132
rect 197412 485120 197418 485172
rect 197464 485092 197492 485200
rect 201494 485188 201500 485200
rect 201552 485188 201558 485240
rect 209774 485228 209780 485240
rect 204732 485200 209780 485228
rect 199378 485120 199384 485172
rect 199436 485160 199442 485172
rect 204732 485160 204760 485200
rect 209774 485188 209780 485200
rect 209832 485188 209838 485240
rect 209866 485188 209872 485240
rect 209924 485228 209930 485240
rect 219894 485228 219900 485240
rect 209924 485200 219900 485228
rect 209924 485188 209930 485200
rect 219894 485188 219900 485200
rect 219952 485188 219958 485240
rect 224034 485188 224040 485240
rect 224092 485228 224098 485240
rect 360838 485228 360844 485240
rect 224092 485200 360844 485228
rect 224092 485188 224098 485200
rect 360838 485188 360844 485200
rect 360896 485188 360902 485240
rect 199436 485132 204760 485160
rect 199436 485120 199442 485132
rect 206830 485120 206836 485172
rect 206888 485160 206894 485172
rect 219158 485160 219164 485172
rect 206888 485132 219164 485160
rect 206888 485120 206894 485132
rect 219158 485120 219164 485132
rect 219216 485120 219222 485172
rect 231762 485120 231768 485172
rect 231820 485160 231826 485172
rect 369118 485160 369124 485172
rect 231820 485132 369124 485160
rect 231820 485120 231826 485132
rect 369118 485120 369124 485132
rect 369176 485120 369182 485172
rect 176626 485064 197492 485092
rect 200206 485052 200212 485104
rect 200264 485092 200270 485104
rect 217410 485092 217416 485104
rect 200264 485064 217416 485092
rect 200264 485052 200270 485064
rect 217410 485052 217416 485064
rect 217468 485052 217474 485104
rect 223482 485052 223488 485104
rect 223540 485092 223546 485104
rect 371878 485092 371884 485104
rect 223540 485064 371884 485092
rect 223540 485052 223546 485064
rect 371878 485052 371884 485064
rect 371936 485052 371942 485104
rect 52178 484984 52184 485036
rect 52236 485024 52242 485036
rect 81710 485024 81716 485036
rect 52236 484996 81716 485024
rect 52236 484984 52242 484996
rect 81710 484984 81716 484996
rect 81768 484984 81774 485036
rect 157426 484984 157432 485036
rect 157484 485024 157490 485036
rect 162210 485024 162216 485036
rect 157484 484996 162216 485024
rect 157484 484984 157490 484996
rect 162210 484984 162216 484996
rect 162268 484984 162274 485036
rect 204254 485024 204260 485036
rect 164206 484996 204260 485024
rect 50614 484916 50620 484968
rect 50672 484956 50678 484968
rect 73246 484956 73252 484968
rect 50672 484928 73252 484956
rect 50672 484916 50678 484928
rect 73246 484916 73252 484928
rect 73304 484916 73310 484968
rect 73798 484916 73804 484968
rect 73856 484956 73862 484968
rect 79318 484956 79324 484968
rect 73856 484928 79324 484956
rect 73856 484916 73862 484928
rect 79318 484916 79324 484928
rect 79376 484916 79382 484968
rect 139394 484916 139400 484968
rect 139452 484956 139458 484968
rect 139452 484928 154574 484956
rect 139452 484916 139458 484928
rect 73890 484848 73896 484900
rect 73948 484888 73954 484900
rect 95326 484888 95332 484900
rect 73948 484860 95332 484888
rect 73948 484848 73954 484860
rect 95326 484848 95332 484860
rect 95384 484848 95390 484900
rect 50890 484780 50896 484832
rect 50948 484820 50954 484832
rect 73338 484820 73344 484832
rect 50948 484792 73344 484820
rect 50948 484780 50954 484792
rect 73338 484780 73344 484792
rect 73396 484780 73402 484832
rect 68278 484712 68284 484764
rect 68336 484752 68342 484764
rect 84378 484752 84384 484764
rect 68336 484724 84384 484752
rect 68336 484712 68342 484724
rect 84378 484712 84384 484724
rect 84436 484712 84442 484764
rect 154546 484752 154574 484928
rect 158714 484916 158720 484968
rect 158772 484956 158778 484968
rect 164206 484956 164234 484996
rect 204254 484984 204260 484996
rect 204312 484984 204318 485036
rect 209774 484984 209780 485036
rect 209832 485024 209838 485036
rect 214742 485024 214748 485036
rect 209832 484996 214748 485024
rect 209832 484984 209838 484996
rect 214742 484984 214748 484996
rect 214800 484984 214806 485036
rect 185578 484956 185584 484968
rect 158772 484928 164234 484956
rect 166966 484928 185584 484956
rect 158772 484916 158778 484928
rect 155586 484848 155592 484900
rect 155644 484888 155650 484900
rect 161474 484888 161480 484900
rect 155644 484860 161480 484888
rect 155644 484848 155650 484860
rect 161474 484848 161480 484860
rect 161532 484848 161538 484900
rect 166966 484888 166994 484928
rect 185578 484916 185584 484928
rect 185636 484916 185642 484968
rect 195330 484916 195336 484968
rect 195388 484956 195394 484968
rect 211614 484956 211620 484968
rect 195388 484928 211620 484956
rect 195388 484916 195394 484928
rect 211614 484916 211620 484928
rect 211672 484916 211678 484968
rect 203518 484888 203524 484900
rect 164206 484860 166994 484888
rect 171106 484860 203524 484888
rect 164206 484752 164234 484860
rect 166258 484780 166264 484832
rect 166316 484820 166322 484832
rect 171106 484820 171134 484860
rect 203518 484848 203524 484860
rect 203576 484848 203582 484900
rect 166316 484792 171134 484820
rect 166316 484780 166322 484792
rect 204898 484780 204904 484832
rect 204956 484820 204962 484832
rect 211154 484820 211160 484832
rect 204956 484792 211160 484820
rect 204956 484780 204962 484792
rect 211154 484780 211160 484792
rect 211212 484780 211218 484832
rect 154546 484724 164234 484752
rect 212534 484440 212540 484492
rect 212592 484480 212598 484492
rect 212718 484480 212724 484492
rect 212592 484452 212724 484480
rect 212592 484440 212598 484452
rect 212718 484440 212724 484452
rect 212776 484440 212782 484492
rect 195146 484372 195152 484424
rect 195204 484412 195210 484424
rect 197078 484412 197084 484424
rect 195204 484384 197084 484412
rect 195204 484372 195210 484384
rect 197078 484372 197084 484384
rect 197136 484372 197142 484424
rect 201954 484372 201960 484424
rect 202012 484412 202018 484424
rect 203978 484412 203984 484424
rect 202012 484384 203984 484412
rect 202012 484372 202018 484384
rect 203978 484372 203984 484384
rect 204036 484372 204042 484424
rect 211890 484372 211896 484424
rect 211948 484412 211954 484424
rect 212902 484412 212908 484424
rect 211948 484384 212908 484412
rect 211948 484372 211954 484384
rect 212902 484372 212908 484384
rect 212960 484372 212966 484424
rect 213362 484372 213368 484424
rect 213420 484412 213426 484424
rect 216214 484412 216220 484424
rect 213420 484384 216220 484412
rect 213420 484372 213426 484384
rect 216214 484372 216220 484384
rect 216272 484372 216278 484424
rect 216582 484372 216588 484424
rect 216640 484412 216646 484424
rect 219158 484412 219164 484424
rect 216640 484384 219164 484412
rect 216640 484372 216646 484384
rect 219158 484372 219164 484384
rect 219216 484372 219222 484424
rect 219986 484372 219992 484424
rect 220044 484412 220050 484424
rect 222654 484412 222660 484424
rect 220044 484384 222660 484412
rect 220044 484372 220050 484384
rect 222654 484372 222660 484384
rect 222712 484372 222718 484424
rect 129826 484304 129832 484356
rect 129884 484344 129890 484356
rect 130010 484344 130016 484356
rect 129884 484316 130016 484344
rect 129884 484304 129890 484316
rect 130010 484304 130016 484316
rect 130068 484304 130074 484356
rect 129734 484236 129740 484288
rect 129792 484276 129798 484288
rect 129918 484276 129924 484288
rect 129792 484248 129924 484276
rect 129792 484236 129798 484248
rect 129918 484236 129924 484248
rect 129976 484236 129982 484288
rect 281626 484236 281632 484288
rect 281684 484236 281690 484288
rect 70486 484168 70492 484220
rect 70544 484208 70550 484220
rect 71222 484208 71228 484220
rect 70544 484180 71228 484208
rect 70544 484168 70550 484180
rect 71222 484168 71228 484180
rect 71280 484168 71286 484220
rect 78674 484168 78680 484220
rect 78732 484208 78738 484220
rect 79134 484208 79140 484220
rect 78732 484180 79140 484208
rect 78732 484168 78738 484180
rect 79134 484168 79140 484180
rect 79192 484168 79198 484220
rect 172514 484168 172520 484220
rect 172572 484208 172578 484220
rect 173526 484208 173532 484220
rect 172572 484180 173532 484208
rect 172572 484168 172578 484180
rect 173526 484168 173532 484180
rect 173584 484168 173590 484220
rect 191834 484168 191840 484220
rect 191892 484208 191898 484220
rect 192386 484208 192392 484220
rect 191892 484180 192392 484208
rect 191892 484168 191898 484180
rect 192386 484168 192392 484180
rect 192444 484168 192450 484220
rect 193214 484168 193220 484220
rect 193272 484208 193278 484220
rect 194134 484208 194140 484220
rect 193272 484180 194140 484208
rect 193272 484168 193278 484180
rect 194134 484168 194140 484180
rect 194192 484168 194198 484220
rect 198734 484168 198740 484220
rect 198792 484208 198798 484220
rect 199470 484208 199476 484220
rect 198792 484180 199476 484208
rect 198792 484168 198798 484180
rect 199470 484168 199476 484180
rect 199528 484168 199534 484220
rect 205726 484168 205732 484220
rect 205784 484208 205790 484220
rect 206462 484208 206468 484220
rect 205784 484180 206468 484208
rect 205784 484168 205790 484180
rect 206462 484168 206468 484180
rect 206520 484168 206526 484220
rect 219526 484168 219532 484220
rect 219584 484208 219590 484220
rect 220078 484208 220084 484220
rect 219584 484180 220084 484208
rect 219584 484168 219590 484180
rect 220078 484168 220084 484180
rect 220136 484168 220142 484220
rect 70394 484100 70400 484152
rect 70452 484140 70458 484152
rect 70854 484140 70860 484152
rect 70452 484112 70860 484140
rect 70452 484100 70458 484112
rect 70854 484100 70860 484112
rect 70912 484100 70918 484152
rect 71866 484100 71872 484152
rect 71924 484140 71930 484152
rect 72602 484140 72608 484152
rect 71924 484112 72608 484140
rect 71924 484100 71930 484112
rect 72602 484100 72608 484112
rect 72660 484100 72666 484152
rect 74626 484100 74632 484152
rect 74684 484140 74690 484152
rect 75270 484140 75276 484152
rect 74684 484112 75276 484140
rect 74684 484100 74690 484112
rect 75270 484100 75276 484112
rect 75328 484100 75334 484152
rect 75914 484100 75920 484152
rect 75972 484140 75978 484152
rect 76558 484140 76564 484152
rect 75972 484112 76564 484140
rect 75972 484100 75978 484112
rect 76558 484100 76564 484112
rect 76616 484100 76622 484152
rect 78766 484100 78772 484152
rect 78824 484140 78830 484152
rect 79686 484140 79692 484152
rect 78824 484112 79692 484140
rect 78824 484100 78830 484112
rect 79686 484100 79692 484112
rect 79744 484100 79750 484152
rect 93854 484100 93860 484152
rect 93912 484140 93918 484152
rect 94590 484140 94596 484152
rect 93912 484112 94596 484140
rect 93912 484100 93918 484112
rect 94590 484100 94596 484112
rect 94648 484100 94654 484152
rect 131114 484100 131120 484152
rect 131172 484140 131178 484152
rect 132126 484140 132132 484152
rect 131172 484112 132132 484140
rect 131172 484100 131178 484112
rect 132126 484100 132132 484112
rect 132184 484100 132190 484152
rect 132586 484100 132592 484152
rect 132644 484140 132650 484152
rect 133414 484140 133420 484152
rect 132644 484112 133420 484140
rect 132644 484100 132650 484112
rect 133414 484100 133420 484112
rect 133472 484100 133478 484152
rect 133874 484100 133880 484152
rect 133932 484140 133938 484152
rect 134702 484140 134708 484152
rect 133932 484112 134708 484140
rect 133932 484100 133938 484112
rect 134702 484100 134708 484112
rect 134760 484100 134766 484152
rect 139394 484100 139400 484152
rect 139452 484140 139458 484152
rect 140038 484140 140044 484152
rect 139452 484112 140044 484140
rect 139452 484100 139458 484112
rect 140038 484100 140044 484112
rect 140096 484100 140102 484152
rect 140866 484100 140872 484152
rect 140924 484140 140930 484152
rect 141326 484140 141332 484152
rect 140924 484112 141332 484140
rect 140924 484100 140930 484112
rect 141326 484100 141332 484112
rect 141384 484100 141390 484152
rect 142154 484100 142160 484152
rect 142212 484140 142218 484152
rect 142614 484140 142620 484152
rect 142212 484112 142620 484140
rect 142212 484100 142218 484112
rect 142614 484100 142620 484112
rect 142672 484100 142678 484152
rect 143534 484100 143540 484152
rect 143592 484140 143598 484152
rect 144454 484140 144460 484152
rect 143592 484112 144460 484140
rect 143592 484100 143598 484112
rect 144454 484100 144460 484112
rect 144512 484100 144518 484152
rect 147674 484100 147680 484152
rect 147732 484140 147738 484152
rect 148318 484140 148324 484152
rect 147732 484112 148324 484140
rect 147732 484100 147738 484112
rect 148318 484100 148324 484112
rect 148376 484100 148382 484152
rect 167086 484100 167092 484152
rect 167144 484140 167150 484152
rect 167730 484140 167736 484152
rect 167144 484112 167736 484140
rect 167144 484100 167150 484112
rect 167730 484100 167736 484112
rect 167788 484100 167794 484152
rect 171134 484100 171140 484152
rect 171192 484140 171198 484152
rect 171686 484140 171692 484152
rect 171192 484112 171692 484140
rect 171192 484100 171198 484112
rect 171686 484100 171692 484112
rect 171744 484100 171750 484152
rect 172606 484100 172612 484152
rect 172664 484140 172670 484152
rect 172974 484140 172980 484152
rect 172664 484112 172980 484140
rect 172664 484100 172670 484112
rect 172974 484100 172980 484112
rect 173032 484100 173038 484152
rect 175274 484100 175280 484152
rect 175332 484140 175338 484152
rect 175734 484140 175740 484152
rect 175332 484112 175740 484140
rect 175332 484100 175338 484112
rect 175734 484100 175740 484112
rect 175792 484100 175798 484152
rect 186314 484100 186320 484152
rect 186372 484140 186378 484152
rect 187142 484140 187148 484152
rect 186372 484112 187148 484140
rect 186372 484100 186378 484112
rect 187142 484100 187148 484112
rect 187200 484100 187206 484152
rect 187786 484100 187792 484152
rect 187844 484140 187850 484152
rect 188430 484140 188436 484152
rect 187844 484112 188436 484140
rect 187844 484100 187850 484112
rect 188430 484100 188436 484112
rect 188488 484100 188494 484152
rect 190454 484100 190460 484152
rect 190512 484140 190518 484152
rect 191006 484140 191012 484152
rect 190512 484112 191012 484140
rect 190512 484100 190518 484112
rect 191006 484100 191012 484112
rect 191064 484100 191070 484152
rect 191926 484100 191932 484152
rect 191984 484140 191990 484152
rect 192110 484140 192116 484152
rect 191984 484112 192116 484140
rect 191984 484100 191990 484112
rect 192110 484100 192116 484112
rect 192168 484100 192174 484152
rect 193306 484100 193312 484152
rect 193364 484140 193370 484152
rect 193766 484140 193772 484152
rect 193364 484112 193772 484140
rect 193364 484100 193370 484112
rect 193766 484100 193772 484112
rect 193824 484100 193830 484152
rect 197446 484100 197452 484152
rect 197504 484140 197510 484152
rect 198182 484140 198188 484152
rect 197504 484112 198188 484140
rect 197504 484100 197510 484112
rect 198182 484100 198188 484112
rect 198240 484100 198246 484152
rect 201586 484100 201592 484152
rect 201644 484140 201650 484152
rect 202046 484140 202052 484152
rect 201644 484112 202052 484140
rect 201644 484100 201650 484112
rect 202046 484100 202052 484112
rect 202104 484100 202110 484152
rect 204438 484100 204444 484152
rect 204496 484140 204502 484152
rect 205174 484140 205180 484152
rect 204496 484112 205180 484140
rect 204496 484100 204502 484112
rect 205174 484100 205180 484112
rect 205232 484100 205238 484152
rect 205634 484100 205640 484152
rect 205692 484140 205698 484152
rect 206094 484140 206100 484152
rect 205692 484112 206100 484140
rect 205692 484100 205698 484112
rect 206094 484100 206100 484112
rect 206152 484100 206158 484152
rect 207014 484100 207020 484152
rect 207072 484140 207078 484152
rect 207750 484140 207756 484152
rect 207072 484112 207756 484140
rect 207072 484100 207078 484112
rect 207750 484100 207756 484112
rect 207808 484100 207814 484152
rect 208486 484100 208492 484152
rect 208544 484140 208550 484152
rect 209130 484140 209136 484152
rect 208544 484112 209136 484140
rect 208544 484100 208550 484112
rect 209130 484100 209136 484112
rect 209188 484100 209194 484152
rect 209774 484100 209780 484152
rect 209832 484140 209838 484152
rect 210510 484140 210516 484152
rect 209832 484112 210516 484140
rect 209832 484100 209838 484112
rect 210510 484100 210516 484112
rect 210568 484100 210574 484152
rect 212626 484100 212632 484152
rect 212684 484140 212690 484152
rect 213454 484140 213460 484152
rect 212684 484112 213460 484140
rect 212684 484100 212690 484112
rect 213454 484100 213460 484112
rect 213512 484100 213518 484152
rect 213914 484100 213920 484152
rect 213972 484140 213978 484152
rect 214926 484140 214932 484152
rect 213972 484112 214932 484140
rect 213972 484100 213978 484112
rect 214926 484100 214932 484112
rect 214984 484100 214990 484152
rect 216766 484100 216772 484152
rect 216824 484140 216830 484152
rect 217502 484140 217508 484152
rect 216824 484112 217508 484140
rect 216824 484100 216830 484112
rect 217502 484100 217508 484112
rect 217560 484100 217566 484152
rect 219434 484100 219440 484152
rect 219492 484140 219498 484152
rect 219710 484140 219716 484152
rect 219492 484112 219716 484140
rect 219492 484100 219498 484112
rect 219710 484100 219716 484112
rect 219768 484100 219774 484152
rect 223574 484100 223580 484152
rect 223632 484140 223638 484152
rect 224126 484140 224132 484152
rect 223632 484112 224132 484140
rect 223632 484100 223638 484112
rect 224126 484100 224132 484112
rect 224184 484100 224190 484152
rect 226334 484100 226340 484152
rect 226392 484140 226398 484152
rect 226702 484140 226708 484152
rect 226392 484112 226708 484140
rect 226392 484100 226398 484112
rect 226702 484100 226708 484112
rect 226760 484100 226766 484152
rect 229094 484100 229100 484152
rect 229152 484140 229158 484152
rect 229462 484140 229468 484152
rect 229152 484112 229468 484140
rect 229152 484100 229158 484112
rect 229462 484100 229468 484112
rect 229520 484100 229526 484152
rect 240226 484100 240232 484152
rect 240284 484140 240290 484152
rect 240870 484140 240876 484152
rect 240284 484112 240876 484140
rect 240284 484100 240290 484112
rect 240870 484100 240876 484112
rect 240928 484100 240934 484152
rect 241514 484100 241520 484152
rect 241572 484140 241578 484152
rect 242158 484140 242164 484152
rect 241572 484112 242164 484140
rect 241572 484100 241578 484112
rect 242158 484100 242164 484112
rect 242216 484100 242222 484152
rect 263686 484100 263692 484152
rect 263744 484140 263750 484152
rect 264238 484140 264244 484152
rect 263744 484112 264244 484140
rect 263744 484100 263750 484112
rect 264238 484100 264244 484112
rect 264296 484100 264302 484152
rect 264974 484100 264980 484152
rect 265032 484140 265038 484152
rect 265526 484140 265532 484152
rect 265032 484112 265532 484140
rect 265032 484100 265038 484112
rect 265526 484100 265532 484112
rect 265584 484100 265590 484152
rect 269114 484100 269120 484152
rect 269172 484140 269178 484152
rect 269942 484140 269948 484152
rect 269172 484112 269948 484140
rect 269172 484100 269178 484112
rect 269942 484100 269948 484112
rect 270000 484100 270006 484152
rect 270494 484100 270500 484152
rect 270552 484140 270558 484152
rect 270862 484140 270868 484152
rect 270552 484112 270868 484140
rect 270552 484100 270558 484112
rect 270862 484100 270868 484112
rect 270920 484100 270926 484152
rect 271966 484100 271972 484152
rect 272024 484140 272030 484152
rect 272518 484140 272524 484152
rect 272024 484112 272524 484140
rect 272024 484100 272030 484112
rect 272518 484100 272524 484112
rect 272576 484100 272582 484152
rect 273346 484100 273352 484152
rect 273404 484140 273410 484152
rect 273806 484140 273812 484152
rect 273404 484112 273812 484140
rect 273404 484100 273410 484112
rect 273806 484100 273812 484112
rect 273864 484100 273870 484152
rect 281644 484072 281672 484236
rect 293954 484100 293960 484152
rect 294012 484140 294018 484152
rect 371694 484140 371700 484152
rect 294012 484112 371700 484140
rect 294012 484100 294018 484112
rect 371694 484100 371700 484112
rect 371752 484100 371758 484152
rect 359458 484072 359464 484084
rect 281644 484044 359464 484072
rect 359458 484032 359464 484044
rect 359516 484032 359522 484084
rect 129826 483964 129832 484016
rect 129884 484004 129890 484016
rect 130286 484004 130292 484016
rect 129884 483976 130292 484004
rect 129884 483964 129890 483976
rect 130286 483964 130292 483976
rect 130344 483964 130350 484016
rect 202966 483964 202972 484016
rect 203024 484004 203030 484016
rect 203886 484004 203892 484016
rect 203024 483976 203892 484004
rect 203024 483964 203030 483976
rect 203886 483964 203892 483976
rect 203944 483964 203950 484016
rect 226426 483964 226432 484016
rect 226484 484004 226490 484016
rect 227254 484004 227260 484016
rect 226484 483976 227260 484004
rect 226484 483964 226490 483976
rect 227254 483964 227260 483976
rect 227312 483964 227318 484016
rect 280062 483964 280068 484016
rect 280120 484004 280126 484016
rect 362770 484004 362776 484016
rect 280120 483976 362776 484004
rect 280120 483964 280126 483976
rect 362770 483964 362776 483976
rect 362828 483964 362834 484016
rect 279786 483896 279792 483948
rect 279844 483936 279850 483948
rect 372338 483936 372344 483948
rect 279844 483908 372344 483936
rect 279844 483896 279850 483908
rect 372338 483896 372344 483908
rect 372396 483896 372402 483948
rect 275554 483828 275560 483880
rect 275612 483868 275618 483880
rect 370406 483868 370412 483880
rect 275612 483840 370412 483868
rect 275612 483828 275618 483840
rect 370406 483828 370412 483840
rect 370464 483828 370470 483880
rect 176562 483760 176568 483812
rect 176620 483800 176626 483812
rect 206370 483800 206376 483812
rect 176620 483772 206376 483800
rect 176620 483760 176626 483772
rect 206370 483760 206376 483772
rect 206428 483760 206434 483812
rect 260098 483760 260104 483812
rect 260156 483800 260162 483812
rect 370682 483800 370688 483812
rect 260156 483772 370688 483800
rect 260156 483760 260162 483772
rect 370682 483760 370688 483772
rect 370740 483760 370746 483812
rect 165522 483692 165528 483744
rect 165580 483732 165586 483744
rect 214558 483732 214564 483744
rect 165580 483704 214564 483732
rect 165580 483692 165586 483704
rect 214558 483692 214564 483704
rect 214616 483692 214622 483744
rect 236730 483692 236736 483744
rect 236788 483732 236794 483744
rect 362310 483732 362316 483744
rect 236788 483704 362316 483732
rect 236788 483692 236794 483704
rect 362310 483692 362316 483704
rect 362368 483692 362374 483744
rect 60642 483624 60648 483676
rect 60700 483664 60706 483676
rect 80698 483664 80704 483676
rect 60700 483636 80704 483664
rect 60700 483624 60706 483636
rect 80698 483624 80704 483636
rect 80756 483624 80762 483676
rect 161566 483624 161572 483676
rect 161624 483664 161630 483676
rect 215938 483664 215944 483676
rect 161624 483636 215944 483664
rect 161624 483624 161630 483636
rect 215938 483624 215944 483636
rect 215996 483624 216002 483676
rect 246942 483624 246948 483676
rect 247000 483664 247006 483676
rect 378778 483664 378784 483676
rect 247000 483636 378784 483664
rect 247000 483624 247006 483636
rect 378778 483624 378784 483636
rect 378836 483624 378842 483676
rect 189074 483352 189080 483404
rect 189132 483392 189138 483404
rect 189350 483392 189356 483404
rect 189132 483364 189356 483392
rect 189132 483352 189138 483364
rect 189350 483352 189356 483364
rect 189408 483352 189414 483404
rect 50430 482944 50436 482996
rect 50488 482984 50494 482996
rect 97166 482984 97172 482996
rect 50488 482956 97172 482984
rect 50488 482944 50494 482956
rect 97166 482944 97172 482956
rect 97224 482944 97230 482996
rect 48038 482876 48044 482928
rect 48096 482916 48102 482928
rect 97534 482916 97540 482928
rect 48096 482888 97540 482916
rect 48096 482876 48102 482888
rect 97534 482876 97540 482888
rect 97592 482876 97598 482928
rect 290090 482876 290096 482928
rect 290148 482916 290154 482928
rect 367002 482916 367008 482928
rect 290148 482888 367008 482916
rect 290148 482876 290154 482888
rect 367002 482876 367008 482888
rect 367060 482876 367066 482928
rect 49234 482808 49240 482860
rect 49292 482848 49298 482860
rect 97994 482848 98000 482860
rect 49292 482820 98000 482848
rect 49292 482808 49298 482820
rect 97994 482808 98000 482820
rect 98052 482808 98058 482860
rect 203702 482808 203708 482860
rect 203760 482848 203766 482860
rect 209406 482848 209412 482860
rect 203760 482820 209412 482848
rect 203760 482808 203766 482820
rect 209406 482808 209412 482820
rect 209464 482808 209470 482860
rect 274818 482808 274824 482860
rect 274876 482848 274882 482860
rect 365530 482848 365536 482860
rect 274876 482820 365536 482848
rect 274876 482808 274882 482820
rect 365530 482808 365536 482820
rect 365588 482808 365594 482860
rect 47854 482740 47860 482792
rect 47912 482780 47918 482792
rect 111702 482780 111708 482792
rect 47912 482752 111708 482780
rect 47912 482740 47918 482752
rect 111702 482740 111708 482752
rect 111760 482740 111766 482792
rect 271782 482740 271788 482792
rect 271840 482780 271846 482792
rect 366910 482780 366916 482792
rect 271840 482752 366916 482780
rect 271840 482740 271846 482752
rect 366910 482740 366916 482752
rect 366968 482740 366974 482792
rect 46566 482672 46572 482724
rect 46624 482712 46630 482724
rect 111242 482712 111248 482724
rect 46624 482684 111248 482712
rect 46624 482672 46630 482684
rect 111242 482672 111248 482684
rect 111300 482672 111306 482724
rect 159266 482672 159272 482724
rect 159324 482712 159330 482724
rect 207750 482712 207756 482724
rect 159324 482684 207756 482712
rect 159324 482672 159330 482684
rect 207750 482672 207756 482684
rect 207808 482672 207814 482724
rect 276658 482672 276664 482724
rect 276716 482712 276722 482724
rect 374454 482712 374460 482724
rect 276716 482684 374460 482712
rect 276716 482672 276722 482684
rect 374454 482672 374460 482684
rect 374512 482672 374518 482724
rect 50522 482604 50528 482656
rect 50580 482644 50586 482656
rect 115658 482644 115664 482656
rect 50580 482616 115664 482644
rect 50580 482604 50586 482616
rect 115658 482604 115664 482616
rect 115716 482604 115722 482656
rect 135622 482604 135628 482656
rect 135680 482644 135686 482656
rect 141786 482644 141792 482656
rect 135680 482616 141792 482644
rect 135680 482604 135686 482616
rect 141786 482604 141792 482616
rect 141844 482604 141850 482656
rect 160554 482604 160560 482656
rect 160612 482644 160618 482656
rect 211798 482644 211804 482656
rect 160612 482616 211804 482644
rect 160612 482604 160618 482616
rect 211798 482604 211804 482616
rect 211856 482604 211862 482656
rect 276842 482604 276848 482656
rect 276900 482644 276906 482656
rect 375834 482644 375840 482656
rect 276900 482616 375840 482644
rect 276900 482604 276906 482616
rect 375834 482604 375840 482616
rect 375892 482604 375898 482656
rect 46382 482536 46388 482588
rect 46440 482576 46446 482588
rect 112530 482576 112536 482588
rect 46440 482548 112536 482576
rect 46440 482536 46446 482548
rect 112530 482536 112536 482548
rect 112588 482536 112594 482588
rect 138474 482536 138480 482588
rect 138532 482576 138538 482588
rect 200298 482576 200304 482588
rect 138532 482548 200304 482576
rect 138532 482536 138538 482548
rect 200298 482536 200304 482548
rect 200356 482536 200362 482588
rect 261386 482536 261392 482588
rect 261444 482576 261450 482588
rect 368014 482576 368020 482588
rect 261444 482548 368020 482576
rect 261444 482536 261450 482548
rect 368014 482536 368020 482548
rect 368072 482536 368078 482588
rect 46474 482468 46480 482520
rect 46532 482508 46538 482520
rect 112070 482508 112076 482520
rect 46532 482480 112076 482508
rect 46532 482468 46538 482480
rect 112070 482468 112076 482480
rect 112128 482468 112134 482520
rect 136818 482468 136824 482520
rect 136876 482508 136882 482520
rect 199102 482508 199108 482520
rect 136876 482480 199108 482508
rect 136876 482468 136882 482480
rect 199102 482468 199108 482480
rect 199160 482468 199166 482520
rect 257522 482468 257528 482520
rect 257580 482508 257586 482520
rect 366634 482508 366640 482520
rect 257580 482480 366640 482508
rect 257580 482468 257586 482480
rect 366634 482468 366640 482480
rect 366692 482468 366698 482520
rect 49142 482400 49148 482452
rect 49200 482440 49206 482452
rect 115198 482440 115204 482452
rect 49200 482412 115204 482440
rect 49200 482400 49206 482412
rect 115198 482400 115204 482412
rect 115256 482400 115262 482452
rect 140774 482400 140780 482452
rect 140832 482440 140838 482452
rect 141694 482440 141700 482452
rect 140832 482412 141700 482440
rect 140832 482400 140838 482412
rect 141694 482400 141700 482412
rect 141752 482400 141758 482452
rect 141786 482400 141792 482452
rect 141844 482440 141850 482452
rect 197998 482440 198004 482452
rect 141844 482412 198004 482440
rect 141844 482400 141850 482412
rect 197998 482400 198004 482412
rect 198056 482400 198062 482452
rect 244642 482400 244648 482452
rect 244700 482440 244706 482452
rect 373350 482440 373356 482452
rect 244700 482412 373356 482440
rect 244700 482400 244706 482412
rect 373350 482400 373356 482412
rect 373408 482400 373414 482452
rect 48130 482332 48136 482384
rect 48188 482372 48194 482384
rect 119614 482372 119620 482384
rect 48188 482344 119620 482372
rect 48188 482332 48194 482344
rect 119614 482332 119620 482344
rect 119672 482332 119678 482384
rect 137922 482332 137928 482384
rect 137980 482372 137986 482384
rect 201862 482372 201868 482384
rect 137980 482344 201868 482372
rect 137980 482332 137986 482344
rect 201862 482332 201868 482344
rect 201920 482332 201926 482384
rect 248322 482332 248328 482384
rect 248380 482372 248386 482384
rect 378962 482372 378968 482384
rect 248380 482344 378968 482372
rect 248380 482332 248386 482344
rect 378962 482332 378968 482344
rect 379020 482332 379026 482384
rect 46658 482264 46664 482316
rect 46716 482304 46722 482316
rect 120074 482304 120080 482316
rect 46716 482276 120080 482304
rect 46716 482264 46722 482276
rect 120074 482264 120080 482276
rect 120132 482264 120138 482316
rect 138566 482264 138572 482316
rect 138624 482304 138630 482316
rect 207290 482304 207296 482316
rect 138624 482276 207296 482304
rect 138624 482264 138630 482276
rect 207290 482264 207296 482276
rect 207348 482264 207354 482316
rect 222562 482264 222568 482316
rect 222620 482304 222626 482316
rect 376018 482304 376024 482316
rect 222620 482276 376024 482304
rect 222620 482264 222626 482276
rect 376018 482264 376024 482276
rect 376076 482264 376082 482316
rect 51902 482196 51908 482248
rect 51960 482236 51966 482248
rect 98454 482236 98460 482248
rect 51960 482208 98460 482236
rect 51960 482196 51966 482208
rect 98454 482196 98460 482208
rect 98512 482196 98518 482248
rect 54846 482128 54852 482180
rect 54904 482168 54910 482180
rect 96706 482168 96712 482180
rect 54904 482140 96712 482168
rect 54904 482128 54910 482140
rect 96706 482128 96712 482140
rect 96764 482128 96770 482180
rect 58710 482060 58716 482112
rect 58768 482100 58774 482112
rect 96246 482100 96252 482112
rect 58768 482072 96252 482100
rect 58768 482060 58774 482072
rect 96246 482060 96252 482072
rect 96304 482060 96310 482112
rect 189166 481720 189172 481772
rect 189224 481760 189230 481772
rect 189718 481760 189724 481772
rect 189224 481732 189724 481760
rect 189224 481720 189230 481732
rect 189718 481720 189724 481732
rect 189776 481720 189782 481772
rect 291286 481448 291292 481500
rect 291344 481488 291350 481500
rect 291470 481488 291476 481500
rect 291344 481460 291476 481488
rect 291344 481448 291350 481460
rect 291470 481448 291476 481460
rect 291528 481448 291534 481500
rect 295518 481448 295524 481500
rect 295576 481488 295582 481500
rect 295702 481488 295708 481500
rect 295576 481460 295708 481488
rect 295576 481448 295582 481460
rect 295702 481448 295708 481460
rect 295760 481448 295766 481500
rect 285490 481380 285496 481432
rect 285548 481420 285554 481432
rect 359734 481420 359740 481432
rect 285548 481392 359740 481420
rect 285548 481380 285554 481392
rect 359734 481380 359740 481392
rect 359792 481380 359798 481432
rect 281442 481312 281448 481364
rect 281500 481352 281506 481364
rect 357066 481352 357072 481364
rect 281500 481324 357072 481352
rect 281500 481312 281506 481324
rect 357066 481312 357072 481324
rect 357124 481312 357130 481364
rect 269022 481244 269028 481296
rect 269080 481284 269086 481296
rect 361390 481284 361396 481296
rect 269080 481256 361396 481284
rect 269080 481244 269086 481256
rect 361390 481244 361396 481256
rect 361448 481244 361454 481296
rect 261202 481176 261208 481228
rect 261260 481216 261266 481228
rect 358354 481216 358360 481228
rect 261260 481188 358360 481216
rect 261260 481176 261266 481188
rect 358354 481176 358360 481188
rect 358412 481176 358418 481228
rect 251358 481108 251364 481160
rect 251416 481148 251422 481160
rect 251542 481148 251548 481160
rect 251416 481120 251548 481148
rect 251416 481108 251422 481120
rect 251542 481108 251548 481120
rect 251600 481108 251606 481160
rect 269298 481108 269304 481160
rect 269356 481148 269362 481160
rect 377490 481148 377496 481160
rect 269356 481120 377496 481148
rect 269356 481108 269362 481120
rect 377490 481108 377496 481120
rect 377548 481108 377554 481160
rect 67726 481040 67732 481092
rect 67784 481080 67790 481092
rect 67910 481080 67916 481092
rect 67784 481052 67916 481080
rect 67784 481040 67790 481052
rect 67910 481040 67916 481052
rect 67968 481040 67974 481092
rect 179598 481040 179604 481092
rect 179656 481080 179662 481092
rect 179782 481080 179788 481092
rect 179656 481052 179788 481080
rect 179656 481040 179662 481052
rect 179782 481040 179788 481052
rect 179840 481040 179846 481092
rect 182358 481040 182364 481092
rect 182416 481080 182422 481092
rect 182542 481080 182548 481092
rect 182416 481052 182548 481080
rect 182416 481040 182422 481052
rect 182542 481040 182548 481052
rect 182600 481040 182606 481092
rect 243078 481040 243084 481092
rect 243136 481080 243142 481092
rect 370498 481080 370504 481092
rect 243136 481052 370504 481080
rect 243136 481040 243142 481052
rect 370498 481040 370504 481052
rect 370556 481040 370562 481092
rect 57882 480972 57888 481024
rect 57940 481012 57946 481024
rect 114278 481012 114284 481024
rect 57940 480984 114284 481012
rect 57940 480972 57946 480984
rect 114278 480972 114284 480984
rect 114336 480972 114342 481024
rect 159082 480972 159088 481024
rect 159140 481012 159146 481024
rect 209038 481012 209044 481024
rect 159140 480984 209044 481012
rect 159140 480972 159146 480984
rect 209038 480972 209044 480984
rect 209096 480972 209102 481024
rect 248046 480972 248052 481024
rect 248104 481012 248110 481024
rect 376110 481012 376116 481024
rect 248104 480984 376116 481012
rect 248104 480972 248110 480984
rect 376110 480972 376116 480984
rect 376168 480972 376174 481024
rect 3786 480904 3792 480956
rect 3844 480944 3850 480956
rect 434806 480944 434812 480956
rect 3844 480916 434812 480944
rect 3844 480904 3850 480916
rect 434806 480904 434812 480916
rect 434864 480904 434870 480956
rect 62114 480836 62120 480888
rect 62172 480876 62178 480888
rect 62942 480876 62948 480888
rect 62172 480848 62948 480876
rect 62172 480836 62178 480848
rect 62942 480836 62948 480848
rect 63000 480836 63006 480888
rect 69106 480836 69112 480888
rect 69164 480876 69170 480888
rect 69934 480876 69940 480888
rect 69164 480848 69940 480876
rect 69164 480836 69170 480848
rect 69934 480836 69940 480848
rect 69992 480836 69998 480888
rect 81526 480836 81532 480888
rect 81584 480876 81590 480888
rect 82262 480876 82268 480888
rect 81584 480848 82268 480876
rect 81584 480836 81590 480848
rect 82262 480836 82268 480848
rect 82320 480836 82326 480888
rect 82814 480836 82820 480888
rect 82872 480876 82878 480888
rect 83550 480876 83556 480888
rect 82872 480848 83556 480876
rect 82872 480836 82878 480848
rect 83550 480836 83556 480848
rect 83608 480836 83614 480888
rect 84286 480836 84292 480888
rect 84344 480876 84350 480888
rect 84930 480876 84936 480888
rect 84344 480848 84936 480876
rect 84344 480836 84350 480848
rect 84930 480836 84936 480848
rect 84988 480836 84994 480888
rect 85574 480836 85580 480888
rect 85632 480876 85638 480888
rect 86310 480876 86316 480888
rect 85632 480848 86316 480876
rect 85632 480836 85638 480848
rect 86310 480836 86316 480848
rect 86368 480836 86374 480888
rect 99466 480836 99472 480888
rect 99524 480876 99530 480888
rect 100294 480876 100300 480888
rect 99524 480848 100300 480876
rect 99524 480836 99530 480848
rect 100294 480836 100300 480848
rect 100352 480836 100358 480888
rect 100754 480836 100760 480888
rect 100812 480876 100818 480888
rect 101582 480876 101588 480888
rect 100812 480848 101588 480876
rect 100812 480836 100818 480848
rect 101582 480836 101588 480848
rect 101640 480836 101646 480888
rect 106366 480836 106372 480888
rect 106424 480876 106430 480888
rect 106918 480876 106924 480888
rect 106424 480848 106924 480876
rect 106424 480836 106430 480848
rect 106918 480836 106924 480848
rect 106976 480836 106982 480888
rect 113266 480836 113272 480888
rect 113324 480876 113330 480888
rect 113542 480876 113548 480888
rect 113324 480848 113548 480876
rect 113324 480836 113330 480848
rect 113542 480836 113548 480848
rect 113600 480836 113606 480888
rect 125594 480836 125600 480888
rect 125652 480876 125658 480888
rect 126330 480876 126336 480888
rect 125652 480848 126336 480876
rect 125652 480836 125658 480848
rect 126330 480836 126336 480848
rect 126388 480836 126394 480888
rect 161474 480836 161480 480888
rect 161532 480876 161538 480888
rect 161934 480876 161940 480888
rect 161532 480848 161940 480876
rect 161532 480836 161538 480848
rect 161934 480836 161940 480848
rect 161992 480836 161998 480888
rect 176654 480836 176660 480888
rect 176712 480876 176718 480888
rect 177390 480876 177396 480888
rect 176712 480848 177396 480876
rect 176712 480836 176718 480848
rect 177390 480836 177396 480848
rect 177448 480836 177454 480888
rect 180794 480836 180800 480888
rect 180852 480876 180858 480888
rect 181438 480876 181444 480888
rect 180852 480848 181444 480876
rect 180852 480836 180858 480848
rect 181438 480836 181444 480848
rect 181496 480836 181502 480888
rect 182174 480836 182180 480888
rect 182232 480876 182238 480888
rect 182726 480876 182732 480888
rect 182232 480848 182732 480876
rect 182232 480836 182238 480848
rect 182726 480836 182732 480848
rect 182784 480836 182790 480888
rect 183554 480836 183560 480888
rect 183612 480876 183618 480888
rect 184382 480876 184388 480888
rect 183612 480848 184388 480876
rect 183612 480836 183618 480848
rect 184382 480836 184388 480848
rect 184440 480836 184446 480888
rect 248414 480836 248420 480888
rect 248472 480876 248478 480888
rect 248782 480876 248788 480888
rect 248472 480848 248788 480876
rect 248472 480836 248478 480848
rect 248782 480836 248788 480848
rect 248840 480836 248846 480888
rect 249794 480836 249800 480888
rect 249852 480876 249858 480888
rect 250530 480876 250536 480888
rect 249852 480848 250536 480876
rect 249852 480836 249858 480848
rect 250530 480836 250536 480848
rect 250588 480836 250594 480888
rect 251174 480836 251180 480888
rect 251232 480876 251238 480888
rect 251910 480876 251916 480888
rect 251232 480848 251916 480876
rect 251232 480836 251238 480848
rect 251910 480836 251916 480848
rect 251968 480836 251974 480888
rect 252554 480836 252560 480888
rect 252612 480876 252618 480888
rect 253198 480876 253204 480888
rect 252612 480848 253204 480876
rect 252612 480836 252618 480848
rect 253198 480836 253204 480848
rect 253256 480836 253262 480888
rect 258074 480836 258080 480888
rect 258132 480876 258138 480888
rect 258534 480876 258540 480888
rect 258132 480848 258540 480876
rect 258132 480836 258138 480848
rect 258534 480836 258540 480848
rect 258592 480836 258598 480888
rect 262306 480836 262312 480888
rect 262364 480876 262370 480888
rect 262858 480876 262864 480888
rect 262364 480848 262864 480876
rect 262364 480836 262370 480848
rect 262858 480836 262864 480848
rect 262916 480836 262922 480888
rect 282914 480836 282920 480888
rect 282972 480876 282978 480888
rect 283558 480876 283564 480888
rect 282972 480848 283564 480876
rect 282972 480836 282978 480848
rect 283558 480836 283564 480848
rect 283616 480836 283622 480888
rect 284294 480836 284300 480888
rect 284352 480876 284358 480888
rect 284478 480876 284484 480888
rect 284352 480848 284484 480876
rect 284352 480836 284358 480848
rect 284478 480836 284484 480848
rect 284536 480836 284542 480888
rect 287054 480836 287060 480888
rect 287112 480876 287118 480888
rect 287974 480876 287980 480888
rect 287112 480848 287980 480876
rect 287112 480836 287118 480848
rect 287974 480836 287980 480848
rect 288032 480836 288038 480888
rect 289814 480836 289820 480888
rect 289872 480876 289878 480888
rect 290550 480876 290556 480888
rect 289872 480848 290556 480876
rect 289872 480836 289878 480848
rect 290550 480836 290556 480848
rect 290608 480836 290614 480888
rect 293954 480836 293960 480888
rect 294012 480876 294018 480888
rect 294598 480876 294604 480888
rect 294012 480848 294604 480876
rect 294012 480836 294018 480848
rect 294598 480836 294604 480848
rect 294656 480836 294662 480888
rect 295334 480836 295340 480888
rect 295392 480876 295398 480888
rect 295886 480876 295892 480888
rect 295392 480848 295892 480876
rect 295392 480836 295398 480848
rect 295886 480836 295892 480848
rect 295944 480836 295950 480888
rect 296714 480836 296720 480888
rect 296772 480876 296778 480888
rect 297174 480876 297180 480888
rect 296772 480848 297180 480876
rect 296772 480836 296778 480848
rect 297174 480836 297180 480848
rect 297232 480836 297238 480888
rect 179506 480700 179512 480752
rect 179564 480740 179570 480752
rect 180058 480740 180064 480752
rect 179564 480712 180064 480740
rect 179564 480700 179570 480712
rect 180058 480700 180064 480712
rect 180116 480700 180122 480752
rect 220814 480224 220820 480276
rect 220872 480264 220878 480276
rect 220998 480264 221004 480276
rect 220872 480236 221004 480264
rect 220872 480224 220878 480236
rect 220998 480224 221004 480236
rect 221056 480224 221062 480276
rect 57238 480156 57244 480208
rect 57296 480196 57302 480208
rect 123018 480196 123024 480208
rect 57296 480168 123024 480196
rect 57296 480156 57302 480168
rect 123018 480156 123024 480168
rect 123076 480156 123082 480208
rect 46750 480088 46756 480140
rect 46808 480128 46814 480140
rect 116210 480128 116216 480140
rect 46808 480100 116216 480128
rect 46808 480088 46814 480100
rect 116210 480088 116216 480100
rect 116268 480088 116274 480140
rect 293310 480088 293316 480140
rect 293368 480128 293374 480140
rect 370314 480128 370320 480140
rect 293368 480100 370320 480128
rect 293368 480088 293374 480100
rect 370314 480088 370320 480100
rect 370372 480088 370378 480140
rect 48222 480020 48228 480072
rect 48280 480060 48286 480072
rect 117498 480060 117504 480072
rect 48280 480032 117504 480060
rect 48280 480020 48286 480032
rect 117498 480020 117504 480032
rect 117556 480020 117562 480072
rect 299474 480020 299480 480072
rect 299532 480060 299538 480072
rect 379238 480060 379244 480072
rect 299532 480032 379244 480060
rect 299532 480020 299538 480032
rect 379238 480020 379244 480032
rect 379296 480020 379302 480072
rect 59722 479952 59728 480004
rect 59780 479992 59786 480004
rect 129826 479992 129832 480004
rect 59780 479964 129832 479992
rect 59780 479952 59786 479964
rect 129826 479952 129832 479964
rect 129884 479952 129890 480004
rect 278774 479952 278780 480004
rect 278832 479992 278838 480004
rect 365622 479992 365628 480004
rect 278832 479964 365628 479992
rect 278832 479952 278838 479964
rect 365622 479952 365628 479964
rect 365680 479952 365686 480004
rect 45462 479884 45468 479936
rect 45520 479924 45526 479936
rect 117590 479924 117596 479936
rect 45520 479896 117596 479924
rect 45520 479884 45526 479896
rect 117590 479884 117596 479896
rect 117648 479884 117654 479936
rect 256326 479884 256332 479936
rect 256384 479924 256390 479936
rect 356882 479924 356888 479936
rect 256384 479896 356888 479924
rect 256384 479884 256390 479896
rect 356882 479884 356888 479896
rect 356940 479884 356946 479936
rect 43714 479816 43720 479868
rect 43772 479856 43778 479868
rect 117958 479856 117964 479868
rect 43772 479828 117964 479856
rect 43772 479816 43778 479828
rect 117958 479816 117964 479828
rect 118016 479816 118022 479868
rect 265894 479816 265900 479868
rect 265952 479856 265958 479868
rect 366726 479856 366732 479868
rect 265952 479828 366732 479856
rect 265952 479816 265958 479828
rect 366726 479816 366732 479828
rect 366784 479816 366790 479868
rect 47670 479748 47676 479800
rect 47728 479788 47734 479800
rect 129734 479788 129740 479800
rect 47728 479760 129740 479788
rect 47728 479748 47734 479760
rect 129734 479748 129740 479760
rect 129792 479748 129798 479800
rect 259546 479748 259552 479800
rect 259604 479788 259610 479800
rect 365346 479788 365352 479800
rect 259604 479760 365352 479788
rect 259604 479748 259610 479760
rect 365346 479748 365352 479760
rect 365404 479748 365410 479800
rect 47762 479680 47768 479732
rect 47820 479720 47826 479732
rect 129918 479720 129924 479732
rect 47820 479692 129924 479720
rect 47820 479680 47826 479692
rect 129918 479680 129924 479692
rect 129976 479680 129982 479732
rect 254486 479680 254492 479732
rect 254544 479720 254550 479732
rect 369486 479720 369492 479732
rect 254544 479692 369492 479720
rect 254544 479680 254550 479692
rect 369486 479680 369492 479692
rect 369544 479680 369550 479732
rect 46106 479612 46112 479664
rect 46164 479652 46170 479664
rect 128906 479652 128912 479664
rect 46164 479624 128912 479652
rect 46164 479612 46170 479624
rect 128906 479612 128912 479624
rect 128964 479612 128970 479664
rect 189258 479612 189264 479664
rect 189316 479652 189322 479664
rect 200758 479652 200764 479664
rect 189316 479624 200764 479652
rect 189316 479612 189322 479624
rect 200758 479612 200764 479624
rect 200816 479612 200822 479664
rect 243446 479612 243452 479664
rect 243504 479652 243510 479664
rect 360930 479652 360936 479664
rect 243504 479624 360936 479652
rect 243504 479612 243510 479624
rect 360930 479612 360936 479624
rect 360988 479612 360994 479664
rect 47578 479544 47584 479596
rect 47636 479584 47642 479596
rect 134334 479584 134340 479596
rect 47636 479556 134340 479584
rect 47636 479544 47642 479556
rect 134334 479544 134340 479556
rect 134392 479544 134398 479596
rect 160186 479544 160192 479596
rect 160244 479584 160250 479596
rect 210510 479584 210516 479596
rect 160244 479556 210516 479584
rect 160244 479544 160250 479556
rect 210510 479544 210516 479556
rect 210568 479544 210574 479596
rect 246114 479544 246120 479596
rect 246172 479584 246178 479596
rect 369210 479584 369216 479596
rect 246172 479556 369216 479584
rect 246172 479544 246178 479556
rect 369210 479544 369216 479556
rect 369268 479544 369274 479596
rect 62390 479476 62396 479528
rect 62448 479516 62454 479528
rect 199286 479516 199292 479528
rect 62448 479488 199292 479516
rect 62448 479476 62454 479488
rect 199286 479476 199292 479488
rect 199344 479476 199350 479528
rect 238202 479476 238208 479528
rect 238260 479516 238266 479528
rect 374730 479516 374736 479528
rect 238260 479488 374736 479516
rect 238260 479476 238266 479488
rect 374730 479476 374736 479488
rect 374788 479476 374794 479528
rect 51718 479408 51724 479460
rect 51776 479448 51782 479460
rect 116118 479448 116124 479460
rect 51776 479420 116124 479448
rect 51776 479408 51782 479420
rect 116118 479408 116124 479420
rect 116176 479408 116182 479460
rect 58526 479340 58532 479392
rect 58584 479380 58590 479392
rect 123662 479380 123668 479392
rect 58584 479352 123668 479380
rect 58584 479340 58590 479352
rect 123662 479340 123668 479352
rect 123720 479340 123726 479392
rect 54754 479272 54760 479324
rect 54812 479312 54818 479324
rect 116670 479312 116676 479324
rect 54812 479284 116676 479312
rect 54812 479272 54818 479284
rect 116670 479272 116676 479284
rect 116728 479272 116734 479324
rect 107746 478524 107752 478576
rect 107804 478564 107810 478576
rect 108206 478564 108212 478576
rect 107804 478536 108212 478564
rect 107804 478524 107810 478536
rect 108206 478524 108212 478536
rect 108264 478524 108270 478576
rect 270586 478524 270592 478576
rect 270644 478564 270650 478576
rect 358538 478564 358544 478576
rect 270644 478536 358544 478564
rect 270644 478524 270650 478536
rect 358538 478524 358544 478536
rect 358596 478524 358602 478576
rect 254854 478456 254860 478508
rect 254912 478496 254918 478508
rect 358446 478496 358452 478508
rect 254912 478468 358452 478496
rect 254912 478456 254918 478468
rect 358446 478456 358452 478468
rect 358504 478456 358510 478508
rect 269390 478388 269396 478440
rect 269448 478428 269454 478440
rect 373902 478428 373908 478440
rect 269448 478400 373908 478428
rect 269448 478388 269454 478400
rect 373902 478388 373908 478400
rect 373960 478388 373966 478440
rect 252738 478320 252744 478372
rect 252796 478360 252802 478372
rect 374914 478360 374920 478372
rect 252796 478332 374920 478360
rect 252796 478320 252802 478332
rect 374914 478320 374920 478332
rect 374972 478320 374978 478372
rect 241698 478252 241704 478304
rect 241756 478292 241762 478304
rect 367830 478292 367836 478304
rect 241756 478264 367836 478292
rect 241756 478252 241762 478264
rect 367830 478252 367836 478264
rect 367888 478252 367894 478304
rect 177022 478184 177028 478236
rect 177080 478224 177086 478236
rect 204990 478224 204996 478236
rect 177080 478196 204996 478224
rect 177080 478184 177086 478196
rect 204990 478184 204996 478196
rect 205048 478184 205054 478236
rect 237466 478184 237472 478236
rect 237524 478224 237530 478236
rect 363874 478224 363880 478236
rect 237524 478196 363880 478224
rect 237524 478184 237530 478196
rect 363874 478184 363880 478196
rect 363932 478184 363938 478236
rect 61654 478116 61660 478168
rect 61712 478156 61718 478168
rect 199378 478156 199384 478168
rect 61712 478128 199384 478156
rect 61712 478116 61718 478128
rect 199378 478116 199384 478128
rect 199436 478116 199442 478168
rect 205818 478116 205824 478168
rect 205876 478156 205882 478168
rect 217318 478156 217324 478168
rect 205876 478128 217324 478156
rect 205876 478116 205882 478128
rect 217318 478116 217324 478128
rect 217376 478116 217382 478168
rect 233326 478116 233332 478168
rect 233384 478156 233390 478168
rect 366358 478156 366364 478168
rect 233384 478128 366364 478156
rect 233384 478116 233390 478128
rect 366358 478116 366364 478128
rect 366416 478116 366422 478168
rect 298002 478048 298008 478100
rect 298060 478088 298066 478100
rect 298278 478088 298284 478100
rect 298060 478060 298284 478088
rect 298060 478048 298066 478060
rect 298278 478048 298284 478060
rect 298336 478048 298342 478100
rect 60734 477912 60740 477964
rect 60792 477952 60798 477964
rect 61102 477952 61108 477964
rect 60792 477924 61108 477952
rect 60792 477912 60798 477924
rect 61102 477912 61108 477924
rect 61160 477912 61166 477964
rect 183646 477640 183652 477692
rect 183704 477680 183710 477692
rect 184014 477680 184020 477692
rect 183704 477652 184020 477680
rect 183704 477640 183710 477652
rect 184014 477640 184020 477652
rect 184072 477640 184078 477692
rect 185026 477640 185032 477692
rect 185084 477680 185090 477692
rect 185854 477680 185860 477692
rect 185084 477652 185860 477680
rect 185084 477640 185090 477652
rect 185854 477640 185860 477652
rect 185912 477640 185918 477692
rect 298186 477572 298192 477624
rect 298244 477612 298250 477624
rect 299014 477612 299020 477624
rect 298244 477584 299020 477612
rect 298244 477572 298250 477584
rect 299014 477572 299020 477584
rect 299072 477572 299078 477624
rect 59630 477436 59636 477488
rect 59688 477476 59694 477488
rect 135990 477476 135996 477488
rect 59688 477448 135996 477476
rect 59688 477436 59694 477448
rect 135990 477436 135996 477448
rect 136048 477436 136054 477488
rect 289262 477436 289268 477488
rect 289320 477476 289326 477488
rect 373810 477476 373816 477488
rect 289320 477448 373816 477476
rect 289320 477436 289326 477448
rect 373810 477436 373816 477448
rect 373868 477436 373874 477488
rect 45370 477368 45376 477420
rect 45428 477408 45434 477420
rect 123294 477408 123300 477420
rect 45428 477380 123300 477408
rect 45428 477368 45434 477380
rect 123294 477368 123300 477380
rect 123352 477368 123358 477420
rect 287330 477368 287336 477420
rect 287388 477408 287394 477420
rect 379330 477408 379336 477420
rect 287388 477380 379336 477408
rect 287388 477368 287394 477380
rect 379330 477368 379336 477380
rect 379388 477368 379394 477420
rect 57422 477300 57428 477352
rect 57480 477340 57486 477352
rect 135254 477340 135260 477352
rect 57480 477312 135260 477340
rect 57480 477300 57486 477312
rect 135254 477300 135260 477312
rect 135312 477300 135318 477352
rect 265158 477300 265164 477352
rect 265216 477340 265222 477352
rect 362586 477340 362592 477352
rect 265216 477312 362592 477340
rect 265216 477300 265222 477312
rect 362586 477300 362592 477312
rect 362644 477300 362650 477352
rect 55950 477232 55956 477284
rect 56008 477272 56014 477284
rect 133874 477272 133880 477284
rect 56008 477244 133880 477272
rect 56008 477232 56014 477244
rect 133874 477232 133880 477244
rect 133932 477232 133938 477284
rect 268102 477232 268108 477284
rect 268160 477272 268166 477284
rect 366266 477272 366272 477284
rect 268160 477244 366272 477272
rect 268160 477232 268166 477244
rect 366266 477232 366272 477244
rect 366324 477232 366330 477284
rect 54478 477164 54484 477216
rect 54536 477204 54542 477216
rect 133966 477204 133972 477216
rect 54536 477176 133972 477204
rect 54536 477164 54542 477176
rect 133966 477164 133972 477176
rect 134024 477164 134030 477216
rect 275646 477164 275652 477216
rect 275704 477204 275710 477216
rect 373718 477204 373724 477216
rect 275704 477176 373724 477204
rect 275704 477164 275710 477176
rect 373718 477164 373724 477176
rect 373776 477164 373782 477216
rect 50062 477096 50068 477148
rect 50120 477136 50126 477148
rect 131206 477136 131212 477148
rect 50120 477108 131212 477136
rect 50120 477096 50126 477108
rect 131206 477096 131212 477108
rect 131264 477096 131270 477148
rect 265066 477096 265072 477148
rect 265124 477136 265130 477148
rect 365438 477136 365444 477148
rect 265124 477108 365444 477136
rect 265124 477096 265130 477108
rect 365438 477096 365444 477108
rect 365496 477096 365502 477148
rect 49050 477028 49056 477080
rect 49108 477068 49114 477080
rect 130654 477068 130660 477080
rect 49108 477040 130660 477068
rect 49108 477028 49114 477040
rect 130654 477028 130660 477040
rect 130712 477028 130718 477080
rect 263686 477028 263692 477080
rect 263744 477068 263750 477080
rect 368106 477068 368112 477080
rect 263744 477040 368112 477068
rect 263744 477028 263750 477040
rect 368106 477028 368112 477040
rect 368164 477028 368170 477080
rect 48958 476960 48964 477012
rect 49016 477000 49022 477012
rect 132586 477000 132592 477012
rect 49016 476972 132592 477000
rect 49016 476960 49022 476972
rect 132586 476960 132592 476972
rect 132644 476960 132650 477012
rect 263778 476960 263784 477012
rect 263836 477000 263842 477012
rect 375006 477000 375012 477012
rect 263836 476972 375012 477000
rect 263836 476960 263842 476972
rect 375006 476960 375012 476972
rect 375064 476960 375070 477012
rect 46290 476892 46296 476944
rect 46348 476932 46354 476944
rect 132862 476932 132868 476944
rect 46348 476904 132868 476932
rect 46348 476892 46354 476904
rect 132862 476892 132868 476904
rect 132920 476892 132926 476944
rect 237374 476892 237380 476944
rect 237432 476932 237438 476944
rect 366450 476932 366456 476944
rect 237432 476904 366456 476932
rect 237432 476892 237438 476904
rect 366450 476892 366456 476904
rect 366508 476892 366514 476944
rect 42150 476824 42156 476876
rect 42208 476864 42214 476876
rect 131574 476864 131580 476876
rect 42208 476836 131580 476864
rect 42208 476824 42214 476836
rect 131574 476824 131580 476836
rect 131632 476824 131638 476876
rect 162946 476824 162952 476876
rect 163004 476864 163010 476876
rect 207658 476864 207664 476876
rect 163004 476836 207664 476864
rect 163004 476824 163010 476836
rect 207658 476824 207664 476836
rect 207716 476824 207722 476876
rect 236822 476824 236828 476876
rect 236880 476864 236886 476876
rect 365070 476864 365076 476876
rect 236880 476836 365076 476864
rect 236880 476824 236886 476836
rect 365070 476824 365076 476836
rect 365128 476824 365134 476876
rect 44726 476756 44732 476808
rect 44784 476796 44790 476808
rect 143626 476796 143632 476808
rect 44784 476768 143632 476796
rect 44784 476756 44790 476768
rect 143626 476756 143632 476768
rect 143684 476756 143690 476808
rect 165706 476756 165712 476808
rect 165764 476796 165770 476808
rect 218790 476796 218796 476808
rect 165764 476768 218796 476796
rect 165764 476756 165770 476768
rect 218790 476756 218796 476768
rect 218848 476756 218854 476808
rect 247034 476756 247040 476808
rect 247092 476796 247098 476808
rect 376294 476796 376300 476808
rect 247092 476768 376300 476796
rect 247092 476756 247098 476768
rect 376294 476756 376300 476768
rect 376352 476756 376358 476808
rect 58434 476688 58440 476740
rect 58492 476728 58498 476740
rect 128446 476728 128452 476740
rect 58492 476700 128452 476728
rect 58492 476688 58498 476700
rect 128446 476688 128452 476700
rect 128504 476688 128510 476740
rect 292758 476688 292764 476740
rect 292816 476728 292822 476740
rect 375742 476728 375748 476740
rect 292816 476700 375748 476728
rect 292816 476688 292822 476700
rect 375742 476688 375748 476700
rect 375800 476688 375806 476740
rect 59814 476620 59820 476672
rect 59872 476660 59878 476672
rect 127618 476660 127624 476672
rect 59872 476632 127624 476660
rect 59872 476620 59878 476632
rect 127618 476620 127624 476632
rect 127676 476620 127682 476672
rect 43990 476552 43996 476604
rect 44048 476592 44054 476604
rect 80974 476592 80980 476604
rect 44048 476564 80980 476592
rect 44048 476552 44054 476564
rect 80974 476552 80980 476564
rect 81032 476552 81038 476604
rect 100846 476484 100852 476536
rect 100904 476524 100910 476536
rect 101214 476524 101220 476536
rect 100904 476496 101220 476524
rect 100904 476484 100910 476496
rect 101214 476484 101220 476496
rect 101272 476484 101278 476536
rect 88426 476416 88432 476468
rect 88484 476456 88490 476468
rect 88886 476456 88892 476468
rect 88484 476428 88892 476456
rect 88484 476416 88490 476428
rect 88886 476416 88892 476428
rect 88944 476416 88950 476468
rect 292574 475736 292580 475788
rect 292632 475776 292638 475788
rect 376754 475776 376760 475788
rect 292632 475748 376760 475776
rect 292632 475736 292638 475748
rect 376754 475736 376760 475748
rect 376812 475736 376818 475788
rect 269114 475668 269120 475720
rect 269172 475708 269178 475720
rect 374362 475708 374368 475720
rect 269172 475680 374368 475708
rect 269172 475668 269178 475680
rect 374362 475668 374368 475680
rect 374420 475668 374426 475720
rect 258902 475600 258908 475652
rect 258960 475640 258966 475652
rect 372154 475640 372160 475652
rect 258960 475612 372160 475640
rect 258960 475600 258966 475612
rect 372154 475600 372160 475612
rect 372212 475600 372218 475652
rect 185026 475532 185032 475584
rect 185084 475572 185090 475584
rect 213178 475572 213184 475584
rect 185084 475544 213184 475572
rect 185084 475532 185090 475544
rect 213178 475532 213184 475544
rect 213236 475532 213242 475584
rect 254026 475532 254032 475584
rect 254084 475572 254090 475584
rect 379054 475572 379060 475584
rect 254084 475544 379060 475572
rect 254084 475532 254090 475544
rect 379054 475532 379060 475544
rect 379112 475532 379118 475584
rect 176746 475464 176752 475516
rect 176804 475504 176810 475516
rect 207842 475504 207848 475516
rect 176804 475476 207848 475504
rect 176804 475464 176810 475476
rect 207842 475464 207848 475476
rect 207900 475464 207906 475516
rect 245286 475464 245292 475516
rect 245344 475504 245350 475516
rect 370590 475504 370596 475516
rect 245344 475476 370596 475504
rect 245344 475464 245350 475476
rect 370590 475464 370596 475476
rect 370648 475464 370654 475516
rect 57606 475396 57612 475448
rect 57664 475436 57670 475448
rect 114738 475436 114744 475448
rect 57664 475408 114744 475436
rect 57664 475396 57670 475408
rect 114738 475396 114744 475408
rect 114796 475396 114802 475448
rect 164602 475396 164608 475448
rect 164660 475436 164666 475448
rect 211890 475436 211896 475448
rect 164660 475408 211896 475436
rect 164660 475396 164666 475408
rect 211890 475396 211896 475408
rect 211948 475396 211954 475448
rect 226610 475396 226616 475448
rect 226668 475436 226674 475448
rect 363598 475436 363604 475448
rect 226668 475408 363604 475436
rect 226668 475396 226674 475408
rect 363598 475396 363604 475408
rect 363656 475396 363662 475448
rect 60826 475328 60832 475380
rect 60884 475368 60890 475380
rect 199470 475368 199476 475380
rect 60884 475340 199476 475368
rect 60884 475328 60890 475340
rect 199470 475328 199476 475340
rect 199528 475328 199534 475380
rect 238754 475328 238760 475380
rect 238812 475368 238818 475380
rect 378870 475368 378876 475380
rect 238812 475340 378876 475368
rect 238812 475328 238818 475340
rect 378870 475328 378876 475340
rect 378928 475328 378934 475380
rect 291930 474648 291936 474700
rect 291988 474688 291994 474700
rect 368382 474688 368388 474700
rect 291988 474660 368388 474688
rect 291988 474648 291994 474660
rect 368382 474648 368388 474660
rect 368440 474648 368446 474700
rect 85666 474580 85672 474632
rect 85724 474620 85730 474632
rect 85850 474620 85856 474632
rect 85724 474592 85856 474620
rect 85724 474580 85730 474592
rect 85850 474580 85856 474592
rect 85908 474580 85914 474632
rect 273438 474580 273444 474632
rect 273496 474620 273502 474632
rect 361482 474620 361488 474632
rect 273496 474592 361488 474620
rect 273496 474580 273502 474592
rect 361482 474580 361488 474592
rect 361540 474580 361546 474632
rect 280430 474512 280436 474564
rect 280488 474552 280494 474564
rect 369670 474552 369676 474564
rect 280488 474524 369676 474552
rect 280488 474512 280494 474524
rect 369670 474512 369676 474524
rect 369728 474512 369734 474564
rect 278222 474444 278228 474496
rect 278280 474484 278286 474496
rect 368290 474484 368296 474496
rect 278280 474456 368296 474484
rect 278280 474444 278286 474456
rect 368290 474444 368296 474456
rect 368348 474444 368354 474496
rect 257614 474376 257620 474428
rect 257672 474416 257678 474428
rect 362678 474416 362684 474428
rect 257672 474388 362684 474416
rect 257672 474376 257678 474388
rect 362678 474376 362684 474388
rect 362736 474376 362742 474428
rect 176654 474308 176660 474360
rect 176712 474348 176718 474360
rect 209222 474348 209228 474360
rect 176712 474320 209228 474348
rect 176712 474308 176718 474320
rect 209222 474308 209228 474320
rect 209280 474308 209286 474360
rect 262582 474308 262588 474360
rect 262640 474348 262646 474360
rect 373534 474348 373540 474360
rect 262640 474320 373540 474348
rect 262640 474308 262646 474320
rect 373534 474308 373540 474320
rect 373592 474308 373598 474360
rect 179782 474240 179788 474292
rect 179840 474280 179846 474292
rect 216122 474280 216128 474292
rect 179840 474252 216128 474280
rect 179840 474240 179846 474252
rect 216122 474240 216128 474252
rect 216180 474240 216186 474292
rect 259454 474240 259460 474292
rect 259512 474280 259518 474292
rect 373626 474280 373632 474292
rect 259512 474252 373632 474280
rect 259512 474240 259518 474252
rect 373626 474240 373632 474252
rect 373684 474240 373690 474292
rect 159358 474172 159364 474224
rect 159416 474212 159422 474224
rect 218882 474212 218888 474224
rect 159416 474184 218888 474212
rect 159416 474172 159422 474184
rect 218882 474172 218888 474184
rect 218940 474172 218946 474224
rect 241606 474172 241612 474224
rect 241664 474212 241670 474224
rect 361022 474212 361028 474224
rect 241664 474184 361028 474212
rect 241664 474172 241670 474184
rect 361022 474172 361028 474184
rect 361080 474172 361086 474224
rect 51626 474104 51632 474156
rect 51684 474144 51690 474156
rect 99558 474144 99564 474156
rect 51684 474116 99564 474144
rect 51684 474104 51690 474116
rect 99558 474104 99564 474116
rect 99616 474104 99622 474156
rect 139486 474104 139492 474156
rect 139544 474144 139550 474156
rect 205818 474144 205824 474156
rect 139544 474116 205824 474144
rect 139544 474104 139550 474116
rect 205818 474104 205824 474116
rect 205876 474104 205882 474156
rect 244274 474104 244280 474156
rect 244332 474144 244338 474156
rect 371970 474144 371976 474156
rect 244332 474116 371976 474144
rect 244332 474104 244338 474116
rect 371970 474104 371976 474116
rect 372028 474104 372034 474156
rect 57790 474036 57796 474088
rect 57848 474076 57854 474088
rect 113266 474076 113272 474088
rect 57848 474048 113272 474076
rect 57848 474036 57854 474048
rect 113266 474036 113272 474048
rect 113324 474036 113330 474088
rect 126974 474036 126980 474088
rect 127032 474076 127038 474088
rect 201494 474076 201500 474088
rect 127032 474048 201500 474076
rect 127032 474036 127038 474048
rect 201494 474036 201500 474048
rect 201552 474036 201558 474088
rect 207198 474036 207204 474088
rect 207256 474076 207262 474088
rect 217226 474076 217232 474088
rect 207256 474048 217232 474076
rect 207256 474036 207262 474048
rect 217226 474036 217232 474048
rect 217284 474036 217290 474088
rect 229830 474036 229836 474088
rect 229888 474076 229894 474088
rect 363782 474076 363788 474088
rect 229888 474048 363788 474076
rect 229888 474036 229894 474048
rect 363782 474036 363788 474048
rect 363840 474036 363846 474088
rect 59354 473968 59360 474020
rect 59412 474008 59418 474020
rect 180150 474008 180156 474020
rect 59412 473980 180156 474008
rect 59412 473968 59418 473980
rect 180150 473968 180156 473980
rect 180208 473968 180214 474020
rect 186406 473968 186412 474020
rect 186464 474008 186470 474020
rect 212074 474008 212080 474020
rect 186464 473980 212080 474008
rect 186464 473968 186470 473980
rect 212074 473968 212080 473980
rect 212132 473968 212138 474020
rect 229186 473968 229192 474020
rect 229244 474008 229250 474020
rect 363690 474008 363696 474020
rect 229244 473980 363696 474008
rect 229244 473968 229250 473980
rect 363690 473968 363696 473980
rect 363748 473968 363754 474020
rect 290182 473900 290188 473952
rect 290240 473940 290246 473952
rect 357158 473940 357164 473952
rect 290240 473912 357164 473940
rect 290240 473900 290246 473912
rect 357158 473900 357164 473912
rect 357216 473900 357222 473952
rect 289814 473016 289820 473068
rect 289872 473056 289878 473068
rect 360746 473056 360752 473068
rect 289872 473028 360752 473056
rect 289872 473016 289878 473028
rect 360746 473016 360752 473028
rect 360804 473016 360810 473068
rect 294046 472948 294052 473000
rect 294104 472988 294110 473000
rect 369762 472988 369768 473000
rect 294104 472960 369768 472988
rect 294104 472948 294110 472960
rect 369762 472948 369768 472960
rect 369820 472948 369826 473000
rect 273346 472880 273352 472932
rect 273404 472920 273410 472932
rect 362862 472920 362868 472932
rect 273404 472892 362868 472920
rect 273404 472880 273410 472892
rect 362862 472880 362868 472892
rect 362920 472880 362926 472932
rect 262306 472812 262312 472864
rect 262364 472852 262370 472864
rect 370774 472852 370780 472864
rect 262364 472824 370780 472852
rect 262364 472812 262370 472824
rect 370774 472812 370780 472824
rect 370832 472812 370838 472864
rect 188062 472744 188068 472796
rect 188120 472784 188126 472796
rect 210694 472784 210700 472796
rect 188120 472756 210700 472784
rect 188120 472744 188126 472756
rect 210694 472744 210700 472756
rect 210752 472744 210758 472796
rect 263594 472744 263600 472796
rect 263652 472784 263658 472796
rect 372246 472784 372252 472796
rect 263652 472756 372252 472784
rect 263652 472744 263658 472756
rect 372246 472744 372252 472756
rect 372304 472744 372310 472796
rect 175366 472676 175372 472728
rect 175424 472716 175430 472728
rect 202138 472716 202144 472728
rect 175424 472688 202144 472716
rect 175424 472676 175430 472688
rect 202138 472676 202144 472688
rect 202196 472676 202202 472728
rect 226426 472676 226432 472728
rect 226484 472716 226490 472728
rect 367738 472716 367744 472728
rect 226484 472688 367744 472716
rect 226484 472676 226490 472688
rect 367738 472676 367744 472688
rect 367796 472676 367802 472728
rect 58618 472608 58624 472660
rect 58676 472648 58682 472660
rect 110598 472648 110604 472660
rect 58676 472620 110604 472648
rect 58676 472608 58682 472620
rect 110598 472608 110604 472620
rect 110656 472608 110662 472660
rect 184934 472608 184940 472660
rect 184992 472648 184998 472660
rect 212166 472648 212172 472660
rect 184992 472620 212172 472648
rect 184992 472608 184998 472620
rect 212166 472608 212172 472620
rect 212224 472608 212230 472660
rect 227714 472608 227720 472660
rect 227772 472648 227778 472660
rect 374638 472648 374644 472660
rect 227772 472620 374644 472648
rect 227772 472608 227778 472620
rect 374638 472608 374644 472620
rect 374696 472608 374702 472660
rect 46198 471928 46204 471980
rect 46256 471968 46262 471980
rect 64874 471968 64880 471980
rect 46256 471940 64880 471968
rect 46256 471928 46262 471940
rect 64874 471928 64880 471940
rect 64932 471928 64938 471980
rect 192754 471928 192760 471980
rect 192812 471968 192818 471980
rect 213454 471968 213460 471980
rect 192812 471940 213460 471968
rect 192812 471928 192818 471940
rect 213454 471928 213460 471940
rect 213512 471928 213518 471980
rect 296254 471928 296260 471980
rect 296312 471968 296318 471980
rect 362034 471968 362040 471980
rect 296312 471940 362040 471968
rect 296312 471928 296318 471940
rect 362034 471928 362040 471940
rect 362092 471928 362098 471980
rect 50982 471860 50988 471912
rect 51040 471900 51046 471912
rect 82814 471900 82820 471912
rect 51040 471872 82820 471900
rect 51040 471860 51046 471872
rect 82814 471860 82820 471872
rect 82872 471860 82878 471912
rect 183094 471860 183100 471912
rect 183152 471900 183158 471912
rect 205082 471900 205088 471912
rect 183152 471872 205088 471900
rect 183152 471860 183158 471872
rect 205082 471860 205088 471872
rect 205140 471860 205146 471912
rect 287146 471860 287152 471912
rect 287204 471900 287210 471912
rect 358722 471900 358728 471912
rect 287204 471872 358728 471900
rect 287204 471860 287210 471872
rect 358722 471860 358728 471872
rect 358780 471860 358786 471912
rect 51534 471792 51540 471844
rect 51592 471832 51598 471844
rect 84470 471832 84476 471844
rect 51592 471804 84476 471832
rect 51592 471792 51598 471804
rect 84470 471792 84476 471804
rect 84528 471792 84534 471844
rect 192018 471792 192024 471844
rect 192076 471832 192082 471844
rect 217686 471832 217692 471844
rect 192076 471804 217692 471832
rect 192076 471792 192082 471804
rect 217686 471792 217692 471804
rect 217744 471792 217750 471844
rect 298186 471792 298192 471844
rect 298244 471832 298250 471844
rect 372430 471832 372436 471844
rect 298244 471804 372436 471832
rect 298244 471792 298250 471804
rect 372430 471792 372436 471804
rect 372488 471792 372494 471844
rect 50614 471724 50620 471776
rect 50672 471764 50678 471776
rect 82906 471764 82912 471776
rect 50672 471736 82912 471764
rect 50672 471724 50678 471736
rect 82906 471724 82912 471736
rect 82964 471724 82970 471776
rect 190638 471724 190644 471776
rect 190696 471764 190702 471776
rect 216398 471764 216404 471776
rect 190696 471736 216404 471764
rect 190696 471724 190702 471736
rect 216398 471724 216404 471736
rect 216456 471724 216462 471776
rect 298094 471724 298100 471776
rect 298152 471764 298158 471776
rect 372614 471764 372620 471776
rect 298152 471736 372620 471764
rect 298152 471724 298158 471736
rect 372614 471724 372620 471736
rect 372672 471724 372678 471776
rect 49418 471656 49424 471708
rect 49476 471696 49482 471708
rect 83182 471696 83188 471708
rect 49476 471668 83188 471696
rect 49476 471656 49482 471668
rect 83182 471656 83188 471668
rect 83240 471656 83246 471708
rect 190546 471656 190552 471708
rect 190604 471696 190610 471708
rect 217502 471696 217508 471708
rect 190604 471668 217508 471696
rect 190604 471656 190610 471668
rect 217502 471656 217508 471668
rect 217560 471656 217566 471708
rect 298278 471656 298284 471708
rect 298336 471696 298342 471708
rect 375190 471696 375196 471708
rect 298336 471668 375196 471696
rect 298336 471656 298342 471668
rect 375190 471656 375196 471668
rect 375248 471656 375254 471708
rect 54662 471588 54668 471640
rect 54720 471628 54726 471640
rect 100754 471628 100760 471640
rect 54720 471600 100760 471628
rect 54720 471588 54726 471600
rect 100754 471588 100760 471600
rect 100812 471588 100818 471640
rect 183646 471588 183652 471640
rect 183704 471628 183710 471640
rect 210786 471628 210792 471640
rect 183704 471600 210792 471628
rect 183704 471588 183710 471600
rect 210786 471588 210792 471600
rect 210844 471588 210850 471640
rect 297726 471588 297732 471640
rect 297784 471628 297790 471640
rect 375098 471628 375104 471640
rect 297784 471600 375104 471628
rect 297784 471588 297790 471600
rect 375098 471588 375104 471600
rect 375156 471588 375162 471640
rect 57330 471520 57336 471572
rect 57388 471560 57394 471572
rect 103606 471560 103612 471572
rect 57388 471532 103612 471560
rect 57388 471520 57394 471532
rect 103606 471520 103612 471532
rect 103664 471520 103670 471572
rect 161566 471520 161572 471572
rect 161624 471560 161630 471572
rect 214650 471560 214656 471572
rect 161624 471532 214656 471560
rect 161624 471520 161630 471532
rect 214650 471520 214656 471532
rect 214708 471520 214714 471572
rect 288526 471520 288532 471572
rect 288584 471560 288590 471572
rect 371142 471560 371148 471572
rect 288584 471532 371148 471560
rect 288584 471520 288590 471532
rect 371142 471520 371148 471532
rect 371200 471520 371206 471572
rect 53282 471452 53288 471504
rect 53340 471492 53346 471504
rect 100846 471492 100852 471504
rect 53340 471464 100852 471492
rect 53340 471452 53346 471464
rect 100846 471452 100852 471464
rect 100904 471452 100910 471504
rect 140958 471452 140964 471504
rect 141016 471492 141022 471504
rect 200390 471492 200396 471504
rect 141016 471464 200396 471492
rect 141016 471452 141022 471464
rect 200390 471452 200396 471464
rect 200448 471452 200454 471504
rect 276934 471452 276940 471504
rect 276992 471492 276998 471504
rect 358630 471492 358636 471504
rect 276992 471464 358636 471492
rect 276992 471452 276998 471464
rect 358630 471452 358636 471464
rect 358688 471452 358694 471504
rect 53190 471384 53196 471436
rect 53248 471424 53254 471436
rect 100938 471424 100944 471436
rect 53248 471396 100944 471424
rect 53248 471384 53254 471396
rect 100938 471384 100944 471396
rect 100996 471384 101002 471436
rect 140866 471384 140872 471436
rect 140924 471424 140930 471436
rect 203150 471424 203156 471436
rect 140924 471396 203156 471424
rect 140924 471384 140930 471396
rect 203150 471384 203156 471396
rect 203208 471384 203214 471436
rect 285858 471384 285864 471436
rect 285916 471424 285922 471436
rect 376478 471424 376484 471436
rect 285916 471396 376484 471424
rect 285916 471384 285922 471396
rect 376478 471384 376484 471396
rect 376536 471384 376542 471436
rect 50246 471316 50252 471368
rect 50304 471356 50310 471368
rect 98638 471356 98644 471368
rect 50304 471328 98644 471356
rect 50304 471316 50310 471328
rect 98638 471316 98644 471328
rect 98696 471316 98702 471368
rect 140774 471316 140780 471368
rect 140832 471356 140838 471368
rect 205910 471356 205916 471368
rect 140832 471328 205916 471356
rect 140832 471316 140838 471328
rect 205910 471316 205916 471328
rect 205968 471316 205974 471368
rect 240134 471316 240140 471368
rect 240192 471356 240198 471368
rect 362402 471356 362408 471368
rect 240192 471328 362408 471356
rect 240192 471316 240198 471328
rect 362402 471316 362408 471328
rect 362460 471316 362466 471368
rect 57698 471248 57704 471300
rect 57756 471288 57762 471300
rect 113358 471288 113364 471300
rect 57756 471260 113364 471288
rect 57756 471248 57762 471260
rect 113358 471248 113364 471260
rect 113416 471248 113422 471300
rect 125686 471248 125692 471300
rect 125744 471288 125750 471300
rect 196894 471288 196900 471300
rect 125744 471260 196900 471288
rect 125744 471248 125750 471260
rect 196894 471248 196900 471260
rect 196952 471248 196958 471300
rect 240226 471248 240232 471300
rect 240284 471288 240290 471300
rect 363966 471288 363972 471300
rect 240284 471260 363972 471288
rect 240284 471248 240290 471260
rect 363966 471248 363972 471260
rect 364024 471248 364030 471300
rect 47394 471180 47400 471232
rect 47452 471220 47458 471232
rect 65518 471220 65524 471232
rect 47452 471192 65524 471220
rect 47452 471180 47458 471192
rect 65518 471180 65524 471192
rect 65576 471180 65582 471232
rect 183554 471180 183560 471232
rect 183612 471220 183618 471232
rect 203794 471220 203800 471232
rect 183612 471192 203800 471220
rect 183612 471180 183618 471192
rect 203794 471180 203800 471192
rect 203852 471180 203858 471232
rect 47486 471112 47492 471164
rect 47544 471152 47550 471164
rect 64966 471152 64972 471164
rect 47544 471124 64972 471152
rect 47544 471112 47550 471124
rect 64966 471112 64972 471124
rect 65024 471112 65030 471164
rect 182358 471112 182364 471164
rect 182416 471152 182422 471164
rect 202414 471152 202420 471164
rect 182416 471124 202420 471152
rect 182416 471112 182422 471124
rect 202414 471112 202420 471124
rect 202472 471112 202478 471164
rect 52086 471044 52092 471096
rect 52144 471084 52150 471096
rect 68278 471084 68284 471096
rect 52144 471056 68284 471084
rect 52144 471044 52150 471056
rect 68278 471044 68284 471056
rect 68336 471044 68342 471096
rect 183738 471044 183744 471096
rect 183796 471084 183802 471096
rect 200850 471084 200856 471096
rect 183796 471056 200856 471084
rect 183796 471044 183802 471056
rect 200850 471044 200856 471056
rect 200908 471044 200914 471096
rect 282914 470432 282920 470484
rect 282972 470472 282978 470484
rect 358078 470472 358084 470484
rect 282972 470444 358084 470472
rect 282972 470432 282978 470444
rect 358078 470432 358084 470444
rect 358136 470432 358142 470484
rect 283098 470364 283104 470416
rect 283156 470404 283162 470416
rect 359918 470404 359924 470416
rect 283156 470376 359924 470404
rect 283156 470364 283162 470376
rect 359918 470364 359924 470376
rect 359976 470364 359982 470416
rect 283006 470296 283012 470348
rect 283064 470336 283070 470348
rect 359826 470336 359832 470348
rect 283064 470308 359832 470336
rect 283064 470296 283070 470308
rect 359826 470296 359832 470308
rect 359884 470296 359890 470348
rect 285674 470228 285680 470280
rect 285732 470268 285738 470280
rect 364242 470268 364248 470280
rect 285732 470240 364248 470268
rect 285732 470228 285738 470240
rect 364242 470228 364248 470240
rect 364300 470228 364306 470280
rect 287054 470160 287060 470212
rect 287112 470200 287118 470212
rect 367646 470200 367652 470212
rect 287112 470172 367652 470200
rect 287112 470160 287118 470172
rect 367646 470160 367652 470172
rect 367704 470160 367710 470212
rect 285766 470092 285772 470144
rect 285824 470132 285830 470144
rect 377674 470132 377680 470144
rect 285824 470104 377680 470132
rect 285824 470092 285830 470104
rect 377674 470092 377680 470104
rect 377732 470092 377738 470144
rect 178126 470024 178132 470076
rect 178184 470064 178190 470076
rect 202322 470064 202328 470076
rect 178184 470036 202328 470064
rect 178184 470024 178190 470036
rect 202322 470024 202328 470036
rect 202380 470024 202386 470076
rect 284294 470024 284300 470076
rect 284352 470064 284358 470076
rect 377398 470064 377404 470076
rect 284352 470036 377404 470064
rect 284352 470024 284358 470036
rect 377398 470024 377404 470036
rect 377456 470024 377462 470076
rect 179506 469956 179512 470008
rect 179564 469996 179570 470008
rect 206462 469996 206468 470008
rect 179564 469968 206468 469996
rect 179564 469956 179570 469968
rect 206462 469956 206468 469968
rect 206520 469956 206526 470008
rect 284386 469956 284392 470008
rect 284444 469996 284450 470008
rect 377582 469996 377588 470008
rect 284444 469968 377588 469996
rect 284444 469956 284450 469968
rect 377582 469956 377588 469968
rect 377640 469956 377646 470008
rect 50798 469888 50804 469940
rect 50856 469928 50862 469940
rect 81618 469928 81624 469940
rect 50856 469900 81624 469928
rect 50856 469888 50862 469900
rect 81618 469888 81624 469900
rect 81676 469888 81682 469940
rect 164234 469888 164240 469940
rect 164292 469928 164298 469940
rect 218974 469928 218980 469940
rect 164292 469900 218980 469928
rect 164292 469888 164298 469900
rect 218974 469888 218980 469900
rect 219032 469888 219038 469940
rect 281534 469888 281540 469940
rect 281592 469928 281598 469940
rect 376570 469928 376576 469940
rect 281592 469900 376576 469928
rect 281592 469888 281598 469900
rect 376570 469888 376576 469900
rect 376628 469888 376634 469940
rect 57514 469820 57520 469872
rect 57572 469860 57578 469872
rect 111978 469860 111984 469872
rect 57572 469832 111984 469860
rect 57572 469820 57578 469832
rect 111978 469820 111984 469832
rect 112036 469820 112042 469872
rect 143534 469820 143540 469872
rect 143592 469860 143598 469872
rect 210418 469860 210424 469872
rect 143592 469832 210424 469860
rect 143592 469820 143598 469832
rect 210418 469820 210424 469832
rect 210476 469820 210482 469872
rect 281626 469820 281632 469872
rect 281684 469860 281690 469872
rect 379974 469860 379980 469872
rect 281684 469832 379980 469860
rect 281684 469820 281690 469832
rect 379974 469820 379980 469832
rect 380032 469820 380038 469872
rect 49510 469140 49516 469192
rect 49568 469180 49574 469192
rect 80054 469180 80060 469192
rect 49568 469152 80060 469180
rect 49568 469140 49574 469152
rect 80054 469140 80060 469152
rect 80112 469140 80118 469192
rect 193398 469140 193404 469192
rect 193456 469180 193462 469192
rect 216490 469180 216496 469192
rect 193456 469152 216496 469180
rect 193456 469140 193462 469152
rect 216490 469140 216496 469152
rect 216548 469140 216554 469192
rect 273254 469140 273260 469192
rect 273312 469180 273318 469192
rect 363414 469180 363420 469192
rect 273312 469152 363420 469180
rect 273312 469140 273318 469152
rect 363414 469140 363420 469152
rect 363472 469140 363478 469192
rect 50706 469072 50712 469124
rect 50764 469112 50770 469124
rect 78766 469112 78772 469124
rect 50764 469084 78772 469112
rect 50764 469072 50770 469084
rect 78766 469072 78772 469084
rect 78824 469072 78830 469124
rect 178034 469072 178040 469124
rect 178092 469112 178098 469124
rect 210878 469112 210884 469124
rect 178092 469084 210884 469112
rect 178092 469072 178098 469084
rect 210878 469072 210884 469084
rect 210936 469072 210942 469124
rect 266538 469072 266544 469124
rect 266596 469112 266602 469124
rect 359550 469112 359556 469124
rect 266596 469084 359556 469112
rect 266596 469072 266602 469084
rect 359550 469072 359556 469084
rect 359608 469072 359614 469124
rect 46014 469004 46020 469056
rect 46072 469044 46078 469056
rect 63586 469044 63592 469056
rect 46072 469016 63592 469044
rect 46072 469004 46078 469016
rect 63586 469004 63592 469016
rect 63644 469004 63650 469056
rect 168558 469004 168564 469056
rect 168616 469044 168622 469056
rect 202230 469044 202236 469056
rect 168616 469016 202236 469044
rect 168616 469004 168622 469016
rect 202230 469004 202236 469016
rect 202288 469004 202294 469056
rect 266446 469004 266452 469056
rect 266504 469044 266510 469056
rect 359642 469044 359648 469056
rect 266504 469016 359648 469044
rect 266504 469004 266510 469016
rect 359642 469004 359648 469016
rect 359700 469004 359706 469056
rect 48774 468936 48780 468988
rect 48832 468976 48838 468988
rect 70578 468976 70584 468988
rect 48832 468948 70584 468976
rect 48832 468936 48838 468948
rect 70578 468936 70584 468948
rect 70636 468936 70642 468988
rect 167086 468936 167092 468988
rect 167144 468976 167150 468988
rect 209130 468976 209136 468988
rect 167144 468948 209136 468976
rect 167144 468936 167150 468948
rect 209130 468936 209136 468948
rect 209188 468936 209194 468988
rect 266354 468936 266360 468988
rect 266412 468976 266418 468988
rect 361298 468976 361304 468988
rect 266412 468948 361304 468976
rect 266412 468936 266418 468948
rect 361298 468936 361304 468948
rect 361356 468936 361362 468988
rect 56134 468868 56140 468920
rect 56192 468908 56198 468920
rect 85574 468908 85580 468920
rect 56192 468880 85580 468908
rect 56192 468868 56198 468880
rect 85574 468868 85580 468880
rect 85632 468868 85638 468920
rect 167178 468868 167184 468920
rect 167236 468908 167242 468920
rect 210602 468908 210608 468920
rect 167236 468880 210608 468908
rect 167236 468868 167242 468880
rect 210602 468868 210608 468880
rect 210660 468868 210666 468920
rect 272058 468868 272064 468920
rect 272116 468908 272122 468920
rect 369026 468908 369032 468920
rect 272116 468880 369032 468908
rect 272116 468868 272122 468880
rect 369026 468868 369032 468880
rect 369084 468868 369090 468920
rect 56226 468800 56232 468852
rect 56284 468840 56290 468852
rect 87138 468840 87144 468852
rect 56284 468812 87144 468840
rect 56284 468800 56290 468812
rect 87138 468800 87144 468812
rect 87196 468800 87202 468852
rect 168466 468800 168472 468852
rect 168524 468840 168530 468852
rect 214742 468840 214748 468852
rect 168524 468812 214748 468840
rect 168524 468800 168530 468812
rect 214742 468800 214748 468812
rect 214800 468800 214806 468852
rect 264974 468800 264980 468852
rect 265032 468840 265038 468852
rect 364058 468840 364064 468852
rect 265032 468812 364064 468840
rect 265032 468800 265038 468812
rect 364058 468800 364064 468812
rect 364116 468800 364122 468852
rect 54938 468732 54944 468784
rect 54996 468772 55002 468784
rect 86954 468772 86960 468784
rect 54996 468744 86960 468772
rect 54996 468732 55002 468744
rect 86954 468732 86960 468744
rect 87012 468732 87018 468784
rect 139394 468732 139400 468784
rect 139452 468772 139458 468784
rect 196986 468772 196992 468784
rect 139452 468744 196992 468772
rect 139452 468732 139458 468744
rect 196986 468732 196992 468744
rect 197044 468732 197050 468784
rect 255314 468732 255320 468784
rect 255372 468772 255378 468784
rect 361206 468772 361212 468784
rect 255372 468744 361212 468772
rect 255372 468732 255378 468744
rect 361206 468732 361212 468744
rect 361264 468732 361270 468784
rect 53374 468664 53380 468716
rect 53432 468704 53438 468716
rect 85666 468704 85672 468716
rect 53432 468676 85672 468704
rect 53432 468664 53438 468676
rect 85666 468664 85672 468676
rect 85724 468664 85730 468716
rect 142338 468664 142344 468716
rect 142396 468704 142402 468716
rect 200482 468704 200488 468716
rect 142396 468676 200488 468704
rect 142396 468664 142402 468676
rect 200482 468664 200488 468676
rect 200540 468664 200546 468716
rect 267734 468664 267740 468716
rect 267792 468704 267798 468716
rect 377306 468704 377312 468716
rect 267792 468676 377312 468704
rect 267792 468664 267798 468676
rect 377306 468664 377312 468676
rect 377364 468664 377370 468716
rect 59906 468596 59912 468648
rect 59964 468636 59970 468648
rect 92566 468636 92572 468648
rect 59964 468608 92572 468636
rect 59964 468596 59970 468608
rect 92566 468596 92572 468608
rect 92624 468596 92630 468648
rect 109034 468596 109040 468648
rect 109092 468636 109098 468648
rect 197722 468636 197728 468648
rect 109092 468608 197728 468636
rect 109092 468596 109098 468608
rect 197722 468596 197728 468608
rect 197780 468596 197786 468648
rect 249978 468596 249984 468648
rect 250036 468636 250042 468648
rect 365162 468636 365168 468648
rect 250036 468608 365168 468636
rect 250036 468596 250042 468608
rect 365162 468596 365168 468608
rect 365220 468596 365226 468648
rect 53466 468528 53472 468580
rect 53524 468568 53530 468580
rect 87046 468568 87052 468580
rect 53524 468540 87052 468568
rect 53524 468528 53530 468540
rect 87046 468528 87052 468540
rect 87104 468528 87110 468580
rect 107838 468528 107844 468580
rect 107896 468568 107902 468580
rect 198918 468568 198924 468580
rect 107896 468540 198924 468568
rect 107896 468528 107902 468540
rect 198918 468528 198924 468540
rect 198976 468528 198982 468580
rect 251358 468528 251364 468580
rect 251416 468568 251422 468580
rect 369302 468568 369308 468580
rect 251416 468540 369308 468568
rect 251416 468528 251422 468540
rect 369302 468528 369308 468540
rect 369360 468528 369366 468580
rect 49326 468460 49332 468512
rect 49384 468500 49390 468512
rect 93946 468500 93952 468512
rect 49384 468472 93952 468500
rect 49384 468460 49390 468472
rect 93946 468460 93952 468472
rect 94004 468460 94010 468512
rect 107746 468460 107752 468512
rect 107804 468500 107810 468512
rect 203058 468500 203064 468512
rect 107804 468472 203064 468500
rect 107804 468460 107810 468472
rect 203058 468460 203064 468472
rect 203116 468460 203122 468512
rect 252554 468460 252560 468512
rect 252612 468500 252618 468512
rect 376202 468500 376208 468512
rect 252612 468472 376208 468500
rect 252612 468460 252618 468472
rect 376202 468460 376208 468472
rect 376260 468460 376266 468512
rect 191926 468392 191932 468444
rect 191984 468432 191990 468444
rect 214374 468432 214380 468444
rect 191984 468404 214380 468432
rect 191984 468392 191990 468404
rect 214374 468392 214380 468404
rect 214432 468392 214438 468444
rect 280154 468392 280160 468444
rect 280212 468432 280218 468444
rect 363506 468432 363512 468444
rect 280212 468404 363512 468432
rect 280212 468392 280218 468404
rect 363506 468392 363512 468404
rect 363564 468392 363570 468444
rect 191834 468324 191840 468376
rect 191892 468364 191898 468376
rect 211522 468364 211528 468376
rect 191892 468336 211528 468364
rect 191892 468324 191898 468336
rect 211522 468324 211528 468336
rect 211580 468324 211586 468376
rect 189166 468256 189172 468308
rect 189224 468296 189230 468308
rect 208026 468296 208032 468308
rect 189224 468268 208032 468296
rect 189224 468256 189230 468268
rect 208026 468256 208032 468268
rect 208084 468256 208090 468308
rect 45094 467780 45100 467832
rect 45152 467820 45158 467832
rect 73798 467820 73804 467832
rect 45152 467792 73804 467820
rect 45152 467780 45158 467792
rect 73798 467780 73804 467792
rect 73856 467780 73862 467832
rect 80698 467780 80704 467832
rect 80756 467820 80762 467832
rect 178034 467820 178040 467832
rect 80756 467792 178040 467820
rect 80756 467780 80762 467792
rect 178034 467780 178040 467792
rect 178092 467780 178098 467832
rect 293954 467780 293960 467832
rect 294012 467820 294018 467832
rect 357986 467820 357992 467832
rect 294012 467792 357992 467820
rect 294012 467780 294018 467792
rect 357986 467780 357992 467792
rect 358044 467780 358050 467832
rect 44818 467712 44824 467764
rect 44876 467752 44882 467764
rect 73982 467752 73988 467764
rect 44876 467724 73988 467752
rect 44876 467712 44882 467724
rect 73982 467712 73988 467724
rect 74040 467712 74046 467764
rect 291286 467712 291292 467764
rect 291344 467752 291350 467764
rect 362126 467752 362132 467764
rect 291344 467724 362132 467752
rect 291344 467712 291350 467724
rect 362126 467712 362132 467724
rect 362184 467712 362190 467764
rect 42518 467644 42524 467696
rect 42576 467684 42582 467696
rect 73890 467684 73896 467696
rect 42576 467656 73896 467684
rect 42576 467644 42582 467656
rect 73890 467644 73896 467656
rect 73948 467644 73954 467696
rect 288434 467644 288440 467696
rect 288492 467684 288498 467696
rect 364794 467684 364800 467696
rect 288492 467656 364800 467684
rect 288492 467644 288498 467656
rect 364794 467644 364800 467656
rect 364852 467644 364858 467696
rect 53098 467576 53104 467628
rect 53156 467616 53162 467628
rect 99650 467616 99656 467628
rect 53156 467588 99656 467616
rect 53156 467576 53162 467588
rect 99650 467576 99656 467588
rect 99708 467576 99714 467628
rect 277486 467576 277492 467628
rect 277544 467616 277550 467628
rect 370222 467616 370228 467628
rect 277544 467588 370228 467616
rect 277544 467576 277550 467588
rect 370222 467576 370228 467588
rect 370280 467576 370286 467628
rect 52362 467508 52368 467560
rect 52420 467548 52426 467560
rect 99466 467548 99472 467560
rect 52420 467520 99472 467548
rect 52420 467508 52426 467520
rect 99466 467508 99472 467520
rect 99524 467508 99530 467560
rect 274634 467508 274640 467560
rect 274692 467548 274698 467560
rect 367554 467548 367560 467560
rect 274692 467520 367560 467548
rect 274692 467508 274698 467520
rect 367554 467508 367560 467520
rect 367612 467508 367618 467560
rect 43898 467440 43904 467492
rect 43956 467480 43962 467492
rect 93854 467480 93860 467492
rect 43956 467452 93860 467480
rect 43956 467440 43962 467452
rect 93854 467440 93860 467452
rect 93912 467440 93918 467492
rect 256694 467440 256700 467492
rect 256752 467480 256758 467492
rect 361114 467480 361120 467492
rect 256752 467452 361120 467480
rect 256752 467440 256758 467452
rect 361114 467440 361120 467452
rect 361172 467440 361178 467492
rect 45002 467372 45008 467424
rect 45060 467412 45066 467424
rect 105078 467412 105084 467424
rect 45060 467384 105084 467412
rect 45060 467372 45066 467384
rect 105078 467372 105084 467384
rect 105136 467372 105142 467424
rect 182174 467372 182180 467424
rect 182232 467412 182238 467424
rect 212258 467412 212264 467424
rect 182232 467384 212264 467412
rect 182232 467372 182238 467384
rect 212258 467372 212264 467384
rect 212316 467372 212322 467424
rect 258166 467372 258172 467424
rect 258224 467412 258230 467424
rect 368198 467412 368204 467424
rect 258224 467384 368204 467412
rect 258224 467372 258230 467384
rect 368198 467372 368204 467384
rect 368256 467372 368262 467424
rect 43438 467304 43444 467356
rect 43496 467344 43502 467356
rect 103698 467344 103704 467356
rect 43496 467316 103704 467344
rect 43496 467304 43502 467316
rect 103698 467304 103704 467316
rect 103756 467304 103762 467356
rect 175274 467304 175280 467356
rect 175332 467344 175338 467356
rect 206554 467344 206560 467356
rect 175332 467316 206560 467344
rect 175332 467304 175338 467316
rect 206554 467304 206560 467316
rect 206612 467304 206618 467356
rect 251266 467304 251272 467356
rect 251324 467344 251330 467356
rect 365254 467344 365260 467356
rect 251324 467316 365260 467344
rect 251324 467304 251330 467316
rect 365254 467304 365260 467316
rect 365312 467304 365318 467356
rect 44910 467236 44916 467288
rect 44968 467276 44974 467288
rect 104986 467276 104992 467288
rect 44968 467248 104992 467276
rect 44968 467236 44974 467248
rect 104986 467236 104992 467248
rect 105044 467236 105050 467288
rect 180150 467236 180156 467288
rect 180208 467276 180214 467288
rect 218054 467276 218060 467288
rect 180208 467248 218060 467276
rect 180208 467236 180214 467248
rect 218054 467236 218060 467248
rect 218112 467236 218118 467288
rect 251174 467236 251180 467288
rect 251232 467276 251238 467288
rect 366818 467276 366824 467288
rect 251232 467248 366824 467276
rect 251232 467236 251238 467248
rect 366818 467236 366824 467248
rect 366876 467236 366882 467288
rect 45278 467168 45284 467220
rect 45336 467208 45342 467220
rect 106366 467208 106372 467220
rect 45336 467180 106372 467208
rect 45336 467168 45342 467180
rect 106366 467168 106372 467180
rect 106424 467168 106430 467220
rect 149054 467168 149060 467220
rect 149112 467208 149118 467220
rect 212902 467208 212908 467220
rect 149112 467180 212908 467208
rect 149112 467168 149118 467180
rect 212902 467168 212908 467180
rect 212960 467168 212966 467220
rect 253934 467168 253940 467220
rect 253992 467208 253998 467220
rect 369578 467208 369584 467220
rect 253992 467180 369584 467208
rect 253992 467168 253998 467180
rect 369578 467168 369584 467180
rect 369636 467168 369642 467220
rect 45186 467100 45192 467152
rect 45244 467140 45250 467152
rect 106458 467140 106464 467152
rect 45244 467112 106464 467140
rect 45244 467100 45250 467112
rect 106458 467100 106464 467112
rect 106516 467100 106522 467152
rect 146294 467100 146300 467152
rect 146352 467140 146358 467152
rect 218698 467140 218704 467152
rect 146352 467112 218704 467140
rect 146352 467100 146358 467112
rect 218698 467100 218704 467112
rect 218756 467100 218762 467152
rect 262214 467100 262220 467152
rect 262272 467140 262278 467152
rect 379146 467140 379152 467152
rect 262272 467112 379152 467140
rect 262272 467100 262278 467112
rect 379146 467100 379152 467112
rect 379204 467100 379210 467152
rect 59262 467032 59268 467084
rect 59320 467072 59326 467084
rect 67726 467072 67732 467084
rect 59320 467044 67732 467072
rect 59320 467032 59326 467044
rect 67726 467032 67732 467044
rect 67784 467032 67790 467084
rect 59170 466964 59176 467016
rect 59228 467004 59234 467016
rect 66346 467004 66352 467016
rect 59228 466976 66352 467004
rect 59228 466964 59234 466976
rect 66346 466964 66352 466976
rect 66404 466964 66410 467016
rect 178034 466556 178040 466608
rect 178092 466596 178098 466608
rect 204622 466596 204628 466608
rect 178092 466568 204628 466596
rect 178092 466556 178098 466568
rect 204622 466556 204628 466568
rect 204680 466596 204686 466608
rect 338482 466596 338488 466608
rect 204680 466568 338488 466596
rect 204680 466556 204686 466568
rect 338482 466556 338488 466568
rect 338540 466596 338546 466608
rect 356974 466596 356980 466608
rect 338540 466568 356980 466596
rect 338540 466556 338546 466568
rect 356974 466556 356980 466568
rect 357032 466596 357038 466608
rect 498470 466596 498476 466608
rect 357032 466568 498476 466596
rect 357032 466556 357038 466568
rect 498470 466556 498476 466568
rect 498528 466596 498534 466608
rect 517790 466596 517796 466608
rect 498528 466568 517796 466596
rect 498528 466556 498534 466568
rect 517790 466556 517796 466568
rect 517848 466556 517854 466608
rect 48866 466488 48872 466540
rect 48924 466528 48930 466540
rect 48924 466500 207152 466528
rect 48924 466488 48930 466500
rect 207124 466472 207152 466500
rect 218054 466488 218060 466540
rect 218112 466528 218118 466540
rect 218238 466528 218244 466540
rect 218112 466500 218244 466528
rect 218112 466488 218118 466500
rect 218238 466488 218244 466500
rect 218296 466528 218302 466540
rect 339770 466528 339776 466540
rect 218296 466500 339776 466528
rect 218296 466488 218302 466500
rect 339770 466488 339776 466500
rect 339828 466528 339834 466540
rect 357526 466528 357532 466540
rect 339828 466500 357532 466528
rect 339828 466488 339834 466500
rect 357526 466488 357532 466500
rect 357584 466528 357590 466540
rect 499758 466528 499764 466540
rect 357584 466500 499764 466528
rect 357584 466488 357590 466500
rect 499758 466488 499764 466500
rect 499816 466528 499822 466540
rect 499816 466500 509234 466528
rect 499816 466488 499822 466500
rect 190914 466420 190920 466472
rect 190972 466460 190978 466472
rect 206278 466460 206284 466472
rect 190972 466432 206284 466460
rect 190972 466420 190978 466432
rect 206278 466420 206284 466432
rect 206336 466420 206342 466472
rect 207106 466420 207112 466472
rect 207164 466460 207170 466472
rect 208118 466460 208124 466472
rect 207164 466432 208124 466460
rect 207164 466420 207170 466432
rect 208118 466420 208124 466432
rect 208176 466420 208182 466472
rect 350994 466420 351000 466472
rect 351052 466460 351058 466472
rect 358814 466460 358820 466472
rect 351052 466432 358820 466460
rect 351052 466420 351058 466432
rect 358814 466420 358820 466432
rect 358872 466420 358878 466472
rect 509206 466460 509234 466500
rect 510890 466488 510896 466540
rect 510948 466528 510954 466540
rect 517514 466528 517520 466540
rect 510948 466500 517520 466528
rect 510948 466488 510954 466500
rect 517514 466488 517520 466500
rect 517572 466488 517578 466540
rect 517882 466460 517888 466472
rect 509206 466432 517888 466460
rect 517882 466420 517888 466432
rect 517940 466420 517946 466472
rect 52270 466352 52276 466404
rect 52328 466392 52334 466404
rect 77294 466392 77300 466404
rect 52328 466364 77300 466392
rect 52328 466352 52334 466364
rect 77294 466352 77300 466364
rect 77352 466352 77358 466404
rect 193306 466352 193312 466404
rect 193364 466392 193370 466404
rect 213086 466392 213092 466404
rect 193364 466364 213092 466392
rect 193364 466352 193370 466364
rect 213086 466352 213092 466364
rect 213144 466352 213150 466404
rect 295426 466352 295432 466404
rect 295484 466392 295490 466404
rect 357250 466392 357256 466404
rect 295484 466364 357256 466392
rect 295484 466352 295490 466364
rect 357250 466352 357256 466364
rect 357308 466352 357314 466404
rect 51994 466284 52000 466336
rect 52052 466324 52058 466336
rect 75914 466324 75920 466336
rect 52052 466296 75920 466324
rect 52052 466284 52058 466296
rect 75914 466284 75920 466296
rect 75972 466284 75978 466336
rect 180978 466284 180984 466336
rect 181036 466324 181042 466336
rect 207934 466324 207940 466336
rect 181036 466296 207940 466324
rect 181036 466284 181042 466296
rect 207934 466284 207940 466296
rect 207992 466284 207998 466336
rect 271966 466284 271972 466336
rect 272024 466324 272030 466336
rect 366174 466324 366180 466336
rect 272024 466296 366180 466324
rect 272024 466284 272030 466296
rect 366174 466284 366180 466296
rect 366232 466284 366238 466336
rect 189074 466216 189080 466268
rect 189132 466256 189138 466268
rect 217594 466256 217600 466268
rect 189132 466228 217600 466256
rect 189132 466216 189138 466228
rect 217594 466216 217600 466228
rect 217652 466216 217658 466268
rect 258074 466216 258080 466268
rect 258132 466256 258138 466268
rect 364150 466256 364156 466268
rect 258132 466228 364156 466256
rect 258132 466216 258138 466228
rect 364150 466216 364156 466228
rect 364208 466216 364214 466268
rect 54386 466148 54392 466200
rect 54444 466188 54450 466200
rect 62114 466188 62120 466200
rect 54444 466160 62120 466188
rect 54444 466148 54450 466160
rect 62114 466148 62120 466160
rect 62172 466148 62178 466200
rect 173894 466148 173900 466200
rect 173952 466188 173958 466200
rect 203886 466188 203892 466200
rect 173952 466160 203892 466188
rect 173952 466148 173958 466160
rect 203886 466148 203892 466160
rect 203944 466148 203950 466200
rect 260834 466148 260840 466200
rect 260892 466188 260898 466200
rect 376386 466188 376392 466200
rect 260892 466160 376392 466188
rect 260892 466148 260898 466160
rect 376386 466148 376392 466160
rect 376444 466148 376450 466200
rect 54294 466080 54300 466132
rect 54352 466120 54358 466132
rect 63494 466120 63500 466132
rect 54352 466092 63500 466120
rect 54352 466080 54358 466092
rect 63494 466080 63500 466092
rect 63552 466080 63558 466132
rect 180886 466080 180892 466132
rect 180944 466120 180950 466132
rect 210970 466120 210976 466132
rect 180944 466092 210976 466120
rect 180944 466080 180950 466092
rect 210970 466080 210976 466092
rect 211028 466080 211034 466132
rect 249794 466080 249800 466132
rect 249852 466120 249858 466132
rect 366542 466120 366548 466132
rect 249852 466092 366548 466120
rect 249852 466080 249858 466092
rect 366542 466080 366548 466092
rect 366600 466080 366606 466132
rect 51442 466012 51448 466064
rect 51500 466052 51506 466064
rect 66254 466052 66260 466064
rect 51500 466024 66260 466052
rect 51500 466012 51506 466024
rect 66254 466012 66260 466024
rect 66312 466012 66318 466064
rect 172514 466012 172520 466064
rect 172572 466052 172578 466064
rect 204898 466052 204904 466064
rect 172572 466024 204904 466052
rect 172572 466012 172578 466024
rect 204898 466012 204904 466024
rect 204956 466012 204962 466064
rect 245654 466012 245660 466064
rect 245712 466052 245718 466064
rect 362494 466052 362500 466064
rect 245712 466024 362500 466052
rect 245712 466012 245718 466024
rect 362494 466012 362500 466024
rect 362552 466012 362558 466064
rect 42058 465944 42064 465996
rect 42116 465984 42122 465996
rect 60734 465984 60740 465996
rect 42116 465956 60740 465984
rect 42116 465944 42122 465956
rect 60734 465944 60740 465956
rect 60792 465944 60798 465996
rect 179414 465944 179420 465996
rect 179472 465984 179478 465996
rect 219066 465984 219072 465996
rect 179472 465956 219072 465984
rect 179472 465944 179478 465956
rect 219066 465944 219072 465956
rect 219124 465944 219130 465996
rect 249886 465944 249892 465996
rect 249944 465984 249950 465996
rect 367922 465984 367928 465996
rect 249944 465956 367928 465984
rect 249944 465944 249950 465956
rect 367922 465944 367928 465956
rect 367980 465944 367986 465996
rect 43346 465876 43352 465928
rect 43404 465916 43410 465928
rect 62206 465916 62212 465928
rect 43404 465888 62212 465916
rect 43404 465876 43410 465888
rect 62206 465876 62212 465888
rect 62264 465876 62270 465928
rect 173986 465876 173992 465928
rect 174044 465916 174050 465928
rect 214834 465916 214840 465928
rect 174044 465888 214840 465916
rect 174044 465876 174050 465888
rect 214834 465876 214840 465888
rect 214892 465876 214898 465928
rect 248506 465876 248512 465928
rect 248564 465916 248570 465928
rect 372062 465916 372068 465928
rect 248564 465888 372068 465916
rect 248564 465876 248570 465888
rect 372062 465876 372068 465888
rect 372120 465876 372126 465928
rect 56042 465808 56048 465860
rect 56100 465848 56106 465860
rect 89806 465848 89812 465860
rect 56100 465820 89812 465848
rect 56100 465808 56106 465820
rect 89806 465808 89812 465820
rect 89864 465808 89870 465860
rect 142246 465808 142252 465860
rect 142304 465848 142310 465860
rect 207106 465848 207112 465860
rect 142304 465820 207112 465848
rect 142304 465808 142310 465820
rect 207106 465808 207112 465820
rect 207164 465808 207170 465860
rect 248598 465808 248604 465860
rect 248656 465848 248662 465860
rect 373442 465848 373448 465860
rect 248656 465820 373448 465848
rect 248656 465808 248662 465820
rect 373442 465808 373448 465820
rect 373500 465808 373506 465860
rect 50798 465740 50804 465792
rect 50856 465780 50862 465792
rect 50982 465780 50988 465792
rect 50856 465752 50988 465780
rect 50856 465740 50862 465752
rect 50982 465740 50988 465752
rect 51040 465740 51046 465792
rect 51534 465740 51540 465792
rect 51592 465780 51598 465792
rect 51994 465780 52000 465792
rect 51592 465752 52000 465780
rect 51592 465740 51598 465752
rect 51994 465740 52000 465752
rect 52052 465740 52058 465792
rect 58802 465740 58808 465792
rect 58860 465780 58866 465792
rect 95418 465780 95424 465792
rect 58860 465752 95424 465780
rect 58860 465740 58866 465752
rect 95418 465740 95424 465752
rect 95476 465740 95482 465792
rect 107654 465740 107660 465792
rect 107712 465780 107718 465792
rect 201770 465780 201776 465792
rect 107712 465752 201776 465780
rect 107712 465740 107718 465752
rect 201770 465740 201776 465752
rect 201828 465740 201834 465792
rect 208302 465740 208308 465792
rect 208360 465780 208366 465792
rect 220998 465780 221004 465792
rect 208360 465752 221004 465780
rect 208360 465740 208366 465752
rect 220998 465740 221004 465752
rect 221056 465740 221062 465792
rect 241514 465740 241520 465792
rect 241572 465780 241578 465792
rect 369394 465780 369400 465792
rect 241572 465752 369400 465780
rect 241572 465740 241578 465752
rect 369394 465740 369400 465752
rect 369452 465740 369458 465792
rect 49510 465672 49516 465724
rect 49568 465712 49574 465724
rect 70394 465712 70400 465724
rect 49568 465684 70400 465712
rect 49568 465672 49574 465684
rect 70394 465672 70400 465684
rect 70452 465672 70458 465724
rect 72418 465672 72424 465724
rect 72476 465712 72482 465724
rect 198826 465712 198832 465724
rect 72476 465684 198832 465712
rect 72476 465672 72482 465684
rect 198826 465672 198832 465684
rect 198884 465672 198890 465724
rect 205358 465672 205364 465724
rect 205416 465712 205422 465724
rect 220906 465712 220912 465724
rect 205416 465684 220912 465712
rect 205416 465672 205422 465684
rect 220906 465672 220912 465684
rect 220964 465672 220970 465724
rect 242894 465672 242900 465724
rect 242952 465712 242958 465724
rect 374822 465712 374828 465724
rect 242952 465684 374828 465712
rect 242952 465672 242958 465684
rect 374822 465672 374828 465684
rect 374880 465672 374886 465724
rect 186314 465604 186320 465656
rect 186372 465644 186378 465656
rect 202506 465644 202512 465656
rect 186372 465616 202512 465644
rect 186372 465604 186378 465616
rect 202506 465604 202512 465616
rect 202564 465604 202570 465656
rect 187786 465536 187792 465588
rect 187844 465576 187850 465588
rect 200942 465576 200948 465588
rect 187844 465548 200948 465576
rect 187844 465536 187850 465548
rect 200942 465536 200948 465548
rect 201000 465536 201006 465588
rect 194594 465468 194600 465520
rect 194652 465508 194658 465520
rect 206646 465508 206652 465520
rect 194652 465480 206652 465508
rect 194652 465468 194658 465480
rect 206646 465468 206652 465480
rect 206704 465468 206710 465520
rect 198826 465060 198832 465112
rect 198884 465100 198890 465112
rect 199010 465100 199016 465112
rect 198884 465072 199016 465100
rect 198884 465060 198890 465072
rect 199010 465060 199016 465072
rect 199068 465100 199074 465112
rect 358906 465100 358912 465112
rect 199068 465072 358912 465100
rect 199068 465060 199074 465072
rect 358906 465060 358912 465072
rect 358964 465100 358970 465112
rect 518894 465100 518900 465112
rect 358964 465072 518900 465100
rect 358964 465060 358970 465072
rect 518894 465060 518900 465072
rect 518952 465060 518958 465112
rect 190454 464788 190460 464840
rect 190512 464828 190518 464840
rect 208946 464828 208952 464840
rect 190512 464800 208952 464828
rect 190512 464788 190518 464800
rect 208946 464788 208952 464800
rect 209004 464788 209010 464840
rect 58986 464720 58992 464772
rect 59044 464760 59050 464772
rect 89898 464760 89904 464772
rect 59044 464732 89904 464760
rect 59044 464720 59050 464732
rect 89898 464720 89904 464732
rect 89956 464720 89962 464772
rect 185578 464720 185584 464772
rect 185636 464760 185642 464772
rect 204714 464760 204720 464772
rect 185636 464732 204720 464760
rect 185636 464720 185642 464732
rect 204714 464720 204720 464732
rect 204772 464720 204778 464772
rect 58894 464652 58900 464704
rect 58952 464692 58958 464704
rect 92658 464692 92664 464704
rect 58952 464664 92664 464692
rect 58952 464652 58958 464664
rect 92658 464652 92664 464664
rect 92716 464652 92722 464704
rect 193214 464652 193220 464704
rect 193272 464692 193278 464704
rect 214282 464692 214288 464704
rect 193272 464664 214288 464692
rect 193272 464652 193278 464664
rect 214282 464652 214288 464664
rect 214340 464652 214346 464704
rect 55858 464584 55864 464636
rect 55916 464624 55922 464636
rect 102318 464624 102324 464636
rect 55916 464596 102324 464624
rect 55916 464584 55922 464596
rect 102318 464584 102324 464596
rect 102376 464584 102382 464636
rect 180794 464584 180800 464636
rect 180852 464624 180858 464636
rect 209314 464624 209320 464636
rect 180852 464596 209320 464624
rect 180852 464584 180858 464596
rect 209314 464584 209320 464596
rect 209372 464584 209378 464636
rect 54570 464516 54576 464568
rect 54628 464556 54634 464568
rect 102226 464556 102232 464568
rect 54628 464528 102232 464556
rect 54628 464516 54634 464528
rect 102226 464516 102232 464528
rect 102284 464516 102290 464568
rect 142154 464516 142160 464568
rect 142212 464556 142218 464568
rect 198090 464556 198096 464568
rect 142212 464528 198096 464556
rect 142212 464516 142218 464528
rect 198090 464516 198096 464528
rect 198148 464516 198154 464568
rect 52914 464448 52920 464500
rect 52972 464488 52978 464500
rect 121454 464488 121460 464500
rect 52972 464460 121460 464488
rect 52972 464448 52978 464460
rect 121454 464448 121460 464460
rect 121512 464448 121518 464500
rect 125594 464448 125600 464500
rect 125652 464488 125658 464500
rect 197814 464488 197820 464500
rect 125652 464460 197820 464488
rect 125652 464448 125658 464460
rect 197814 464448 197820 464460
rect 197872 464448 197878 464500
rect 295334 464448 295340 464500
rect 295392 464488 295398 464500
rect 360654 464488 360660 464500
rect 295392 464460 360660 464488
rect 295392 464448 295398 464460
rect 360654 464448 360660 464460
rect 360712 464448 360718 464500
rect 57054 464380 57060 464432
rect 57112 464420 57118 464432
rect 131114 464420 131120 464432
rect 57112 464392 131120 464420
rect 57112 464380 57118 464392
rect 131114 464380 131120 464392
rect 131172 464380 131178 464432
rect 138014 464380 138020 464432
rect 138072 464420 138078 464432
rect 200574 464420 200580 464432
rect 138072 464392 200580 464420
rect 138072 464380 138078 464392
rect 200574 464380 200580 464392
rect 200632 464380 200638 464432
rect 291194 464380 291200 464432
rect 291252 464420 291258 464432
rect 364886 464420 364892 464432
rect 291252 464392 364892 464420
rect 291252 464380 291258 464392
rect 364886 464380 364892 464392
rect 364944 464380 364950 464432
rect 57146 464312 57152 464364
rect 57204 464352 57210 464364
rect 132494 464352 132500 464364
rect 57204 464324 132500 464352
rect 57204 464312 57210 464324
rect 132494 464312 132500 464324
rect 132552 464312 132558 464364
rect 136634 464312 136640 464364
rect 136692 464352 136698 464364
rect 199562 464352 199568 464364
rect 136692 464324 199568 464352
rect 136692 464312 136698 464324
rect 199562 464312 199568 464324
rect 199620 464312 199626 464364
rect 271874 464312 271880 464364
rect 271932 464352 271938 464364
rect 371602 464352 371608 464364
rect 271932 464324 371608 464352
rect 271932 464312 271938 464324
rect 371602 464312 371608 464324
rect 371660 464312 371666 464364
rect 519538 460164 519544 460216
rect 519596 460204 519602 460216
rect 580350 460204 580356 460216
rect 519596 460176 580356 460204
rect 519596 460164 519602 460176
rect 580350 460164 580356 460176
rect 580408 460164 580414 460216
rect 48866 418072 48872 418124
rect 48924 418112 48930 418124
rect 57054 418112 57060 418124
rect 48924 418084 57060 418112
rect 48924 418072 48930 418084
rect 57054 418072 57060 418084
rect 57112 418072 57118 418124
rect 204530 417732 204536 417784
rect 204588 417772 204594 417784
rect 208210 417772 208216 417784
rect 204588 417744 208216 417772
rect 204588 417732 204594 417744
rect 208210 417732 208216 417744
rect 208268 417732 208274 417784
rect 208118 417392 208124 417444
rect 208176 417432 208182 417444
rect 216674 417432 216680 417444
rect 208176 417404 216680 417432
rect 208176 417392 208182 417404
rect 216674 417392 216680 417404
rect 216732 417392 216738 417444
rect 359734 417392 359740 417444
rect 359792 417432 359798 417444
rect 377214 417432 377220 417444
rect 359792 417404 377220 417432
rect 359792 417392 359798 417404
rect 377214 417392 377220 417404
rect 377272 417392 377278 417444
rect 55766 417120 55772 417172
rect 55824 417160 55830 417172
rect 57238 417160 57244 417172
rect 55824 417132 57244 417160
rect 55824 417120 55830 417132
rect 57238 417120 57244 417132
rect 57296 417120 57302 417172
rect 44634 416780 44640 416832
rect 44692 416820 44698 416832
rect 57238 416820 57244 416832
rect 44692 416792 57244 416820
rect 44692 416780 44698 416792
rect 57238 416780 57244 416792
rect 57296 416780 57302 416832
rect 56870 416168 56876 416220
rect 56928 416208 56934 416220
rect 59630 416208 59636 416220
rect 56928 416180 59636 416208
rect 56928 416168 56934 416180
rect 59630 416168 59636 416180
rect 59688 416168 59694 416220
rect 205726 414808 205732 414860
rect 205784 414848 205790 414860
rect 217134 414848 217140 414860
rect 205784 414820 217140 414848
rect 205784 414808 205790 414820
rect 217134 414808 217140 414820
rect 217192 414808 217198 414860
rect 205450 414672 205456 414724
rect 205508 414712 205514 414724
rect 216766 414712 216772 414724
rect 205508 414684 216772 414712
rect 205508 414672 205514 414684
rect 216766 414672 216772 414684
rect 216824 414672 216830 414724
rect 51534 413992 51540 414044
rect 51592 414032 51598 414044
rect 57054 414032 57060 414044
rect 51592 414004 57060 414032
rect 51592 413992 51598 414004
rect 57054 413992 57060 414004
rect 57112 413992 57118 414044
rect 55674 413924 55680 413976
rect 55732 413964 55738 413976
rect 56962 413964 56968 413976
rect 55732 413936 56968 413964
rect 55732 413924 55738 413936
rect 56962 413924 56968 413936
rect 57020 413924 57026 413976
rect 205634 413244 205640 413296
rect 205692 413284 205698 413296
rect 216858 413284 216864 413296
rect 205692 413256 216864 413284
rect 205692 413244 205698 413256
rect 216858 413244 216864 413256
rect 216916 413244 216922 413296
rect 50154 412700 50160 412752
rect 50212 412740 50218 412752
rect 57238 412740 57244 412752
rect 50212 412712 57244 412740
rect 50212 412700 50218 412712
rect 57238 412700 57244 412712
rect 57296 412700 57302 412752
rect 358078 411884 358084 411936
rect 358136 411924 358142 411936
rect 377214 411924 377220 411936
rect 358136 411896 377220 411924
rect 358136 411884 358142 411896
rect 377214 411884 377220 411896
rect 377272 411884 377278 411936
rect 204438 411544 204444 411596
rect 204496 411584 204502 411596
rect 205634 411584 205640 411596
rect 204496 411556 205640 411584
rect 204496 411544 204502 411556
rect 205634 411544 205640 411556
rect 205692 411544 205698 411596
rect 49602 411272 49608 411324
rect 49660 411312 49666 411324
rect 57238 411312 57244 411324
rect 49660 411284 57244 411312
rect 49660 411272 49666 411284
rect 57238 411272 57244 411284
rect 57296 411272 57302 411324
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 15838 411244 15844 411256
rect 3016 411216 15844 411244
rect 3016 411204 3022 411216
rect 15838 411204 15844 411216
rect 15896 411204 15902 411256
rect 52270 411068 52276 411120
rect 52328 411108 52334 411120
rect 53006 411108 53012 411120
rect 52328 411080 53012 411108
rect 52328 411068 52334 411080
rect 53006 411068 53012 411080
rect 53064 411068 53070 411120
rect 206738 410660 206744 410712
rect 206796 410700 206802 410712
rect 216950 410700 216956 410712
rect 206796 410672 216956 410700
rect 206796 410660 206802 410672
rect 216950 410660 216956 410672
rect 217008 410660 217014 410712
rect 205634 410524 205640 410576
rect 205692 410564 205698 410576
rect 216674 410564 216680 410576
rect 205692 410536 216680 410564
rect 205692 410524 205698 410536
rect 216674 410524 216680 410536
rect 216732 410524 216738 410576
rect 359918 410524 359924 410576
rect 359976 410564 359982 410576
rect 377214 410564 377220 410576
rect 359976 410536 377220 410564
rect 359976 410524 359982 410536
rect 377214 410524 377220 410536
rect 377272 410564 377278 410576
rect 377674 410564 377680 410576
rect 377272 410536 377680 410564
rect 377272 410524 377278 410536
rect 377674 410524 377680 410536
rect 377732 410524 377738 410576
rect 217686 410048 217692 410100
rect 217744 410088 217750 410100
rect 219250 410088 219256 410100
rect 217744 410060 219256 410088
rect 217744 410048 217750 410060
rect 219250 410048 219256 410060
rect 219308 410048 219314 410100
rect 48866 409844 48872 409896
rect 48924 409884 48930 409896
rect 56686 409884 56692 409896
rect 48924 409856 56692 409884
rect 48924 409844 48930 409856
rect 56686 409844 56692 409856
rect 56744 409844 56750 409896
rect 208210 409096 208216 409148
rect 208268 409136 208274 409148
rect 216674 409136 216680 409148
rect 208268 409108 216680 409136
rect 208268 409096 208274 409108
rect 216674 409096 216680 409108
rect 216732 409096 216738 409148
rect 359826 409096 359832 409148
rect 359884 409136 359890 409148
rect 377398 409136 377404 409148
rect 359884 409108 377404 409136
rect 359884 409096 359890 409108
rect 377398 409096 377404 409108
rect 377456 409096 377462 409148
rect 52362 408484 52368 408536
rect 52420 408524 52426 408536
rect 57238 408524 57244 408536
rect 52420 408496 57244 408524
rect 52420 408484 52426 408496
rect 57238 408484 57244 408496
rect 57296 408484 57302 408536
rect 198826 400868 198832 400920
rect 198884 400908 198890 400920
rect 199470 400908 199476 400920
rect 198884 400880 199476 400908
rect 198884 400868 198890 400880
rect 199470 400868 199476 400880
rect 199528 400908 199534 400920
rect 207198 400908 207204 400920
rect 199528 400880 207204 400908
rect 199528 400868 199534 400880
rect 207198 400868 207204 400880
rect 207256 400868 207262 400920
rect 520918 396720 520924 396772
rect 520976 396760 520982 396772
rect 580350 396760 580356 396772
rect 520976 396732 580356 396760
rect 520976 396720 520982 396732
rect 580350 396720 580356 396732
rect 580408 396720 580414 396772
rect 198182 396312 198188 396364
rect 198240 396352 198246 396364
rect 199194 396352 199200 396364
rect 198240 396324 199200 396352
rect 198240 396312 198246 396324
rect 199194 396312 199200 396324
rect 199252 396312 199258 396364
rect 197998 395972 198004 396024
rect 198056 396012 198062 396024
rect 198826 396012 198832 396024
rect 198056 395984 198832 396012
rect 198056 395972 198062 395984
rect 198826 395972 198832 395984
rect 198884 395972 198890 396024
rect 198274 395496 198280 395548
rect 198332 395536 198338 395548
rect 199562 395536 199568 395548
rect 198332 395508 199568 395536
rect 198332 395496 198338 395508
rect 199562 395496 199568 395508
rect 199620 395496 199626 395548
rect 44726 391892 44732 391944
rect 44784 391932 44790 391944
rect 57238 391932 57244 391944
rect 44784 391904 57244 391932
rect 44784 391892 44790 391904
rect 57238 391892 57244 391904
rect 57296 391892 57302 391944
rect 209406 391892 209412 391944
rect 209464 391932 209470 391944
rect 216674 391932 216680 391944
rect 209464 391904 216680 391932
rect 209464 391892 209470 391904
rect 216674 391892 216680 391904
rect 216732 391892 216738 391944
rect 359458 391892 359464 391944
rect 359516 391932 359522 391944
rect 376938 391932 376944 391944
rect 359516 391904 376944 391932
rect 359516 391892 359522 391904
rect 376938 391892 376944 391904
rect 376996 391892 377002 391944
rect 358814 390464 358820 390516
rect 358872 390504 358878 390516
rect 376938 390504 376944 390516
rect 358872 390476 376944 390504
rect 358872 390464 358878 390476
rect 376938 390464 376944 390476
rect 376996 390464 377002 390516
rect 206278 389784 206284 389836
rect 206336 389824 206342 389836
rect 216674 389824 216680 389836
rect 206336 389796 216680 389824
rect 206336 389784 206342 389796
rect 216674 389784 216680 389796
rect 216732 389784 216738 389836
rect 57054 389512 57060 389564
rect 57112 389552 57118 389564
rect 57422 389552 57428 389564
rect 57112 389524 57428 389552
rect 57112 389512 57118 389524
rect 57422 389512 57428 389524
rect 57480 389512 57486 389564
rect 358078 389172 358084 389224
rect 358136 389212 358142 389224
rect 358814 389212 358820 389224
rect 358136 389184 358820 389212
rect 358136 389172 358142 389184
rect 358814 389172 358820 389184
rect 358872 389172 358878 389224
rect 53742 389104 53748 389156
rect 53800 389144 53806 389156
rect 57238 389144 57244 389156
rect 53800 389116 57244 389144
rect 53800 389104 53806 389116
rect 57238 389104 57244 389116
rect 57296 389144 57302 389156
rect 57514 389144 57520 389156
rect 57296 389116 57520 389144
rect 57296 389104 57302 389116
rect 57514 389104 57520 389116
rect 57572 389104 57578 389156
rect 200758 389104 200764 389156
rect 200816 389144 200822 389156
rect 217686 389144 217692 389156
rect 200816 389116 217692 389144
rect 200816 389104 200822 389116
rect 217686 389104 217692 389116
rect 217744 389104 217750 389156
rect 359642 389104 359648 389156
rect 359700 389144 359706 389156
rect 376938 389144 376944 389156
rect 359700 389116 376944 389144
rect 359700 389104 359706 389116
rect 376938 389104 376944 389116
rect 376996 389104 377002 389156
rect 46106 389036 46112 389088
rect 46164 389076 46170 389088
rect 57146 389076 57152 389088
rect 46164 389048 57152 389076
rect 46164 389036 46170 389048
rect 57146 389036 57152 389048
rect 57204 389036 57210 389088
rect 57054 388356 57060 388408
rect 57112 388396 57118 388408
rect 57422 388396 57428 388408
rect 57112 388368 57428 388396
rect 57112 388356 57118 388368
rect 57422 388356 57428 388368
rect 57480 388356 57486 388408
rect 199286 384276 199292 384328
rect 199344 384316 199350 384328
rect 199654 384316 199660 384328
rect 199344 384288 199660 384316
rect 199344 384276 199350 384288
rect 199654 384276 199660 384288
rect 199712 384276 199718 384328
rect 197170 382168 197176 382220
rect 197228 382208 197234 382220
rect 197906 382208 197912 382220
rect 197228 382180 197912 382208
rect 197228 382168 197234 382180
rect 197906 382168 197912 382180
rect 197964 382168 197970 382220
rect 58526 381828 58532 381880
rect 58584 381868 58590 381880
rect 59630 381868 59636 381880
rect 58584 381840 59636 381868
rect 58584 381828 58590 381840
rect 59630 381828 59636 381840
rect 59688 381828 59694 381880
rect 55858 381692 55864 381744
rect 55916 381732 55922 381744
rect 59354 381732 59360 381744
rect 55916 381704 59360 381732
rect 55916 381692 55922 381704
rect 59354 381692 59360 381704
rect 59412 381692 59418 381744
rect 205542 381488 205548 381540
rect 205600 381528 205606 381540
rect 212902 381528 212908 381540
rect 205600 381500 212908 381528
rect 205600 381488 205606 381500
rect 212902 381488 212908 381500
rect 212960 381488 212966 381540
rect 362034 381488 362040 381540
rect 362092 381528 362098 381540
rect 369854 381528 369860 381540
rect 362092 381500 369860 381528
rect 362092 381488 362098 381500
rect 369854 381488 369860 381500
rect 369912 381488 369918 381540
rect 218238 381052 218244 381064
rect 195900 381024 218244 381052
rect 195900 380996 195928 381024
rect 218238 381012 218244 381024
rect 218296 381012 218302 381064
rect 57330 380944 57336 380996
rect 57388 380984 57394 380996
rect 59446 380984 59452 380996
rect 57388 380956 59452 380984
rect 57388 380944 57394 380956
rect 59446 380944 59452 380956
rect 59504 380944 59510 380996
rect 195882 380944 195888 380996
rect 195940 380944 195946 380996
rect 219526 380944 219532 380996
rect 219584 380984 219590 380996
rect 220078 380984 220084 380996
rect 219584 380956 220084 380984
rect 219584 380944 219590 380956
rect 220078 380944 220084 380956
rect 220136 380944 220142 380996
rect 58434 380876 58440 380928
rect 58492 380916 58498 380928
rect 60734 380916 60740 380928
rect 58492 380888 60740 380916
rect 58492 380876 58498 380888
rect 60734 380876 60740 380888
rect 60792 380876 60798 380928
rect 208394 380876 208400 380928
rect 208452 380916 208458 380928
rect 208670 380916 208676 380928
rect 208452 380888 208676 380916
rect 208452 380876 208458 380888
rect 208670 380876 208676 380888
rect 208728 380876 208734 380928
rect 217594 380876 217600 380928
rect 217652 380916 217658 380928
rect 248230 380916 248236 380928
rect 217652 380888 248236 380916
rect 217652 380876 217658 380888
rect 248230 380876 248236 380888
rect 248288 380876 248294 380928
rect 369854 380876 369860 380928
rect 369912 380916 369918 380928
rect 371050 380916 371056 380928
rect 369912 380888 371056 380916
rect 369912 380876 369918 380888
rect 371050 380876 371056 380888
rect 371108 380916 371114 380928
rect 431126 380916 431132 380928
rect 371108 380888 431132 380916
rect 371108 380876 371114 380888
rect 431126 380876 431132 380888
rect 431184 380876 431190 380928
rect 44634 380808 44640 380860
rect 44692 380848 44698 380860
rect 217226 380848 217232 380860
rect 44692 380820 217232 380848
rect 44692 380808 44698 380820
rect 217226 380808 217232 380820
rect 217284 380808 217290 380860
rect 219158 380808 219164 380860
rect 219216 380848 219222 380860
rect 219342 380848 219348 380860
rect 219216 380820 219348 380848
rect 219216 380808 219222 380820
rect 219342 380808 219348 380820
rect 219400 380808 219406 380860
rect 219894 380808 219900 380860
rect 219952 380848 219958 380860
rect 220722 380848 220728 380860
rect 219952 380820 220728 380848
rect 219952 380808 219958 380820
rect 220722 380808 220728 380820
rect 220780 380808 220786 380860
rect 52914 380740 52920 380792
rect 52972 380780 52978 380792
rect 55858 380780 55864 380792
rect 52972 380752 55864 380780
rect 52972 380740 52978 380752
rect 55858 380740 55864 380752
rect 55916 380740 55922 380792
rect 216858 380780 216864 380792
rect 64846 380752 216864 380780
rect 50154 380672 50160 380724
rect 50212 380712 50218 380724
rect 64846 380712 64874 380752
rect 216858 380740 216864 380752
rect 216916 380780 216922 380792
rect 217686 380780 217692 380792
rect 216916 380752 217692 380780
rect 216916 380740 216922 380752
rect 217686 380740 217692 380752
rect 217744 380740 217750 380792
rect 367002 380740 367008 380792
rect 367060 380780 367066 380792
rect 380986 380780 380992 380792
rect 367060 380752 380992 380780
rect 367060 380740 367066 380752
rect 380986 380740 380992 380752
rect 381044 380740 381050 380792
rect 50212 380684 64874 380712
rect 50212 380672 50218 380684
rect 155954 380672 155960 380724
rect 156012 380712 156018 380724
rect 203150 380712 203156 380724
rect 156012 380684 203156 380712
rect 156012 380672 156018 380684
rect 203150 380672 203156 380684
rect 203208 380672 203214 380724
rect 357986 380672 357992 380724
rect 358044 380712 358050 380724
rect 380894 380712 380900 380724
rect 358044 380684 380900 380712
rect 358044 380672 358050 380684
rect 380894 380672 380900 380684
rect 380952 380672 380958 380724
rect 158530 380604 158536 380656
rect 158588 380644 158594 380656
rect 205910 380644 205916 380656
rect 158588 380616 205916 380644
rect 158588 380604 158594 380616
rect 205910 380604 205916 380616
rect 205968 380604 205974 380656
rect 377306 380604 377312 380656
rect 377364 380644 377370 380656
rect 410702 380644 410708 380656
rect 377364 380616 410708 380644
rect 377364 380604 377370 380616
rect 410702 380604 410708 380616
rect 410760 380604 410766 380656
rect 140958 380536 140964 380588
rect 141016 380576 141022 380588
rect 200574 380576 200580 380588
rect 141016 380548 200580 380576
rect 141016 380536 141022 380548
rect 200574 380536 200580 380548
rect 200632 380536 200638 380588
rect 373902 380536 373908 380588
rect 373960 380576 373966 380588
rect 421098 380576 421104 380588
rect 373960 380548 421104 380576
rect 373960 380536 373966 380548
rect 421098 380536 421104 380548
rect 421156 380536 421162 380588
rect 54478 380468 54484 380520
rect 54536 380508 54542 380520
rect 113542 380508 113548 380520
rect 54536 380480 113548 380508
rect 54536 380468 54542 380480
rect 113542 380468 113548 380480
rect 113600 380468 113606 380520
rect 146018 380468 146024 380520
rect 146076 380508 146082 380520
rect 205818 380508 205824 380520
rect 146076 380480 205824 380508
rect 146076 380468 146082 380480
rect 205818 380468 205824 380480
rect 205876 380468 205882 380520
rect 371602 380468 371608 380520
rect 371660 380508 371666 380520
rect 433610 380508 433616 380520
rect 371660 380480 433616 380508
rect 371660 380468 371666 380480
rect 433610 380468 433616 380480
rect 433668 380468 433674 380520
rect 55950 380400 55956 380452
rect 56008 380440 56014 380452
rect 118418 380440 118424 380452
rect 56008 380412 118424 380440
rect 56008 380400 56014 380412
rect 118418 380400 118424 380412
rect 118476 380400 118482 380452
rect 143534 380400 143540 380452
rect 143592 380440 143598 380452
rect 204714 380440 204720 380452
rect 143592 380412 204720 380440
rect 143592 380400 143598 380412
rect 204714 380400 204720 380412
rect 204772 380400 204778 380452
rect 369026 380400 369032 380452
rect 369084 380440 369090 380452
rect 436002 380440 436008 380452
rect 369084 380412 436008 380440
rect 369084 380400 369090 380412
rect 436002 380400 436008 380412
rect 436060 380400 436066 380452
rect 48958 380332 48964 380384
rect 49016 380372 49022 380384
rect 110966 380372 110972 380384
rect 49016 380344 110972 380372
rect 49016 380332 49022 380344
rect 110966 380332 110972 380344
rect 111024 380332 111030 380384
rect 133506 380332 133512 380384
rect 133564 380372 133570 380384
rect 201862 380372 201868 380384
rect 133564 380344 201868 380372
rect 133564 380332 133570 380344
rect 201862 380332 201868 380344
rect 201920 380332 201926 380384
rect 213638 380332 213644 380384
rect 213696 380372 213702 380384
rect 222010 380372 222016 380384
rect 213696 380344 222016 380372
rect 213696 380332 213702 380344
rect 222010 380332 222016 380344
rect 222068 380332 222074 380384
rect 366174 380332 366180 380384
rect 366232 380372 366238 380384
rect 438486 380372 438492 380384
rect 366232 380344 438492 380372
rect 366232 380332 366238 380344
rect 438486 380332 438492 380344
rect 438544 380332 438550 380384
rect 57422 380264 57428 380316
rect 57480 380304 57486 380316
rect 123478 380304 123484 380316
rect 57480 380276 123484 380304
rect 57480 380264 57486 380276
rect 123478 380264 123484 380276
rect 123536 380264 123542 380316
rect 131022 380264 131028 380316
rect 131080 380304 131086 380316
rect 198274 380304 198280 380316
rect 131080 380276 198280 380304
rect 131080 380264 131086 380276
rect 198274 380264 198280 380276
rect 198332 380264 198338 380316
rect 200114 380264 200120 380316
rect 200172 380304 200178 380316
rect 295334 380304 295340 380316
rect 200172 380276 295340 380304
rect 200172 380264 200178 380276
rect 295334 380264 295340 380276
rect 295392 380264 295398 380316
rect 363414 380264 363420 380316
rect 363472 380304 363478 380316
rect 440878 380304 440884 380316
rect 363472 380276 440884 380304
rect 363472 380264 363478 380276
rect 440878 380264 440884 380276
rect 440936 380264 440942 380316
rect 56870 380196 56876 380248
rect 56928 380236 56934 380248
rect 125962 380236 125968 380248
rect 56928 380208 125968 380236
rect 56928 380196 56934 380208
rect 125962 380196 125968 380208
rect 126020 380196 126026 380248
rect 128354 380196 128360 380248
rect 128412 380236 128418 380248
rect 199102 380236 199108 380248
rect 128412 380208 199108 380236
rect 128412 380196 128418 380208
rect 199102 380196 199108 380208
rect 199160 380196 199166 380248
rect 200206 380196 200212 380248
rect 200264 380236 200270 380248
rect 301498 380236 301504 380248
rect 200264 380208 301504 380236
rect 200264 380196 200270 380208
rect 301498 380196 301504 380208
rect 301556 380196 301562 380248
rect 361482 380196 361488 380248
rect 361540 380236 361546 380248
rect 443454 380236 443460 380248
rect 361540 380208 443460 380236
rect 361540 380196 361546 380208
rect 443454 380196 443460 380208
rect 443512 380196 443518 380248
rect 47578 380128 47584 380180
rect 47636 380168 47642 380180
rect 116026 380168 116032 380180
rect 47636 380140 116032 380168
rect 47636 380128 47642 380140
rect 116026 380128 116032 380140
rect 116084 380128 116090 380180
rect 120994 380128 121000 380180
rect 121052 380168 121058 380180
rect 198826 380168 198832 380180
rect 121052 380140 198832 380168
rect 121052 380128 121058 380140
rect 198826 380128 198832 380140
rect 198884 380128 198890 380180
rect 201678 380128 201684 380180
rect 201736 380168 201742 380180
rect 310422 380168 310428 380180
rect 201736 380140 310428 380168
rect 201736 380128 201742 380140
rect 310422 380128 310428 380140
rect 310480 380128 310486 380180
rect 357066 380128 357072 380180
rect 357124 380168 357130 380180
rect 485958 380168 485964 380180
rect 357124 380140 485964 380168
rect 357124 380128 357130 380140
rect 485958 380128 485964 380140
rect 486016 380128 486022 380180
rect 160922 380060 160928 380112
rect 160980 380100 160986 380112
rect 207106 380100 207112 380112
rect 160980 380072 207112 380100
rect 160980 380060 160986 380072
rect 207106 380060 207112 380072
rect 207164 380060 207170 380112
rect 213546 380060 213552 380112
rect 213604 380100 213610 380112
rect 213822 380100 213828 380112
rect 213604 380072 213828 380100
rect 213604 380060 213610 380072
rect 213822 380060 213828 380072
rect 213880 380100 213886 380112
rect 235994 380100 236000 380112
rect 213880 380072 236000 380100
rect 213880 380060 213886 380072
rect 235994 380060 236000 380072
rect 236052 380060 236058 380112
rect 163406 379992 163412 380044
rect 163464 380032 163470 380044
rect 198090 380032 198096 380044
rect 163464 380004 198096 380032
rect 163464 379992 163470 380004
rect 198090 379992 198096 380004
rect 198148 379992 198154 380044
rect 215846 379992 215852 380044
rect 215904 380032 215910 380044
rect 237098 380032 237104 380044
rect 215904 380004 237104 380032
rect 215904 379992 215910 380004
rect 237098 379992 237104 380004
rect 237156 379992 237162 380044
rect 239122 379992 239128 380044
rect 239180 380032 239186 380044
rect 259454 380032 259460 380044
rect 239180 380004 259460 380032
rect 239180 379992 239186 380004
rect 259454 379992 259460 380004
rect 259512 379992 259518 380044
rect 165982 379924 165988 379976
rect 166040 379964 166046 379976
rect 200482 379964 200488 379976
rect 166040 379936 200488 379964
rect 166040 379924 166046 379936
rect 200482 379924 200488 379936
rect 200540 379924 200546 379976
rect 213822 379924 213828 379976
rect 213880 379964 213886 379976
rect 243078 379964 243084 379976
rect 213880 379936 243084 379964
rect 213880 379924 213886 379936
rect 243078 379924 243084 379936
rect 243136 379924 243142 379976
rect 219802 379856 219808 379908
rect 219860 379896 219866 379908
rect 254486 379896 254492 379908
rect 219860 379868 254492 379896
rect 219860 379856 219866 379868
rect 254486 379856 254492 379868
rect 254544 379856 254550 379908
rect 215294 379788 215300 379840
rect 215352 379828 215358 379840
rect 216214 379828 216220 379840
rect 215352 379800 216220 379828
rect 215352 379788 215358 379800
rect 216214 379788 216220 379800
rect 216272 379828 216278 379840
rect 256970 379828 256976 379840
rect 216272 379800 256976 379828
rect 216272 379788 216278 379800
rect 256970 379788 256976 379800
rect 257028 379788 257034 379840
rect 376478 379788 376484 379840
rect 376536 379828 376542 379840
rect 405458 379828 405464 379840
rect 376536 379800 405464 379828
rect 376536 379788 376542 379800
rect 405458 379788 405464 379800
rect 405516 379788 405522 379840
rect 212534 379720 212540 379772
rect 212592 379760 212598 379772
rect 255866 379760 255872 379772
rect 212592 379732 255872 379760
rect 212592 379720 212598 379732
rect 255866 379720 255872 379732
rect 255924 379720 255930 379772
rect 380986 379720 380992 379772
rect 381044 379760 381050 379772
rect 381354 379760 381360 379772
rect 381044 379732 381360 379760
rect 381044 379720 381050 379732
rect 381354 379720 381360 379732
rect 381412 379760 381418 379772
rect 413462 379760 413468 379772
rect 381412 379732 413468 379760
rect 381412 379720 381418 379732
rect 413462 379720 413468 379732
rect 413520 379720 413526 379772
rect 212626 379652 212632 379704
rect 212684 379692 212690 379704
rect 258074 379692 258080 379704
rect 212684 379664 258080 379692
rect 212684 379652 212690 379664
rect 258074 379652 258080 379664
rect 258132 379652 258138 379704
rect 380894 379652 380900 379704
rect 380952 379692 380958 379704
rect 426434 379692 426440 379704
rect 380952 379664 426440 379692
rect 380952 379652 380958 379664
rect 426434 379652 426440 379664
rect 426492 379652 426498 379704
rect 212718 379584 212724 379636
rect 212776 379624 212782 379636
rect 219802 379624 219808 379636
rect 212776 379596 219808 379624
rect 212776 379584 212782 379596
rect 219802 379584 219808 379596
rect 219860 379584 219866 379636
rect 219894 379584 219900 379636
rect 219952 379624 219958 379636
rect 263870 379624 263876 379636
rect 219952 379596 263876 379624
rect 219952 379584 219958 379596
rect 263870 379584 263876 379596
rect 263928 379584 263934 379636
rect 368382 379584 368388 379636
rect 368440 379624 368446 379636
rect 372522 379624 372528 379636
rect 368440 379596 372528 379624
rect 368440 379584 368446 379596
rect 372522 379584 372528 379596
rect 372580 379624 372586 379636
rect 419442 379624 419448 379636
rect 372580 379596 419448 379624
rect 372580 379584 372586 379596
rect 419442 379584 419448 379596
rect 419500 379584 419506 379636
rect 207106 379516 207112 379568
rect 207164 379556 207170 379568
rect 213822 379556 213828 379568
rect 207164 379528 213828 379556
rect 207164 379516 207170 379528
rect 213822 379516 213828 379528
rect 213880 379516 213886 379568
rect 265250 379556 265256 379568
rect 220004 379528 265256 379556
rect 86586 379448 86592 379500
rect 86644 379488 86650 379500
rect 208486 379488 208492 379500
rect 86644 379460 208492 379488
rect 86644 379448 86650 379460
rect 208486 379448 208492 379460
rect 208544 379488 208550 379500
rect 212442 379488 212448 379500
rect 208544 379460 212448 379488
rect 208544 379448 208550 379460
rect 212442 379448 212448 379460
rect 212500 379448 212506 379500
rect 219342 379448 219348 379500
rect 219400 379488 219406 379500
rect 220004 379488 220032 379528
rect 265250 379516 265256 379528
rect 265308 379516 265314 379568
rect 374546 379516 374552 379568
rect 374604 379556 374610 379568
rect 375098 379556 375104 379568
rect 374604 379528 375104 379556
rect 374604 379516 374610 379528
rect 375098 379516 375104 379528
rect 375156 379556 375162 379568
rect 434346 379556 434352 379568
rect 375156 379528 434352 379556
rect 375156 379516 375162 379528
rect 434346 379516 434352 379528
rect 434404 379516 434410 379568
rect 219400 379460 220032 379488
rect 219400 379448 219406 379460
rect 220078 379448 220084 379500
rect 220136 379488 220142 379500
rect 275646 379488 275652 379500
rect 220136 379460 275652 379488
rect 220136 379448 220142 379460
rect 275646 379448 275652 379460
rect 275704 379448 275710 379500
rect 301498 379448 301504 379500
rect 301556 379488 301562 379500
rect 313366 379488 313372 379500
rect 301556 379460 313372 379488
rect 301556 379448 301562 379460
rect 313366 379448 313372 379460
rect 313424 379448 313430 379500
rect 359550 379448 359556 379500
rect 359608 379488 359614 379500
rect 408310 379488 408316 379500
rect 359608 379460 408316 379488
rect 359608 379448 359614 379460
rect 408310 379448 408316 379460
rect 408368 379448 408374 379500
rect 47762 379380 47768 379432
rect 47820 379420 47826 379432
rect 88334 379420 88340 379432
rect 47820 379392 88340 379420
rect 47820 379380 47826 379392
rect 88334 379380 88340 379392
rect 88392 379380 88398 379432
rect 92382 379380 92388 379432
rect 92440 379420 92446 379432
rect 212810 379420 212816 379432
rect 92440 379392 212816 379420
rect 92440 379380 92446 379392
rect 212810 379380 212816 379392
rect 212868 379420 212874 379432
rect 213822 379420 213828 379432
rect 212868 379392 213828 379420
rect 212868 379380 212874 379392
rect 213822 379380 213828 379392
rect 213880 379380 213886 379432
rect 219434 379380 219440 379432
rect 219492 379420 219498 379432
rect 274358 379420 274364 379432
rect 219492 379392 274364 379420
rect 219492 379380 219498 379392
rect 274358 379380 274364 379392
rect 274416 379380 274422 379432
rect 310422 379380 310428 379432
rect 310480 379420 310486 379432
rect 315758 379420 315764 379432
rect 310480 379392 315764 379420
rect 310480 379380 310486 379392
rect 315758 379380 315764 379392
rect 315816 379380 315822 379432
rect 372430 379380 372436 379432
rect 372488 379420 372494 379432
rect 377398 379420 377404 379432
rect 372488 379392 377404 379420
rect 372488 379380 372494 379392
rect 377398 379380 377404 379392
rect 377456 379380 377462 379432
rect 88794 379312 88800 379364
rect 88852 379352 88858 379364
rect 88852 379324 195974 379352
rect 88852 379312 88858 379324
rect 47670 379244 47676 379296
rect 47728 379284 47734 379296
rect 90634 379284 90640 379296
rect 47728 379256 90640 379284
rect 47728 379244 47734 379256
rect 90634 379244 90640 379256
rect 90692 379244 90698 379296
rect 195946 379284 195974 379324
rect 208486 379312 208492 379364
rect 208544 379352 208550 379364
rect 209590 379352 209596 379364
rect 208544 379324 209596 379352
rect 208544 379312 208550 379324
rect 209590 379312 209596 379324
rect 209648 379352 209654 379364
rect 209648 379324 215294 379352
rect 209648 379312 209654 379324
rect 209866 379284 209872 379296
rect 195946 379256 209872 379284
rect 209866 379244 209872 379256
rect 209924 379284 209930 379296
rect 215266 379284 215294 379324
rect 219618 379312 219624 379364
rect 219676 379352 219682 379364
rect 273254 379352 273260 379364
rect 219676 379324 273260 379352
rect 219676 379312 219682 379324
rect 273254 379312 273260 379324
rect 273312 379312 273318 379364
rect 295334 379312 295340 379364
rect 295392 379352 295398 379364
rect 310974 379352 310980 379364
rect 295392 379324 310980 379352
rect 295392 379312 295398 379324
rect 310974 379312 310980 379324
rect 311032 379312 311038 379364
rect 218330 379284 218336 379296
rect 209924 379256 213040 379284
rect 215266 379256 218336 379284
rect 209924 379244 209930 379256
rect 91370 379176 91376 379228
rect 91428 379216 91434 379228
rect 211338 379216 211344 379228
rect 91428 379188 211344 379216
rect 91428 379176 91434 379188
rect 211338 379176 211344 379188
rect 211396 379216 211402 379228
rect 213012 379216 213040 379256
rect 218330 379244 218336 379256
rect 218388 379284 218394 379296
rect 271046 379284 271052 379296
rect 218388 379256 271052 379284
rect 218388 379244 218394 379256
rect 271046 379244 271052 379256
rect 271104 379244 271110 379296
rect 219526 379216 219532 379228
rect 211396 379188 212948 379216
rect 213012 379188 219532 379216
rect 211396 379176 211402 379188
rect 59722 379108 59728 379160
rect 59780 379148 59786 379160
rect 93486 379148 93492 379160
rect 59780 379120 93492 379148
rect 59780 379108 59786 379120
rect 93486 379108 93492 379120
rect 93544 379108 93550 379160
rect 93578 379108 93584 379160
rect 93636 379148 93642 379160
rect 201402 379148 201408 379160
rect 93636 379120 201408 379148
rect 93636 379108 93642 379120
rect 201402 379108 201408 379120
rect 201460 379108 201466 379160
rect 46290 379040 46296 379092
rect 46348 379080 46354 379092
rect 108206 379080 108212 379092
rect 46348 379052 108212 379080
rect 46348 379040 46354 379052
rect 108206 379040 108212 379052
rect 108264 379040 108270 379092
rect 108850 379040 108856 379092
rect 108908 379080 108914 379092
rect 205450 379080 205456 379092
rect 108908 379052 205456 379080
rect 108908 379040 108914 379052
rect 205450 379040 205456 379052
rect 205508 379080 205514 379092
rect 210326 379080 210332 379092
rect 205508 379052 210332 379080
rect 205508 379040 205514 379052
rect 210326 379040 210332 379052
rect 210384 379040 210390 379092
rect 212920 379080 212948 379188
rect 219526 379176 219532 379188
rect 219584 379216 219590 379228
rect 220170 379216 220176 379228
rect 219584 379188 220176 379216
rect 219584 379176 219590 379188
rect 220170 379176 220176 379188
rect 220228 379176 220234 379228
rect 220998 379080 221004 379092
rect 212920 379052 221004 379080
rect 220998 379040 221004 379052
rect 221056 379040 221062 379092
rect 373810 379040 373816 379092
rect 373868 379080 373874 379092
rect 380894 379080 380900 379092
rect 373868 379052 380900 379080
rect 373868 379040 373874 379052
rect 380894 379040 380900 379052
rect 380952 379040 380958 379092
rect 42150 378972 42156 379024
rect 42208 379012 42214 379024
rect 101030 379012 101036 379024
rect 42208 378984 101036 379012
rect 42208 378972 42214 378984
rect 101030 378972 101036 378984
rect 101088 378972 101094 379024
rect 112346 378972 112352 379024
rect 112404 379012 112410 379024
rect 206830 379012 206836 379024
rect 112404 378984 206836 379012
rect 112404 378972 112410 378984
rect 206830 378972 206836 378984
rect 206888 379012 206894 379024
rect 212350 379012 212356 379024
rect 206888 378984 212356 379012
rect 206888 378972 206894 378984
rect 212350 378972 212356 378984
rect 212408 379012 212414 379024
rect 272150 379012 272156 379024
rect 212408 378984 272156 379012
rect 212408 378972 212414 378984
rect 272150 378972 272156 378984
rect 272208 378972 272214 379024
rect 379790 378972 379796 379024
rect 379848 379012 379854 379024
rect 379974 379012 379980 379024
rect 379848 378984 379980 379012
rect 379848 378972 379854 378984
rect 379974 378972 379980 378984
rect 380032 379012 380038 379024
rect 397086 379012 397092 379024
rect 380032 378984 397092 379012
rect 380032 378972 380038 378984
rect 397086 378972 397092 378984
rect 397144 378972 397150 379024
rect 55674 378904 55680 378956
rect 55732 378944 55738 378956
rect 103514 378944 103520 378956
rect 55732 378916 103520 378944
rect 55732 378904 55738 378916
rect 103514 378904 103520 378916
rect 103572 378904 103578 378956
rect 201402 378904 201408 378956
rect 201460 378944 201466 378956
rect 220906 378944 220912 378956
rect 201460 378916 220912 378944
rect 201460 378904 201466 378916
rect 220906 378904 220912 378916
rect 220964 378904 220970 378956
rect 371142 378904 371148 378956
rect 371200 378944 371206 378956
rect 379514 378944 379520 378956
rect 371200 378916 379520 378944
rect 371200 378904 371206 378916
rect 379514 378904 379520 378916
rect 379572 378904 379578 378956
rect 57054 378836 57060 378888
rect 57112 378876 57118 378888
rect 104894 378876 104900 378888
rect 57112 378848 104900 378876
rect 57112 378836 57118 378848
rect 104894 378836 104900 378848
rect 104952 378836 104958 378888
rect 205634 378836 205640 378888
rect 205692 378876 205698 378888
rect 206830 378876 206836 378888
rect 205692 378848 206836 378876
rect 205692 378836 205698 378848
rect 206830 378836 206836 378848
rect 206888 378876 206894 378888
rect 219434 378876 219440 378888
rect 206888 378848 219440 378876
rect 206888 378836 206894 378848
rect 219434 378836 219440 378848
rect 219492 378836 219498 378888
rect 220722 378836 220728 378888
rect 220780 378876 220786 378888
rect 247586 378876 247592 378888
rect 220780 378848 247592 378876
rect 220780 378836 220786 378848
rect 247586 378836 247592 378848
rect 247644 378836 247650 378888
rect 376570 378836 376576 378888
rect 376628 378876 376634 378888
rect 396074 378876 396080 378888
rect 376628 378848 396080 378876
rect 376628 378836 376634 378848
rect 396074 378836 396080 378848
rect 396132 378836 396138 378888
rect 55766 378768 55772 378820
rect 55824 378808 55830 378820
rect 56962 378808 56968 378820
rect 55824 378780 56968 378808
rect 55824 378768 55830 378780
rect 56962 378768 56968 378780
rect 57020 378768 57026 378820
rect 222010 378768 222016 378820
rect 222068 378808 222074 378820
rect 245378 378808 245384 378820
rect 222068 378780 245384 378808
rect 222068 378768 222074 378780
rect 245378 378768 245384 378780
rect 245436 378768 245442 378820
rect 358722 378768 358728 378820
rect 358780 378808 358786 378820
rect 372614 378808 372620 378820
rect 358780 378780 372620 378808
rect 358780 378768 358786 378780
rect 372614 378768 372620 378780
rect 372672 378768 372678 378820
rect 377398 378768 377404 378820
rect 377456 378808 377462 378820
rect 437842 378808 437848 378820
rect 377456 378780 437848 378808
rect 377456 378768 377462 378780
rect 437842 378768 437848 378780
rect 437900 378768 437906 378820
rect 50062 378700 50068 378752
rect 50120 378740 50126 378752
rect 98454 378740 98460 378752
rect 50120 378712 98460 378740
rect 50120 378700 50126 378712
rect 98454 378700 98460 378712
rect 98512 378700 98518 378752
rect 211062 378700 211068 378752
rect 211120 378740 211126 378752
rect 219710 378740 219716 378752
rect 211120 378712 219716 378740
rect 211120 378700 211126 378712
rect 219710 378700 219716 378712
rect 219768 378740 219774 378752
rect 219768 378712 220032 378740
rect 219768 378700 219774 378712
rect 49050 378632 49056 378684
rect 49108 378672 49114 378684
rect 96062 378672 96068 378684
rect 49108 378644 96068 378672
rect 49108 378632 49114 378644
rect 96062 378632 96068 378644
rect 96120 378632 96126 378684
rect 46198 378564 46204 378616
rect 46256 378604 46262 378616
rect 47670 378604 47676 378616
rect 46256 378576 47676 378604
rect 46256 378564 46262 378576
rect 47670 378564 47676 378576
rect 47728 378564 47734 378616
rect 113450 378564 113456 378616
rect 113508 378604 113514 378616
rect 214190 378604 214196 378616
rect 113508 378576 214196 378604
rect 113508 378564 113514 378576
rect 214190 378564 214196 378576
rect 214248 378604 214254 378616
rect 219618 378604 219624 378616
rect 214248 378576 219624 378604
rect 214248 378564 214254 378576
rect 219618 378564 219624 378576
rect 219676 378564 219682 378616
rect 220004 378604 220032 378712
rect 375282 378700 375288 378752
rect 375340 378740 375346 378752
rect 400398 378740 400404 378752
rect 375340 378712 400404 378740
rect 375340 378700 375346 378712
rect 400398 378700 400404 378712
rect 400456 378700 400462 378752
rect 220170 378632 220176 378684
rect 220228 378672 220234 378684
rect 248598 378672 248604 378684
rect 220228 378644 248604 378672
rect 220228 378632 220234 378644
rect 248598 378632 248604 378644
rect 248656 378632 248662 378684
rect 372706 378632 372712 378684
rect 372764 378672 372770 378684
rect 373166 378672 373172 378684
rect 372764 378644 373172 378672
rect 372764 378632 372770 378644
rect 373166 378632 373172 378644
rect 373224 378672 373230 378684
rect 399478 378672 399484 378684
rect 373224 378644 399484 378672
rect 373224 378632 373230 378644
rect 399478 378632 399484 378644
rect 399536 378632 399542 378684
rect 250070 378604 250076 378616
rect 220004 378576 250076 378604
rect 250070 378564 250076 378576
rect 250128 378564 250134 378616
rect 379330 378564 379336 378616
rect 379388 378604 379394 378616
rect 379882 378604 379888 378616
rect 379388 378576 379888 378604
rect 379388 378564 379394 378576
rect 379882 378564 379888 378576
rect 379940 378604 379946 378616
rect 405826 378604 405832 378616
rect 379940 378576 405832 378604
rect 379940 378564 379946 378576
rect 405826 378564 405832 378576
rect 405884 378564 405890 378616
rect 114462 378496 114468 378548
rect 114520 378536 114526 378548
rect 205634 378536 205640 378548
rect 114520 378508 205640 378536
rect 114520 378496 114526 378508
rect 205634 378496 205640 378508
rect 205692 378496 205698 378548
rect 213822 378496 213828 378548
rect 213880 378536 213886 378548
rect 213880 378508 220400 378536
rect 213880 378496 213886 378508
rect 115842 378428 115848 378480
rect 115900 378468 115906 378480
rect 213362 378468 213368 378480
rect 115900 378440 213368 378468
rect 115900 378428 115906 378440
rect 213362 378428 213368 378440
rect 213420 378468 213426 378480
rect 220078 378468 220084 378480
rect 213420 378440 220084 378468
rect 213420 378428 213426 378440
rect 220078 378428 220084 378440
rect 220136 378428 220142 378480
rect 220372 378468 220400 378508
rect 220998 378496 221004 378548
rect 221056 378536 221062 378548
rect 251174 378536 251180 378548
rect 221056 378508 251180 378536
rect 221056 378496 221062 378508
rect 251174 378496 251180 378508
rect 251232 378496 251238 378548
rect 380894 378496 380900 378548
rect 380952 378536 380958 378548
rect 381170 378536 381176 378548
rect 380952 378508 381176 378536
rect 380952 378496 380958 378508
rect 381170 378496 381176 378508
rect 381228 378536 381234 378548
rect 412358 378536 412364 378548
rect 381228 378508 412364 378536
rect 381228 378496 381234 378508
rect 412358 378496 412364 378508
rect 412416 378496 412422 378548
rect 220814 378468 220820 378480
rect 220372 378440 220820 378468
rect 220814 378428 220820 378440
rect 220872 378468 220878 378480
rect 252278 378468 252284 378480
rect 220872 378440 252284 378468
rect 220872 378428 220878 378440
rect 252278 378428 252284 378440
rect 252336 378428 252342 378480
rect 379514 378428 379520 378480
rect 379572 378468 379578 378480
rect 411254 378468 411260 378480
rect 379572 378440 411260 378468
rect 379572 378428 379578 378440
rect 411254 378428 411260 378440
rect 411312 378428 411318 378480
rect 111334 378360 111340 378412
rect 111392 378400 111398 378412
rect 208486 378400 208492 378412
rect 111392 378372 208492 378400
rect 111392 378360 111398 378372
rect 208486 378360 208492 378372
rect 208544 378360 208550 378412
rect 210326 378360 210332 378412
rect 210384 378400 210390 378412
rect 268654 378400 268660 378412
rect 210384 378372 268660 378400
rect 210384 378360 210390 378372
rect 268654 378360 268660 378372
rect 268712 378360 268718 378412
rect 372614 378360 372620 378412
rect 372672 378400 372678 378412
rect 373902 378400 373908 378412
rect 372672 378372 373908 378400
rect 372672 378360 372678 378372
rect 373902 378360 373908 378372
rect 373960 378400 373966 378412
rect 407574 378400 407580 378412
rect 373960 378372 407580 378400
rect 373960 378360 373966 378372
rect 407574 378360 407580 378372
rect 407632 378360 407638 378412
rect 90082 378292 90088 378344
rect 90140 378332 90146 378344
rect 209774 378332 209780 378344
rect 90140 378304 209780 378332
rect 90140 378292 90146 378304
rect 209774 378292 209780 378304
rect 209832 378332 209838 378344
rect 211062 378332 211068 378344
rect 209832 378304 211068 378332
rect 209832 378292 209838 378304
rect 211062 378292 211068 378304
rect 211120 378292 211126 378344
rect 211706 378292 211712 378344
rect 211764 378332 211770 378344
rect 212442 378332 212448 378344
rect 211764 378304 212448 378332
rect 211764 378292 211770 378304
rect 212442 378292 212448 378304
rect 212500 378332 212506 378344
rect 246206 378332 246212 378344
rect 212500 378304 246212 378332
rect 212500 378292 212506 378304
rect 246206 378292 246212 378304
rect 246264 378292 246270 378344
rect 273254 378292 273260 378344
rect 273312 378332 273318 378344
rect 300854 378332 300860 378344
rect 273312 378304 300860 378332
rect 273312 378292 273318 378304
rect 300854 378292 300860 378304
rect 300912 378292 300918 378344
rect 342254 378292 342260 378344
rect 342312 378332 342318 378344
rect 343174 378332 343180 378344
rect 342312 378304 343180 378332
rect 342312 378292 342318 378304
rect 343174 378292 343180 378304
rect 343232 378332 343238 378344
rect 360194 378332 360200 378344
rect 343232 378304 360200 378332
rect 343232 378292 343238 378304
rect 360194 378292 360200 378304
rect 360252 378332 360258 378344
rect 360252 378304 364334 378332
rect 360252 378292 360258 378304
rect 85482 378224 85488 378276
rect 85540 378264 85546 378276
rect 208578 378264 208584 378276
rect 85540 378236 208584 378264
rect 85540 378224 85546 378236
rect 208578 378224 208584 378236
rect 208636 378264 208642 378276
rect 212994 378264 213000 378276
rect 208636 378236 213000 378264
rect 208636 378224 208642 378236
rect 212994 378224 213000 378236
rect 213052 378264 213058 378276
rect 213638 378264 213644 378276
rect 213052 378236 213644 378264
rect 213052 378224 213058 378236
rect 213638 378224 213644 378236
rect 213696 378224 213702 378276
rect 276014 378224 276020 378276
rect 276072 378264 276078 378276
rect 277026 378264 277032 378276
rect 276072 378236 277032 378264
rect 276072 378224 276078 378236
rect 277026 378224 277032 378236
rect 277084 378264 277090 378276
rect 356606 378264 356612 378276
rect 277084 378236 356612 378264
rect 277084 378224 277090 378236
rect 356606 378224 356612 378236
rect 356664 378224 356670 378276
rect 364306 378264 364334 378304
rect 375374 378292 375380 378344
rect 375432 378332 375438 378344
rect 435174 378332 435180 378344
rect 375432 378304 435180 378332
rect 375432 378292 375438 378304
rect 435174 378292 435180 378304
rect 435232 378292 435238 378344
rect 503070 378264 503076 378276
rect 364306 378236 503076 378264
rect 503070 378224 503076 378236
rect 503128 378264 503134 378276
rect 517606 378264 517612 378276
rect 503128 378236 517612 378264
rect 503128 378224 503134 378236
rect 517606 378224 517612 378236
rect 517664 378264 517670 378276
rect 580258 378264 580264 378276
rect 517664 378236 580264 378264
rect 517664 378224 517670 378236
rect 580258 378224 580264 378236
rect 580316 378224 580322 378276
rect 47670 378156 47676 378208
rect 47728 378196 47734 378208
rect 80422 378196 80428 378208
rect 47728 378168 80428 378196
rect 47728 378156 47734 378168
rect 80422 378156 80428 378168
rect 80480 378156 80486 378208
rect 87874 378156 87880 378208
rect 87932 378196 87938 378208
rect 219618 378196 219624 378208
rect 87932 378168 219624 378196
rect 87932 378156 87938 378168
rect 219618 378156 219624 378168
rect 219676 378196 219682 378208
rect 220722 378196 220728 378208
rect 219676 378168 220728 378196
rect 219676 378156 219682 378168
rect 220722 378156 220728 378168
rect 220780 378156 220786 378208
rect 220906 378156 220912 378208
rect 220964 378196 220970 378208
rect 221182 378196 221188 378208
rect 220964 378168 221188 378196
rect 220964 378156 220970 378168
rect 221182 378156 221188 378168
rect 221240 378196 221246 378208
rect 253382 378196 253388 378208
rect 221240 378168 253388 378196
rect 221240 378156 221246 378168
rect 253382 378156 253388 378168
rect 253440 378156 253446 378208
rect 271782 378156 271788 378208
rect 271840 378196 271846 378208
rect 305822 378196 305828 378208
rect 271840 378168 305828 378196
rect 271840 378156 271846 378168
rect 305822 378156 305828 378168
rect 305880 378156 305886 378208
rect 343542 378156 343548 378208
rect 343600 378196 343606 378208
rect 503530 378196 503536 378208
rect 343600 378168 503536 378196
rect 343600 378156 343606 378168
rect 503530 378156 503536 378168
rect 503588 378196 503594 378208
rect 517698 378196 517704 378208
rect 503588 378168 517704 378196
rect 503588 378156 503594 378168
rect 517698 378156 517704 378168
rect 517756 378196 517762 378208
rect 580166 378196 580172 378208
rect 517756 378168 580172 378196
rect 517756 378156 517762 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 196710 378088 196716 378140
rect 196768 378128 196774 378140
rect 287606 378128 287612 378140
rect 196768 378100 287612 378128
rect 196768 378088 196774 378100
rect 287606 378088 287612 378100
rect 287664 378088 287670 378140
rect 372338 378088 372344 378140
rect 372396 378128 372402 378140
rect 474826 378128 474832 378140
rect 372396 378100 474832 378128
rect 372396 378088 372402 378100
rect 474826 378088 474832 378100
rect 474884 378088 474890 378140
rect 42058 378020 42064 378072
rect 42116 378060 42122 378072
rect 199470 378060 199476 378072
rect 42116 378032 199476 378060
rect 42116 378020 42122 378032
rect 199470 378020 199476 378032
rect 199528 378020 199534 378072
rect 203978 378020 203984 378072
rect 204036 378060 204042 378072
rect 317414 378060 317420 378072
rect 204036 378032 317420 378060
rect 204036 378020 204042 378032
rect 317414 378020 317420 378032
rect 317472 378020 317478 378072
rect 364242 378020 364248 378072
rect 364300 378060 364306 378072
rect 375282 378060 375288 378072
rect 364300 378032 375288 378060
rect 364300 378020 364306 378032
rect 375282 378020 375288 378032
rect 375340 378020 375346 378072
rect 375834 378020 375840 378072
rect 375892 378060 375898 378072
rect 460934 378060 460940 378072
rect 375892 378032 460940 378060
rect 375892 378020 375898 378032
rect 460934 378020 460940 378032
rect 460992 378020 460998 378072
rect 197446 377952 197452 378004
rect 197504 377992 197510 378004
rect 298462 377992 298468 378004
rect 197504 377964 298468 377992
rect 197504 377952 197510 377964
rect 298462 377952 298468 377964
rect 298520 377952 298526 378004
rect 374454 377952 374460 378004
rect 374512 377992 374518 378004
rect 458358 377992 458364 378004
rect 374512 377964 458364 377992
rect 374512 377952 374518 377964
rect 458358 377952 458364 377964
rect 458416 377952 458422 378004
rect 54386 377884 54392 377936
rect 54444 377924 54450 377936
rect 183462 377924 183468 377936
rect 54444 377896 183468 377924
rect 54444 377884 54450 377896
rect 183462 377884 183468 377896
rect 183520 377884 183526 377936
rect 197630 377884 197636 377936
rect 197688 377924 197694 377936
rect 295426 377924 295432 377936
rect 197688 377896 295432 377924
rect 197688 377884 197694 377896
rect 295426 377884 295432 377896
rect 295484 377884 295490 377936
rect 362862 377884 362868 377936
rect 362920 377924 362926 377936
rect 445846 377924 445852 377936
rect 362920 377896 445852 377924
rect 362920 377884 362926 377896
rect 445846 377884 445852 377896
rect 445904 377884 445910 377936
rect 54294 377816 54300 377868
rect 54352 377856 54358 377868
rect 182266 377856 182272 377868
rect 54352 377828 182272 377856
rect 54352 377816 54358 377828
rect 182266 377816 182272 377828
rect 182324 377856 182330 377868
rect 182818 377856 182824 377868
rect 182324 377828 182824 377856
rect 182324 377816 182330 377828
rect 182818 377816 182824 377828
rect 182876 377816 182882 377868
rect 197538 377816 197544 377868
rect 197596 377856 197602 377868
rect 292666 377856 292672 377868
rect 197596 377828 292672 377856
rect 197596 377816 197602 377828
rect 292666 377816 292672 377828
rect 292724 377816 292730 377868
rect 367554 377816 367560 377868
rect 367612 377856 367618 377868
rect 450998 377856 451004 377868
rect 367612 377828 451004 377856
rect 367612 377816 367618 377828
rect 450998 377816 451004 377828
rect 451056 377816 451062 377868
rect 95970 377748 95976 377800
rect 96028 377788 96034 377800
rect 212534 377788 212540 377800
rect 96028 377760 212540 377788
rect 96028 377748 96034 377760
rect 212534 377748 212540 377760
rect 212592 377788 212598 377800
rect 213270 377788 213276 377800
rect 212592 377760 213276 377788
rect 212592 377748 212598 377760
rect 213270 377748 213276 377760
rect 213328 377748 213334 377800
rect 215754 377788 215760 377800
rect 214852 377760 215760 377788
rect 98270 377680 98276 377732
rect 98328 377720 98334 377732
rect 212626 377720 212632 377732
rect 98328 377692 212632 377720
rect 98328 377680 98334 377692
rect 212626 377680 212632 377692
rect 212684 377720 212690 377732
rect 214852 377720 214880 377760
rect 215754 377748 215760 377760
rect 215812 377748 215818 377800
rect 217410 377748 217416 377800
rect 217468 377788 217474 377800
rect 307846 377788 307852 377800
rect 217468 377760 307852 377788
rect 217468 377748 217474 377760
rect 307846 377748 307852 377760
rect 307904 377748 307910 377800
rect 370406 377748 370412 377800
rect 370464 377788 370470 377800
rect 453022 377788 453028 377800
rect 370464 377760 453028 377788
rect 370464 377748 370470 377760
rect 453022 377748 453028 377760
rect 453080 377748 453086 377800
rect 212684 377692 214880 377720
rect 212684 377680 212690 377692
rect 214926 377680 214932 377732
rect 214984 377720 214990 377732
rect 303246 377720 303252 377732
rect 214984 377692 303252 377720
rect 214984 377680 214990 377692
rect 303246 377680 303252 377692
rect 303304 377680 303310 377732
rect 373718 377680 373724 377732
rect 373776 377720 373782 377732
rect 455506 377720 455512 377732
rect 373776 377692 455512 377720
rect 373776 377680 373782 377692
rect 455506 377680 455512 377692
rect 455564 377680 455570 377732
rect 196802 377612 196808 377664
rect 196860 377652 196866 377664
rect 290918 377652 290924 377664
rect 196860 377624 290924 377652
rect 196860 377612 196866 377624
rect 290918 377612 290924 377624
rect 290976 377612 290982 377664
rect 365530 377612 365536 377664
rect 365588 377652 365594 377664
rect 447502 377652 447508 377664
rect 365588 377624 447508 377652
rect 365588 377612 365594 377624
rect 447502 377612 447508 377624
rect 447560 377612 447566 377664
rect 196618 377544 196624 377596
rect 196676 377584 196682 377596
rect 285950 377584 285956 377596
rect 196676 377556 285956 377584
rect 196676 377544 196682 377556
rect 285950 377544 285956 377556
rect 286008 377544 286014 377596
rect 358538 377544 358544 377596
rect 358596 377584 358602 377596
rect 425974 377584 425980 377596
rect 358596 377556 425980 377584
rect 358596 377544 358602 377556
rect 425974 377544 425980 377556
rect 426032 377544 426038 377596
rect 197078 377476 197084 377528
rect 197136 377516 197142 377528
rect 278222 377516 278228 377528
rect 197136 377488 278228 377516
rect 197136 377476 197142 377488
rect 278222 377476 278228 377488
rect 278280 377476 278286 377528
rect 361390 377476 361396 377528
rect 361448 377516 361454 377528
rect 415670 377516 415676 377528
rect 361448 377488 415676 377516
rect 361448 377476 361454 377488
rect 415670 377476 415676 377488
rect 415728 377476 415734 377528
rect 43346 377408 43352 377460
rect 43404 377448 43410 377460
rect 199562 377448 199568 377460
rect 43404 377420 199568 377448
rect 43404 377408 43410 377420
rect 199562 377408 199568 377420
rect 199620 377408 199626 377460
rect 199746 377408 199752 377460
rect 199804 377448 199810 377460
rect 273254 377448 273260 377460
rect 199804 377420 273260 377448
rect 199804 377408 199810 377420
rect 273254 377408 273260 377420
rect 273312 377408 273318 377460
rect 360746 377408 360752 377460
rect 360804 377448 360810 377460
rect 360804 377420 373994 377448
rect 360804 377408 360810 377420
rect 150986 377340 150992 377392
rect 151044 377380 151050 377392
rect 198182 377380 198188 377392
rect 151044 377352 198188 377380
rect 151044 377340 151050 377352
rect 198182 377340 198188 377352
rect 198240 377340 198246 377392
rect 198734 377340 198740 377392
rect 198792 377380 198798 377392
rect 271782 377380 271788 377392
rect 198792 377352 271788 377380
rect 198792 377340 198798 377352
rect 271782 377340 271788 377352
rect 271840 377340 271846 377392
rect 373966 377380 373994 377420
rect 376662 377408 376668 377460
rect 376720 377448 376726 377460
rect 416866 377448 416872 377460
rect 376720 377420 416872 377448
rect 376720 377408 376726 377420
rect 416866 377408 416872 377420
rect 416924 377408 416930 377460
rect 375190 377380 375196 377392
rect 373966 377352 375196 377380
rect 375190 377340 375196 377352
rect 375248 377380 375254 377392
rect 415854 377380 415860 377392
rect 375248 377352 415860 377380
rect 375248 377340 375254 377352
rect 415854 377340 415860 377352
rect 415912 377340 415918 377392
rect 138474 377272 138480 377324
rect 138532 377312 138538 377324
rect 207290 377312 207296 377324
rect 138532 377284 207296 377312
rect 138532 377272 138538 377284
rect 207290 377272 207296 377284
rect 207348 377272 207354 377324
rect 211614 377272 211620 377324
rect 211672 377312 211678 377324
rect 280246 377312 280252 377324
rect 211672 377284 280252 377312
rect 211672 377272 211678 377284
rect 280246 377272 280252 377284
rect 280304 377272 280310 377324
rect 364794 377272 364800 377324
rect 364852 377312 364858 377324
rect 379330 377312 379336 377324
rect 364852 377284 379336 377312
rect 364852 377272 364858 377284
rect 379330 377272 379336 377284
rect 379388 377312 379394 377324
rect 409966 377312 409972 377324
rect 379388 377284 409972 377312
rect 379388 377272 379394 377284
rect 409966 377272 409972 377284
rect 410024 377272 410030 377324
rect 48866 377204 48872 377256
rect 48924 377244 48930 377256
rect 216766 377244 216772 377256
rect 48924 377216 216772 377244
rect 48924 377204 48930 377216
rect 216766 377204 216772 377216
rect 216824 377244 216830 377256
rect 216950 377244 216956 377256
rect 216824 377216 216956 377244
rect 216824 377204 216830 377216
rect 216950 377204 216956 377216
rect 217008 377204 217014 377256
rect 374546 377204 374552 377256
rect 374604 377244 374610 377256
rect 375282 377244 375288 377256
rect 374604 377216 375288 377244
rect 374604 377204 374610 377216
rect 375282 377204 375288 377216
rect 375340 377244 375346 377256
rect 402974 377244 402980 377256
rect 375340 377216 402980 377244
rect 375340 377204 375346 377216
rect 402974 377204 402980 377216
rect 403032 377204 403038 377256
rect 154022 377136 154028 377188
rect 154080 377176 154086 377188
rect 200390 377176 200396 377188
rect 154080 377148 200396 377176
rect 154080 377136 154086 377148
rect 200390 377136 200396 377148
rect 200448 377136 200454 377188
rect 212994 377136 213000 377188
rect 213052 377176 213058 377188
rect 213546 377176 213552 377188
rect 213052 377148 213552 377176
rect 213052 377136 213058 377148
rect 213546 377136 213552 377148
rect 213604 377136 213610 377188
rect 362126 377136 362132 377188
rect 362184 377176 362190 377188
rect 375926 377176 375932 377188
rect 362184 377148 375932 377176
rect 362184 377136 362190 377148
rect 375926 377136 375932 377148
rect 375984 377176 375990 377188
rect 376662 377176 376668 377188
rect 375984 377148 376668 377176
rect 375984 377136 375990 377148
rect 376662 377136 376668 377148
rect 376720 377136 376726 377188
rect 380986 377136 380992 377188
rect 381044 377176 381050 377188
rect 381354 377176 381360 377188
rect 381044 377148 381360 377176
rect 381044 377136 381050 377148
rect 381354 377136 381360 377148
rect 381412 377136 381418 377188
rect 374454 377068 374460 377120
rect 374512 377108 374518 377120
rect 375282 377108 375288 377120
rect 374512 377080 375288 377108
rect 374512 377068 374518 377080
rect 375282 377068 375288 377080
rect 375340 377068 375346 377120
rect 376478 377000 376484 377052
rect 376536 377040 376542 377052
rect 376662 377040 376668 377052
rect 376536 377012 376668 377040
rect 376536 377000 376542 377012
rect 376662 377000 376668 377012
rect 376720 377000 376726 377052
rect 375374 376864 375380 376916
rect 375432 376904 375438 376916
rect 376478 376904 376484 376916
rect 375432 376876 376484 376904
rect 375432 376864 375438 376876
rect 376478 376864 376484 376876
rect 376536 376864 376542 376916
rect 368382 376728 368388 376780
rect 368440 376768 368446 376780
rect 372614 376768 372620 376780
rect 368440 376740 372620 376768
rect 368440 376728 368446 376740
rect 372614 376728 372620 376740
rect 372672 376728 372678 376780
rect 77202 376660 77208 376712
rect 77260 376700 77266 376712
rect 204346 376700 204352 376712
rect 77260 376672 204352 376700
rect 77260 376660 77266 376672
rect 204346 376660 204352 376672
rect 204404 376700 204410 376712
rect 215846 376700 215852 376712
rect 204404 376672 215852 376700
rect 204404 376660 204410 376672
rect 215846 376660 215852 376672
rect 215904 376660 215910 376712
rect 362770 376660 362776 376712
rect 362828 376700 362834 376712
rect 477586 376700 477592 376712
rect 362828 376672 477592 376700
rect 362828 376660 362834 376672
rect 477586 376660 477592 376672
rect 477644 376660 477650 376712
rect 206646 376592 206652 376644
rect 206704 376632 206710 376644
rect 283374 376632 283380 376644
rect 206704 376604 283380 376632
rect 206704 376592 206710 376604
rect 283374 376592 283380 376604
rect 283432 376592 283438 376644
rect 369670 376592 369676 376644
rect 369728 376632 369734 376644
rect 483382 376632 483388 376644
rect 369728 376604 483388 376632
rect 369728 376592 369734 376604
rect 483382 376592 483388 376604
rect 483440 376592 483446 376644
rect 135898 376524 135904 376576
rect 135956 376564 135962 376576
rect 200298 376564 200304 376576
rect 135956 376536 200304 376564
rect 135956 376524 135962 376536
rect 200298 376524 200304 376536
rect 200356 376524 200362 376576
rect 201586 376524 201592 376576
rect 201644 376564 201650 376576
rect 320910 376564 320916 376576
rect 201644 376536 320916 376564
rect 201644 376524 201650 376536
rect 320910 376524 320916 376536
rect 320968 376524 320974 376576
rect 365622 376524 365628 376576
rect 365680 376564 365686 376576
rect 473446 376564 473452 376576
rect 365680 376536 473452 376564
rect 365680 376524 365686 376536
rect 473446 376524 473452 376536
rect 473504 376524 473510 376576
rect 94682 376456 94688 376508
rect 94740 376496 94746 376508
rect 212718 376496 212724 376508
rect 94740 376468 212724 376496
rect 94740 376456 94746 376468
rect 212718 376456 212724 376468
rect 212776 376456 212782 376508
rect 214282 376456 214288 376508
rect 214340 376496 214346 376508
rect 276106 376496 276112 376508
rect 214340 376468 276112 376496
rect 214340 376456 214346 376468
rect 276106 376456 276112 376468
rect 276164 376456 276170 376508
rect 358630 376456 358636 376508
rect 358688 376496 358694 376508
rect 463510 376496 463516 376508
rect 358688 376468 463516 376496
rect 358688 376456 358694 376468
rect 463510 376456 463516 376468
rect 463568 376456 463574 376508
rect 83274 376388 83280 376440
rect 83332 376428 83338 376440
rect 207106 376428 207112 376440
rect 83332 376400 207112 376428
rect 83332 376388 83338 376400
rect 207106 376388 207112 376400
rect 207164 376388 207170 376440
rect 213086 376388 213092 376440
rect 213144 376428 213150 376440
rect 273438 376428 273444 376440
rect 213144 376400 273444 376428
rect 213144 376388 213150 376400
rect 273438 376388 273444 376400
rect 273496 376388 273502 376440
rect 368290 376388 368296 376440
rect 368348 376428 368354 376440
rect 470778 376428 470784 376440
rect 368348 376400 470784 376428
rect 368348 376388 368354 376400
rect 470778 376388 470784 376400
rect 470836 376388 470842 376440
rect 99466 376320 99472 376372
rect 99524 376360 99530 376372
rect 214006 376360 214012 376372
rect 99524 376332 214012 376360
rect 99524 376320 99530 376332
rect 214006 376320 214012 376332
rect 214064 376320 214070 376372
rect 216490 376320 216496 376372
rect 216548 376360 216554 376372
rect 270954 376360 270960 376372
rect 216548 376332 270960 376360
rect 216548 376320 216554 376332
rect 270954 376320 270960 376332
rect 271012 376320 271018 376372
rect 370222 376320 370228 376372
rect 370280 376360 370286 376372
rect 467926 376360 467932 376372
rect 370280 376332 467932 376360
rect 370280 376320 370286 376332
rect 467926 376320 467932 376332
rect 467984 376320 467990 376372
rect 148686 376252 148692 376304
rect 148744 376292 148750 376304
rect 196986 376292 196992 376304
rect 148744 376264 196992 376292
rect 148744 376252 148750 376264
rect 196986 376252 196992 376264
rect 197044 376252 197050 376304
rect 213454 376252 213460 376304
rect 213512 376292 213518 376304
rect 268102 376292 268108 376304
rect 213512 376264 268108 376292
rect 213512 376252 213518 376264
rect 268102 376252 268108 376264
rect 268160 376252 268166 376304
rect 366910 376252 366916 376304
rect 366968 376292 366974 376304
rect 430666 376292 430672 376304
rect 366968 376264 430672 376292
rect 366968 376252 366974 376264
rect 430666 376252 430672 376264
rect 430724 376252 430730 376304
rect 211522 376184 211528 376236
rect 211580 376224 211586 376236
rect 265894 376224 265900 376236
rect 211580 376196 265900 376224
rect 211580 376184 211586 376196
rect 265894 376184 265900 376196
rect 265952 376184 265958 376236
rect 372614 376184 372620 376236
rect 372672 376224 372678 376236
rect 436186 376224 436192 376236
rect 372672 376196 436192 376224
rect 372672 376184 372678 376196
rect 436186 376184 436192 376196
rect 436244 376184 436250 376236
rect 214374 376116 214380 376168
rect 214432 376156 214438 376168
rect 263594 376156 263600 376168
rect 214432 376128 263600 376156
rect 214432 376116 214438 376128
rect 263594 376116 263600 376128
rect 263652 376116 263658 376168
rect 374362 376116 374368 376168
rect 374420 376156 374426 376168
rect 422846 376156 422852 376168
rect 374420 376128 422852 376156
rect 374420 376116 374426 376128
rect 422846 376116 422852 376128
rect 422904 376116 422910 376168
rect 208026 376048 208032 376100
rect 208084 376088 208090 376100
rect 250622 376088 250628 376100
rect 208084 376060 250628 376088
rect 208084 376048 208090 376060
rect 250622 376048 250628 376060
rect 250680 376048 250686 376100
rect 366266 376048 366272 376100
rect 366324 376088 366330 376100
rect 413278 376088 413284 376100
rect 366324 376060 413284 376088
rect 366324 376048 366330 376060
rect 413278 376048 413284 376060
rect 413336 376048 413342 376100
rect 97810 375980 97816 376032
rect 97868 376020 97874 376032
rect 215018 376020 215024 376032
rect 97868 375992 215024 376020
rect 97868 375980 97874 375992
rect 215018 375980 215024 375992
rect 215076 376020 215082 376032
rect 215294 376020 215300 376032
rect 215076 375992 215300 376020
rect 215076 375980 215082 375992
rect 215294 375980 215300 375992
rect 215352 375980 215358 376032
rect 219250 375980 219256 376032
rect 219308 376020 219314 376032
rect 260926 376020 260932 376032
rect 219308 375992 260932 376020
rect 219308 375980 219314 375992
rect 260926 375980 260932 375992
rect 260984 375980 260990 376032
rect 377490 375980 377496 376032
rect 377548 376020 377554 376032
rect 418430 376020 418436 376032
rect 377548 375992 418436 376020
rect 377548 375980 377554 375992
rect 418430 375980 418436 375992
rect 418488 375980 418494 376032
rect 208946 375912 208952 375964
rect 209004 375952 209010 375964
rect 258350 375952 258356 375964
rect 209004 375924 258356 375952
rect 209004 375912 209010 375924
rect 258350 375912 258356 375924
rect 258408 375912 258414 375964
rect 357158 375912 357164 375964
rect 357216 375952 357222 375964
rect 379974 375952 379980 375964
rect 357216 375924 379980 375952
rect 357216 375912 357222 375924
rect 379974 375912 379980 375924
rect 380032 375952 380038 375964
rect 414566 375952 414572 375964
rect 380032 375924 414572 375952
rect 380032 375912 380038 375924
rect 414566 375912 414572 375924
rect 414624 375912 414630 375964
rect 100846 375844 100852 375896
rect 100904 375884 100910 375896
rect 214466 375884 214472 375896
rect 100904 375856 214472 375884
rect 100904 375844 100910 375856
rect 214466 375844 214472 375856
rect 214524 375844 214530 375896
rect 216398 375844 216404 375896
rect 216456 375884 216462 375896
rect 255958 375884 255964 375896
rect 216456 375856 255964 375884
rect 216456 375844 216462 375856
rect 255958 375844 255964 375856
rect 256016 375844 256022 375896
rect 217502 375776 217508 375828
rect 217560 375816 217566 375828
rect 253566 375816 253572 375828
rect 217560 375788 253572 375816
rect 217560 375776 217566 375788
rect 253566 375776 253572 375788
rect 253624 375776 253630 375828
rect 202874 375708 202880 375760
rect 202932 375748 202938 375760
rect 325878 375748 325884 375760
rect 202932 375720 325884 375748
rect 202932 375708 202938 375720
rect 325878 375708 325884 375720
rect 325936 375708 325942 375760
rect 105722 375640 105728 375692
rect 105780 375680 105786 375692
rect 218514 375680 218520 375692
rect 105780 375652 218520 375680
rect 105780 375640 105786 375652
rect 218514 375640 218520 375652
rect 218572 375680 218578 375692
rect 219342 375680 219348 375692
rect 218572 375652 219348 375680
rect 218572 375640 218578 375652
rect 219342 375640 219348 375652
rect 219400 375640 219406 375692
rect 372982 375368 372988 375420
rect 373040 375408 373046 375420
rect 376754 375408 376760 375420
rect 373040 375380 376760 375408
rect 373040 375368 373046 375380
rect 376754 375368 376760 375380
rect 376812 375408 376818 375420
rect 377398 375408 377404 375420
rect 376812 375380 377404 375408
rect 376812 375368 376818 375380
rect 377398 375368 377404 375380
rect 377456 375368 377462 375420
rect 84378 375300 84384 375352
rect 84436 375340 84442 375352
rect 208394 375340 208400 375352
rect 84436 375312 208400 375340
rect 84436 375300 84442 375312
rect 208394 375300 208400 375312
rect 208452 375340 208458 375352
rect 208670 375340 208676 375352
rect 208452 375312 208676 375340
rect 208452 375300 208458 375312
rect 208670 375300 208676 375312
rect 208728 375300 208734 375352
rect 215386 375340 215392 375352
rect 209746 375312 215392 375340
rect 102962 375232 102968 375284
rect 103020 375272 103026 375284
rect 209746 375272 209774 375312
rect 215386 375300 215392 375312
rect 215444 375340 215450 375352
rect 217226 375340 217232 375352
rect 215444 375312 217232 375340
rect 215444 375300 215450 375312
rect 217226 375300 217232 375312
rect 217284 375300 217290 375352
rect 372430 375300 372436 375352
rect 372488 375340 372494 375352
rect 379698 375340 379704 375352
rect 372488 375312 379704 375340
rect 372488 375300 372494 375312
rect 379698 375300 379704 375312
rect 379756 375340 379762 375352
rect 432230 375340 432236 375352
rect 379756 375312 432236 375340
rect 379756 375300 379762 375312
rect 432230 375300 432236 375312
rect 432288 375300 432294 375352
rect 103020 375244 209774 375272
rect 103020 375232 103026 375244
rect 213914 375232 213920 375284
rect 213972 375272 213978 375284
rect 216490 375272 216496 375284
rect 213972 375244 216496 375272
rect 213972 375232 213978 375244
rect 216490 375232 216496 375244
rect 216548 375232 216554 375284
rect 369762 375232 369768 375284
rect 369820 375272 369826 375284
rect 376754 375272 376760 375284
rect 369820 375244 376760 375272
rect 369820 375232 369826 375244
rect 376754 375232 376760 375244
rect 376812 375272 376818 375284
rect 425146 375272 425152 375284
rect 376812 375244 425152 375272
rect 376812 375232 376818 375244
rect 425146 375232 425152 375244
rect 425204 375232 425210 375284
rect 101858 375164 101864 375216
rect 101916 375204 101922 375216
rect 213932 375204 213960 375232
rect 101916 375176 213960 375204
rect 101916 375164 101922 375176
rect 375742 375164 375748 375216
rect 375800 375204 375806 375216
rect 421190 375204 421196 375216
rect 375800 375176 421196 375204
rect 375800 375164 375806 375176
rect 421190 375164 421196 375176
rect 421248 375164 421254 375216
rect 107562 375096 107568 375148
rect 107620 375136 107626 375148
rect 107620 375108 205634 375136
rect 107620 375096 107626 375108
rect 106458 375028 106464 375080
rect 106516 375068 106522 375080
rect 106516 375040 195974 375068
rect 106516 375028 106522 375040
rect 195946 374728 195974 375040
rect 205606 374796 205634 375108
rect 377398 375096 377404 375148
rect 377456 375136 377462 375148
rect 420638 375136 420644 375148
rect 377456 375108 420644 375136
rect 377456 375096 377462 375108
rect 420638 375096 420644 375108
rect 420696 375096 420702 375148
rect 367646 375028 367652 375080
rect 367704 375068 367710 375080
rect 377490 375068 377496 375080
rect 367704 375040 377496 375068
rect 367704 375028 367710 375040
rect 377490 375028 377496 375040
rect 377548 375068 377554 375080
rect 408678 375068 408684 375080
rect 377548 375040 408684 375068
rect 377548 375028 377554 375040
rect 408678 375028 408684 375040
rect 408736 375028 408742 375080
rect 216398 375000 216404 375012
rect 215266 374972 216404 375000
rect 208394 374824 208400 374876
rect 208452 374864 208458 374876
rect 215266 374864 215294 374972
rect 216398 374960 216404 374972
rect 216456 375000 216462 375012
rect 244274 375000 244280 375012
rect 216456 374972 244280 375000
rect 216456 374960 216462 374972
rect 244274 374960 244280 374972
rect 244332 374960 244338 375012
rect 377122 375000 377128 375012
rect 373966 374972 377128 375000
rect 216490 374892 216496 374944
rect 216548 374932 216554 374944
rect 261662 374932 261668 374944
rect 216548 374904 261668 374932
rect 216548 374892 216554 374904
rect 261662 374892 261668 374904
rect 261720 374892 261726 374944
rect 364886 374892 364892 374944
rect 364944 374932 364950 374944
rect 373966 374932 373994 374972
rect 377122 374960 377128 374972
rect 377180 375000 377186 375012
rect 418154 375000 418160 375012
rect 377180 374972 418160 375000
rect 377180 374960 377186 374972
rect 418154 374960 418160 374972
rect 418212 374960 418218 375012
rect 364944 374904 373994 374932
rect 364944 374892 364950 374904
rect 378134 374892 378140 374944
rect 378192 374932 378198 374944
rect 423950 374932 423956 374944
rect 378192 374904 423956 374932
rect 378192 374892 378198 374904
rect 423950 374892 423956 374904
rect 424008 374892 424014 374944
rect 208452 374836 215294 374864
rect 208452 374824 208458 374836
rect 217226 374824 217232 374876
rect 217284 374864 217290 374876
rect 262766 374864 262772 374876
rect 217284 374836 262772 374864
rect 217284 374824 217290 374836
rect 262766 374824 262772 374836
rect 262824 374824 262830 374876
rect 370314 374824 370320 374876
rect 370372 374864 370378 374876
rect 373994 374864 374000 374876
rect 370372 374836 374000 374864
rect 370372 374824 370378 374836
rect 373994 374824 374000 374836
rect 374052 374864 374058 374876
rect 422662 374864 422668 374876
rect 374052 374836 422668 374864
rect 374052 374824 374058 374836
rect 422662 374824 422668 374836
rect 422720 374824 422726 374876
rect 211062 374796 211068 374808
rect 205606 374768 211068 374796
rect 211062 374756 211068 374768
rect 211120 374796 211126 374808
rect 219434 374796 219440 374808
rect 211120 374768 219440 374796
rect 211120 374756 211126 374768
rect 219434 374756 219440 374768
rect 219492 374796 219498 374808
rect 267550 374796 267556 374808
rect 219492 374768 267556 374796
rect 219492 374756 219498 374768
rect 267550 374756 267556 374768
rect 267608 374756 267614 374808
rect 360654 374756 360660 374808
rect 360712 374796 360718 374808
rect 372338 374796 372344 374808
rect 360712 374768 372344 374796
rect 360712 374756 360718 374768
rect 372338 374756 372344 374768
rect 372396 374796 372402 374808
rect 429654 374796 429660 374808
rect 372396 374768 429660 374796
rect 372396 374756 372402 374768
rect 429654 374756 429660 374768
rect 429712 374756 429718 374808
rect 206738 374728 206744 374740
rect 195946 374700 206744 374728
rect 206738 374688 206744 374700
rect 206796 374728 206802 374740
rect 219342 374728 219348 374740
rect 206796 374700 219348 374728
rect 206796 374688 206802 374700
rect 219342 374688 219348 374700
rect 219400 374728 219406 374740
rect 266354 374728 266360 374740
rect 219400 374700 266360 374728
rect 219400 374688 219406 374700
rect 266354 374688 266360 374700
rect 266412 374688 266418 374740
rect 428550 374728 428556 374740
rect 369688 374700 428556 374728
rect 369688 374672 369716 374700
rect 428550 374688 428556 374700
rect 428608 374688 428614 374740
rect 183462 374620 183468 374672
rect 183520 374660 183526 374672
rect 197630 374660 197636 374672
rect 183520 374632 197636 374660
rect 183520 374620 183526 374632
rect 197630 374620 197636 374632
rect 197688 374660 197694 374672
rect 342254 374660 342260 374672
rect 197688 374632 342260 374660
rect 197688 374620 197694 374632
rect 342254 374620 342260 374632
rect 342312 374620 342318 374672
rect 357250 374620 357256 374672
rect 357308 374660 357314 374672
rect 369670 374660 369676 374672
rect 357308 374632 369676 374660
rect 357308 374620 357314 374632
rect 369670 374620 369676 374632
rect 369728 374620 369734 374672
rect 371694 374620 371700 374672
rect 371752 374660 371758 374672
rect 378134 374660 378140 374672
rect 371752 374632 378140 374660
rect 371752 374620 371758 374632
rect 378134 374620 378140 374632
rect 378192 374620 378198 374672
rect 379422 374620 379428 374672
rect 379480 374660 379486 374672
rect 439038 374660 439044 374672
rect 379480 374632 439044 374660
rect 379480 374620 379486 374632
rect 439038 374620 439044 374632
rect 439096 374620 439102 374672
rect 519354 371940 519360 371952
rect 509206 371912 519360 371940
rect 199378 371832 199384 371884
rect 199436 371872 199442 371884
rect 199562 371872 199568 371884
rect 199436 371844 199568 371872
rect 199436 371832 199442 371844
rect 199562 371832 199568 371844
rect 199620 371872 199626 371884
rect 359182 371872 359188 371884
rect 199620 371844 359188 371872
rect 199620 371832 199626 371844
rect 359182 371832 359188 371844
rect 359240 371872 359246 371884
rect 359458 371872 359464 371884
rect 359240 371844 359464 371872
rect 359240 371832 359246 371844
rect 359458 371832 359464 371844
rect 359516 371832 359522 371884
rect 359734 371832 359740 371884
rect 359792 371872 359798 371884
rect 509206 371872 509234 371912
rect 519354 371900 519360 371912
rect 519412 371940 519418 371952
rect 519538 371940 519544 371952
rect 519412 371912 519544 371940
rect 519412 371900 519418 371912
rect 519538 371900 519544 371912
rect 519596 371900 519602 371952
rect 359792 371844 509234 371872
rect 359792 371832 359798 371844
rect 199470 370472 199476 370524
rect 199528 370512 199534 370524
rect 359090 370512 359096 370524
rect 199528 370484 359096 370512
rect 199528 370472 199534 370484
rect 359090 370472 359096 370484
rect 359148 370472 359154 370524
rect 359090 369860 359096 369912
rect 359148 369900 359154 369912
rect 359642 369900 359648 369912
rect 359148 369872 359648 369900
rect 359148 369860 359154 369872
rect 359642 369860 359648 369872
rect 359700 369860 359706 369912
rect 207014 369792 207020 369844
rect 207072 369832 207078 369844
rect 207198 369832 207204 369844
rect 207072 369804 207204 369832
rect 207072 369792 207078 369804
rect 207198 369792 207204 369804
rect 207256 369832 207262 369844
rect 358998 369832 359004 369844
rect 207256 369804 359004 369832
rect 207256 369792 207262 369804
rect 358998 369792 359004 369804
rect 359056 369792 359062 369844
rect 199562 369112 199568 369164
rect 199620 369152 199626 369164
rect 207014 369152 207020 369164
rect 199620 369124 207020 369152
rect 199620 369112 199626 369124
rect 207014 369112 207020 369124
rect 207072 369112 207078 369164
rect 359458 369112 359464 369164
rect 359516 369152 359522 369164
rect 519170 369152 519176 369164
rect 359516 369124 519176 369152
rect 359516 369112 359522 369124
rect 519170 369112 519176 369124
rect 519228 369112 519234 369164
rect 358998 366324 359004 366376
rect 359056 366364 359062 366376
rect 359550 366364 359556 366376
rect 359056 366336 359556 366364
rect 359056 366324 359062 366336
rect 359550 366324 359556 366336
rect 359608 366364 359614 366376
rect 519078 366364 519084 366376
rect 359608 366336 519084 366364
rect 359608 366324 359614 366336
rect 519078 366324 519084 366336
rect 519136 366364 519142 366376
rect 519354 366364 519360 366376
rect 519136 366336 519360 366364
rect 519136 366324 519142 366336
rect 519354 366324 519360 366336
rect 519412 366324 519418 366376
rect 359642 363672 359648 363724
rect 359700 363712 359706 363724
rect 518894 363712 518900 363724
rect 359700 363684 518900 363712
rect 359700 363672 359706 363684
rect 518894 363672 518900 363684
rect 518952 363672 518958 363724
rect 199746 363604 199752 363656
rect 199804 363644 199810 363656
rect 358998 363644 359004 363656
rect 199804 363616 359004 363644
rect 199804 363604 199810 363616
rect 358998 363604 359004 363616
rect 359056 363604 359062 363656
rect 358998 362924 359004 362976
rect 359056 362964 359062 362976
rect 359734 362964 359740 362976
rect 359056 362936 359740 362964
rect 359056 362924 359062 362936
rect 359734 362924 359740 362936
rect 359792 362924 359798 362976
rect 199654 362176 199660 362228
rect 199712 362216 199718 362228
rect 359182 362216 359188 362228
rect 199712 362188 359188 362216
rect 199712 362176 199718 362188
rect 359182 362176 359188 362188
rect 359240 362216 359246 362228
rect 519078 362216 519084 362228
rect 359240 362188 519084 362216
rect 359240 362176 359246 362188
rect 519078 362176 519084 362188
rect 519136 362216 519142 362228
rect 519262 362216 519268 362228
rect 519136 362188 519268 362216
rect 519136 362176 519142 362188
rect 519262 362176 519268 362188
rect 519320 362176 519326 362228
rect 201402 360204 201408 360256
rect 201460 360244 201466 360256
rect 206278 360244 206284 360256
rect 201460 360216 206284 360244
rect 201460 360204 201466 360216
rect 206278 360204 206284 360216
rect 206336 360204 206342 360256
rect 180150 360136 180156 360188
rect 180208 360176 180214 360188
rect 195882 360176 195888 360188
rect 180208 360148 195888 360176
rect 180208 360136 180214 360148
rect 195882 360136 195888 360148
rect 195940 360136 195946 360188
rect 195882 359660 195888 359712
rect 195940 359700 195946 359712
rect 197538 359700 197544 359712
rect 195940 359672 197544 359700
rect 195940 359660 195946 359672
rect 197538 359660 197544 359672
rect 197596 359660 197602 359712
rect 340046 359592 340052 359644
rect 340104 359632 340110 359644
rect 357526 359632 357532 359644
rect 340104 359604 357532 359632
rect 340104 359592 340110 359604
rect 357526 359592 357532 359604
rect 357584 359592 357590 359644
rect 500402 359592 500408 359644
rect 500460 359632 500466 359644
rect 517974 359632 517980 359644
rect 500460 359604 517980 359632
rect 500460 359592 500466 359604
rect 517974 359592 517980 359604
rect 518032 359592 518038 359644
rect 197354 359524 197360 359576
rect 197412 359564 197418 359576
rect 204622 359564 204628 359576
rect 197412 359536 204628 359564
rect 197412 359524 197418 359536
rect 204622 359524 204628 359536
rect 204680 359524 204686 359576
rect 338482 359524 338488 359576
rect 338540 359564 338546 359576
rect 356974 359564 356980 359576
rect 338540 359536 356980 359564
rect 338540 359524 338546 359536
rect 356974 359524 356980 359536
rect 357032 359524 357038 359576
rect 498930 359524 498936 359576
rect 498988 359564 498994 359576
rect 517790 359564 517796 359576
rect 498988 359536 517796 359564
rect 498988 359524 498994 359536
rect 517790 359524 517796 359536
rect 517848 359524 517854 359576
rect 190914 359456 190920 359508
rect 190972 359496 190978 359508
rect 200758 359496 200764 359508
rect 190972 359468 200764 359496
rect 190972 359456 190978 359468
rect 200758 359456 200764 359468
rect 200816 359496 200822 359508
rect 201402 359496 201408 359508
rect 200816 359468 201408 359496
rect 200816 359456 200822 359468
rect 201402 359456 201408 359468
rect 201460 359456 201466 359508
rect 351730 359456 351736 359508
rect 351788 359496 351794 359508
rect 358078 359496 358084 359508
rect 351788 359468 358084 359496
rect 351788 359456 351794 359468
rect 358078 359456 358084 359468
rect 358136 359456 358142 359508
rect 178586 358776 178592 358828
rect 178644 358816 178650 358828
rect 197354 358816 197360 358828
rect 178644 358788 197360 358816
rect 178644 358776 178650 358788
rect 197354 358776 197360 358788
rect 197412 358776 197418 358828
rect 342254 358776 342260 358828
rect 342312 358816 342318 358828
rect 343542 358816 343548 358828
rect 342312 358788 343548 358816
rect 342312 358776 342318 358788
rect 343542 358776 343548 358788
rect 343600 358816 343606 358828
rect 358814 358816 358820 358828
rect 343600 358788 358820 358816
rect 343600 358776 343606 358788
rect 358814 358776 358820 358788
rect 358872 358776 358878 358828
rect 510890 358776 510896 358828
rect 510948 358816 510954 358828
rect 517514 358816 517520 358828
rect 510948 358788 517520 358816
rect 510948 358776 510954 358788
rect 517514 358776 517520 358788
rect 517572 358776 517578 358828
rect 219250 358708 219256 358760
rect 219308 358748 219314 358760
rect 220814 358748 220820 358760
rect 219308 358720 220820 358748
rect 219308 358708 219314 358720
rect 220814 358708 220820 358720
rect 220872 358708 220878 358760
rect 57146 358640 57152 358692
rect 57204 358680 57210 358692
rect 59446 358680 59452 358692
rect 57204 358652 59452 358680
rect 57204 358640 57210 358652
rect 59446 358640 59452 358652
rect 59504 358640 59510 358692
rect 218606 358640 218612 358692
rect 218664 358680 218670 358692
rect 220998 358680 221004 358692
rect 218664 358652 221004 358680
rect 218664 358640 218670 358652
rect 220998 358640 221004 358652
rect 221056 358640 221062 358692
rect 377030 358572 377036 358624
rect 377088 358612 377094 358624
rect 381170 358612 381176 358624
rect 377088 358584 381176 358612
rect 377088 358572 377094 358584
rect 381170 358572 381176 358584
rect 381228 358572 381234 358624
rect 217134 358232 217140 358284
rect 217192 358272 217198 358284
rect 219434 358272 219440 358284
rect 217192 358244 219440 358272
rect 217192 358232 217198 358244
rect 219434 358232 219440 358244
rect 219492 358232 219498 358284
rect 379238 358096 379244 358148
rect 379296 358136 379302 358148
rect 380986 358136 380992 358148
rect 379296 358108 380992 358136
rect 379296 358096 379302 358108
rect 380986 358096 380992 358108
rect 381044 358096 381050 358148
rect 54478 358028 54484 358080
rect 54536 358068 54542 358080
rect 59354 358068 59360 358080
rect 54536 358040 59360 358068
rect 54536 358028 54542 358040
rect 59354 358028 59360 358040
rect 59412 358028 59418 358080
rect 182818 358028 182824 358080
rect 182876 358068 182882 358080
rect 201586 358068 201592 358080
rect 182876 358040 201592 358068
rect 182876 358028 182882 358040
rect 201586 358028 201592 358040
rect 201644 358068 201650 358080
rect 342254 358068 342260 358080
rect 201644 358040 342260 358068
rect 201644 358028 201650 358040
rect 342254 358028 342260 358040
rect 342312 358028 342318 358080
rect 373810 358028 373816 358080
rect 373868 358068 373874 358080
rect 381078 358068 381084 358080
rect 373868 358040 381084 358068
rect 373868 358028 373874 358040
rect 381078 358028 381084 358040
rect 381136 358028 381142 358080
rect 379422 357960 379428 358012
rect 379480 358000 379486 358012
rect 381262 358000 381268 358012
rect 379480 357972 381268 358000
rect 379480 357960 379486 357972
rect 381262 357960 381268 357972
rect 381320 357960 381326 358012
rect 219158 357824 219164 357876
rect 219216 357864 219222 357876
rect 220906 357864 220912 357876
rect 219216 357836 220912 357864
rect 219216 357824 219222 357836
rect 220906 357824 220912 357836
rect 220964 357824 220970 357876
rect 378686 357824 378692 357876
rect 378744 357864 378750 357876
rect 380894 357864 380900 357876
rect 378744 357836 380900 357864
rect 378744 357824 378750 357836
rect 380894 357824 380900 357836
rect 380952 357824 380958 357876
rect 58526 357348 58532 357400
rect 58584 357388 58590 357400
rect 60734 357388 60740 357400
rect 58584 357360 60740 357388
rect 58584 357348 58590 357360
rect 60734 357348 60740 357360
rect 60792 357348 60798 357400
rect 46382 303560 46388 303612
rect 46440 303600 46446 303612
rect 57330 303600 57336 303612
rect 46440 303572 57336 303600
rect 46440 303560 46446 303572
rect 57330 303560 57336 303572
rect 57388 303600 57394 303612
rect 57514 303600 57520 303612
rect 57388 303572 57520 303600
rect 57388 303560 57394 303572
rect 57514 303560 57520 303572
rect 57572 303560 57578 303612
rect 46474 300772 46480 300824
rect 46532 300812 46538 300824
rect 56778 300812 56784 300824
rect 46532 300784 56784 300812
rect 46532 300772 46538 300784
rect 56778 300772 56784 300784
rect 56836 300772 56842 300824
rect 56962 300772 56968 300824
rect 57020 300812 57026 300824
rect 58434 300812 58440 300824
rect 57020 300784 58440 300812
rect 57020 300772 57026 300784
rect 58434 300772 58440 300784
rect 58492 300772 58498 300824
rect 56796 300744 56824 300772
rect 57054 300744 57060 300756
rect 56796 300716 57060 300744
rect 57054 300704 57060 300716
rect 57112 300704 57118 300756
rect 520182 288396 520188 288448
rect 520240 288436 520246 288448
rect 580258 288436 580264 288448
rect 520240 288408 580264 288436
rect 520240 288396 520246 288408
rect 580258 288396 580264 288408
rect 580316 288396 580322 288448
rect 518986 287036 518992 287088
rect 519044 287076 519050 287088
rect 580350 287076 580356 287088
rect 519044 287048 580356 287076
rect 519044 287036 519050 287048
rect 580350 287036 580356 287048
rect 580408 287036 580414 287088
rect 200942 284248 200948 284300
rect 201000 284288 201006 284300
rect 216674 284288 216680 284300
rect 201000 284260 216680 284288
rect 201000 284248 201006 284260
rect 216674 284248 216680 284260
rect 216732 284248 216738 284300
rect 361298 284248 361304 284300
rect 361356 284288 361362 284300
rect 376846 284288 376852 284300
rect 361356 284260 376852 284288
rect 361356 284248 361362 284260
rect 376846 284248 376852 284260
rect 376904 284248 376910 284300
rect 203886 282820 203892 282872
rect 203944 282860 203950 282872
rect 216766 282860 216772 282872
rect 203944 282832 216772 282860
rect 203944 282820 203950 282832
rect 216766 282820 216772 282832
rect 216824 282820 216830 282872
rect 366818 282820 366824 282872
rect 366876 282860 366882 282872
rect 377582 282860 377588 282872
rect 366876 282832 377588 282860
rect 366876 282820 366882 282832
rect 377582 282820 377588 282832
rect 377640 282820 377646 282872
rect 55858 282616 55864 282668
rect 55916 282656 55922 282668
rect 58618 282656 58624 282668
rect 55916 282628 58624 282656
rect 55916 282616 55922 282628
rect 58618 282616 58624 282628
rect 58676 282616 58682 282668
rect 51534 282140 51540 282192
rect 51592 282180 51598 282192
rect 58342 282180 58348 282192
rect 51592 282152 58348 282180
rect 51592 282140 51598 282152
rect 58342 282140 58348 282152
rect 58400 282140 58406 282192
rect 200758 282140 200764 282192
rect 200816 282180 200822 282192
rect 201402 282180 201408 282192
rect 200816 282152 201408 282180
rect 200816 282140 200822 282152
rect 201402 282140 201408 282152
rect 201460 282180 201466 282192
rect 216674 282180 216680 282192
rect 201460 282152 216680 282180
rect 201460 282140 201466 282152
rect 216674 282140 216680 282152
rect 216732 282140 216738 282192
rect 358078 282140 358084 282192
rect 358136 282180 358142 282192
rect 376938 282180 376944 282192
rect 358136 282152 376944 282180
rect 358136 282140 358142 282152
rect 376938 282140 376944 282152
rect 376996 282140 377002 282192
rect 370406 273912 370412 273964
rect 370464 273952 370470 273964
rect 370866 273952 370872 273964
rect 370464 273924 370872 273952
rect 370464 273912 370470 273924
rect 370866 273912 370872 273924
rect 370924 273912 370930 273964
rect 43622 273572 43628 273624
rect 43680 273612 43686 273624
rect 133414 273612 133420 273624
rect 43680 273584 133420 273612
rect 43680 273572 43686 273584
rect 133414 273572 133420 273584
rect 133472 273572 133478 273624
rect 371050 273572 371056 273624
rect 371108 273612 371114 273624
rect 378134 273612 378140 273624
rect 371108 273584 378140 273612
rect 371108 273572 371114 273584
rect 378134 273572 378140 273584
rect 378192 273572 378198 273624
rect 378686 273572 378692 273624
rect 378744 273612 378750 273624
rect 379698 273612 379704 273624
rect 378744 273584 379704 273612
rect 378744 273572 378750 273584
rect 379698 273572 379704 273584
rect 379756 273612 379762 273624
rect 426434 273612 426440 273624
rect 379756 273584 426440 273612
rect 379756 273572 379762 273584
rect 426434 273572 426440 273584
rect 426492 273572 426498 273624
rect 44818 273504 44824 273556
rect 44876 273544 44882 273556
rect 135898 273544 135904 273556
rect 44876 273516 135904 273544
rect 44876 273504 44882 273516
rect 135898 273504 135904 273516
rect 135956 273504 135962 273556
rect 369486 273504 369492 273556
rect 369544 273544 369550 273556
rect 421098 273544 421104 273556
rect 369544 273516 421104 273544
rect 369544 273504 369550 273516
rect 421098 273504 421104 273516
rect 421156 273504 421162 273556
rect 44910 273436 44916 273488
rect 44968 273476 44974 273488
rect 138474 273476 138480 273488
rect 44968 273448 138480 273476
rect 44968 273436 44974 273448
rect 138474 273436 138480 273448
rect 138532 273436 138538 273488
rect 370958 273436 370964 273488
rect 371016 273476 371022 273488
rect 373074 273476 373080 273488
rect 371016 273448 373080 273476
rect 371016 273436 371022 273448
rect 373074 273436 373080 273448
rect 373132 273476 373138 273488
rect 431126 273476 431132 273488
rect 373132 273448 431132 273476
rect 373132 273436 373138 273448
rect 431126 273436 431132 273448
rect 431184 273436 431190 273488
rect 45002 273368 45008 273420
rect 45060 273408 45066 273420
rect 140866 273408 140872 273420
rect 45060 273380 140872 273408
rect 45060 273368 45066 273380
rect 140866 273368 140872 273380
rect 140924 273368 140930 273420
rect 219342 273368 219348 273420
rect 219400 273408 219406 273420
rect 219894 273408 219900 273420
rect 219400 273380 219900 273408
rect 219400 273368 219406 273380
rect 219894 273368 219900 273380
rect 219952 273408 219958 273420
rect 266354 273408 266360 273420
rect 219952 273380 266360 273408
rect 219952 273368 219958 273380
rect 266354 273368 266360 273380
rect 266412 273368 266418 273420
rect 373810 273368 373816 273420
rect 373868 273408 373874 273420
rect 433334 273408 433340 273420
rect 373868 273380 433340 273408
rect 373868 273368 373874 273380
rect 433334 273368 433340 273380
rect 433392 273368 433398 273420
rect 45094 273300 45100 273352
rect 45152 273340 45158 273352
rect 143534 273340 143540 273352
rect 45152 273312 143540 273340
rect 45152 273300 45158 273312
rect 143534 273300 143540 273312
rect 143592 273300 143598 273352
rect 214190 273300 214196 273352
rect 214248 273340 214254 273352
rect 214926 273340 214932 273352
rect 214248 273312 214932 273340
rect 214248 273300 214254 273312
rect 214926 273300 214932 273312
rect 214984 273340 214990 273352
rect 273254 273340 273260 273352
rect 214984 273312 273260 273340
rect 214984 273300 214990 273312
rect 273254 273300 273260 273312
rect 273312 273300 273318 273352
rect 356882 273300 356888 273352
rect 356940 273340 356946 273352
rect 430942 273340 430948 273352
rect 356940 273312 430948 273340
rect 356940 273300 356946 273312
rect 430942 273300 430948 273312
rect 431000 273300 431006 273352
rect 45186 273232 45192 273284
rect 45244 273272 45250 273284
rect 145926 273272 145932 273284
rect 45244 273244 145932 273272
rect 45244 273232 45250 273244
rect 145926 273232 145932 273244
rect 145984 273232 145990 273284
rect 210970 273232 210976 273284
rect 211028 273272 211034 273284
rect 283466 273272 283472 273284
rect 211028 273244 283472 273272
rect 211028 273232 211034 273244
rect 283466 273232 283472 273244
rect 283524 273232 283530 273284
rect 369762 273232 369768 273284
rect 369820 273272 369826 273284
rect 369820 273244 373580 273272
rect 369820 273232 369826 273244
rect 373552 273204 373580 273244
rect 373626 273232 373632 273284
rect 373684 273272 373690 273284
rect 453390 273272 453396 273284
rect 373684 273244 453396 273272
rect 373684 273232 373690 273244
rect 453390 273232 453396 273244
rect 453448 273232 453454 273284
rect 373994 273204 374000 273216
rect 373552 273176 374000 273204
rect 373994 273164 374000 273176
rect 374052 273204 374058 273216
rect 422846 273204 422852 273216
rect 374052 273176 422852 273204
rect 374052 273164 374058 273176
rect 422846 273164 422852 273176
rect 422904 273164 422910 273216
rect 361206 273096 361212 273148
rect 361264 273136 361270 273148
rect 425974 273136 425980 273148
rect 361264 273108 425980 273136
rect 361264 273096 361270 273108
rect 425974 273096 425980 273108
rect 426032 273096 426038 273148
rect 46658 273028 46664 273080
rect 46716 273068 46722 273080
rect 51534 273068 51540 273080
rect 46716 273040 51540 273068
rect 46716 273028 46722 273040
rect 51534 273028 51540 273040
rect 51592 273068 51598 273080
rect 95878 273068 95884 273080
rect 51592 273040 95884 273068
rect 51592 273028 51598 273040
rect 95878 273028 95884 273040
rect 95936 273028 95942 273080
rect 209314 273028 209320 273080
rect 209372 273068 209378 273080
rect 288158 273068 288164 273080
rect 209372 273040 288164 273068
rect 209372 273028 209378 273040
rect 288158 273028 288164 273040
rect 288216 273028 288222 273080
rect 358446 273028 358452 273080
rect 358504 273068 358510 273080
rect 423398 273068 423404 273080
rect 358504 273040 423404 273068
rect 358504 273028 358510 273040
rect 423398 273028 423404 273040
rect 423456 273028 423462 273080
rect 49142 272960 49148 273012
rect 49200 273000 49206 273012
rect 54294 273000 54300 273012
rect 49200 272972 54300 273000
rect 49200 272960 49206 272972
rect 54294 272960 54300 272972
rect 54352 273000 54358 273012
rect 82998 273000 83004 273012
rect 54352 272972 83004 273000
rect 54352 272960 54358 272972
rect 82998 272960 83004 272972
rect 83056 272960 83062 273012
rect 207934 272960 207940 273012
rect 207992 273000 207998 273012
rect 285950 273000 285956 273012
rect 207992 272972 285956 273000
rect 207992 272960 207998 272972
rect 285950 272960 285956 272972
rect 286008 272960 286014 273012
rect 370774 272960 370780 273012
rect 370832 273000 370838 273012
rect 468478 273000 468484 273012
rect 370832 272972 468484 273000
rect 370832 272960 370838 272972
rect 468478 272960 468484 272972
rect 468536 272960 468542 273012
rect 58434 272892 58440 272944
rect 58492 272932 58498 272944
rect 61010 272932 61016 272944
rect 58492 272904 61016 272932
rect 58492 272892 58498 272904
rect 61010 272892 61016 272904
rect 61068 272932 61074 272944
rect 61470 272932 61476 272944
rect 61068 272904 61476 272932
rect 61068 272892 61074 272904
rect 61470 272892 61476 272904
rect 61528 272892 61534 272944
rect 212258 272892 212264 272944
rect 212316 272932 212322 272944
rect 295886 272932 295892 272944
rect 212316 272904 295892 272932
rect 212316 272892 212322 272904
rect 295886 272892 295892 272904
rect 295944 272892 295950 272944
rect 372246 272892 372252 272944
rect 372304 272932 372310 272944
rect 470870 272932 470876 272944
rect 372304 272904 470876 272932
rect 372304 272892 372310 272904
rect 470870 272892 470876 272904
rect 470928 272892 470934 272944
rect 202414 272824 202420 272876
rect 202472 272864 202478 272876
rect 290918 272864 290924 272876
rect 202472 272836 290924 272864
rect 202472 272824 202478 272836
rect 290918 272824 290924 272836
rect 290976 272824 290982 272876
rect 375006 272824 375012 272876
rect 375064 272864 375070 272876
rect 473446 272864 473452 272876
rect 375064 272836 473452 272864
rect 375064 272824 375070 272836
rect 473446 272824 473452 272836
rect 473504 272824 473510 272876
rect 50338 272756 50344 272808
rect 50396 272796 50402 272808
rect 53834 272796 53840 272808
rect 50396 272768 53840 272796
rect 50396 272756 50402 272768
rect 53834 272756 53840 272768
rect 53892 272756 53898 272808
rect 210786 272756 210792 272808
rect 210844 272796 210850 272808
rect 303430 272796 303436 272808
rect 210844 272768 303436 272796
rect 210844 272756 210850 272768
rect 303430 272756 303436 272768
rect 303488 272756 303494 272808
rect 368106 272756 368112 272808
rect 368164 272796 368170 272808
rect 475838 272796 475844 272808
rect 368164 272768 475844 272796
rect 368164 272756 368170 272768
rect 475838 272756 475844 272768
rect 475896 272756 475902 272808
rect 50430 272688 50436 272740
rect 50488 272728 50494 272740
rect 90726 272728 90732 272740
rect 50488 272700 90732 272728
rect 50488 272688 50494 272700
rect 90726 272688 90732 272700
rect 90784 272688 90790 272740
rect 205082 272688 205088 272740
rect 205140 272728 205146 272740
rect 298462 272728 298468 272740
rect 205140 272700 298468 272728
rect 205140 272688 205146 272700
rect 298462 272688 298468 272700
rect 298520 272688 298526 272740
rect 365438 272688 365444 272740
rect 365496 272728 365502 272740
rect 478414 272728 478420 272740
rect 365496 272700 478420 272728
rect 365496 272688 365502 272700
rect 478414 272688 478420 272700
rect 478472 272688 478478 272740
rect 48038 272620 48044 272672
rect 48096 272660 48102 272672
rect 93670 272660 93676 272672
rect 48096 272632 93676 272660
rect 48096 272620 48102 272632
rect 93670 272620 93676 272632
rect 93728 272620 93734 272672
rect 200850 272620 200856 272672
rect 200908 272660 200914 272672
rect 300854 272660 300860 272672
rect 200908 272632 300860 272660
rect 200908 272620 200914 272632
rect 300854 272620 300860 272632
rect 300912 272620 300918 272672
rect 362586 272620 362592 272672
rect 362644 272660 362650 272672
rect 480806 272660 480812 272672
rect 362644 272632 480812 272660
rect 362644 272620 362650 272632
rect 480806 272620 480812 272632
rect 480864 272620 480870 272672
rect 49234 272552 49240 272604
rect 49292 272592 49298 272604
rect 96062 272592 96068 272604
rect 49292 272564 96068 272592
rect 49292 272552 49298 272564
rect 96062 272552 96068 272564
rect 96120 272552 96126 272604
rect 203794 272552 203800 272604
rect 203852 272592 203858 272604
rect 305822 272592 305828 272604
rect 203852 272564 305828 272592
rect 203852 272552 203858 272564
rect 305822 272552 305828 272564
rect 305880 272552 305886 272604
rect 364058 272552 364064 272604
rect 364116 272592 364122 272604
rect 483198 272592 483204 272604
rect 364116 272564 483204 272592
rect 364116 272552 364122 272564
rect 483198 272552 483204 272564
rect 483256 272552 483262 272604
rect 51902 272484 51908 272536
rect 51960 272524 51966 272536
rect 98454 272524 98460 272536
rect 51960 272496 98460 272524
rect 51960 272484 51966 272496
rect 98454 272484 98460 272496
rect 98512 272484 98518 272536
rect 197170 272524 197176 272536
rect 103486 272496 197176 272524
rect 47854 272416 47860 272468
rect 47912 272456 47918 272468
rect 77110 272456 77116 272468
rect 47912 272428 77116 272456
rect 47912 272416 47918 272428
rect 77110 272416 77116 272428
rect 77168 272416 77174 272468
rect 98086 272416 98092 272468
rect 98144 272456 98150 272468
rect 103486 272456 103514 272496
rect 197170 272484 197176 272496
rect 197228 272484 197234 272536
rect 202506 272484 202512 272536
rect 202564 272524 202570 272536
rect 320910 272524 320916 272536
rect 202564 272496 320916 272524
rect 202564 272484 202570 272496
rect 320910 272484 320916 272496
rect 320968 272484 320974 272536
rect 366726 272484 366732 272536
rect 366784 272524 366790 272536
rect 485958 272524 485964 272536
rect 366784 272496 485964 272524
rect 366784 272484 366790 272496
rect 485958 272484 485964 272496
rect 486016 272484 486022 272536
rect 98144 272428 103514 272456
rect 98144 272416 98150 272428
rect 378134 272416 378140 272468
rect 378192 272456 378198 272468
rect 423766 272456 423772 272468
rect 378192 272428 423772 272456
rect 378192 272416 378198 272428
rect 423766 272416 423772 272428
rect 423824 272416 423830 272468
rect 46566 272348 46572 272400
rect 46624 272388 46630 272400
rect 76006 272388 76012 272400
rect 46624 272360 76012 272388
rect 46624 272348 46630 272360
rect 76006 272348 76012 272360
rect 76064 272348 76070 272400
rect 59630 272280 59636 272332
rect 59688 272320 59694 272332
rect 60826 272320 60832 272332
rect 59688 272292 60832 272320
rect 59688 272280 59694 272292
rect 60826 272280 60832 272292
rect 60884 272280 60890 272332
rect 62206 272280 62212 272332
rect 62264 272320 62270 272332
rect 94406 272320 94412 272332
rect 62264 272292 94412 272320
rect 62264 272280 62270 272292
rect 94406 272280 94412 272292
rect 94464 272280 94470 272332
rect 54110 272212 54116 272264
rect 54168 272252 54174 272264
rect 54754 272252 54760 272264
rect 54168 272224 54760 272252
rect 54168 272212 54174 272224
rect 54754 272212 54760 272224
rect 54812 272252 54818 272264
rect 87598 272252 87604 272264
rect 54812 272224 87604 272252
rect 54812 272212 54818 272224
rect 87598 272212 87604 272224
rect 87656 272212 87662 272264
rect 58342 272144 58348 272196
rect 58400 272184 58406 272196
rect 59722 272184 59728 272196
rect 58400 272156 59728 272184
rect 58400 272144 58406 272156
rect 59722 272144 59728 272156
rect 59780 272184 59786 272196
rect 99374 272184 99380 272196
rect 59780 272156 99380 272184
rect 59780 272144 59786 272156
rect 99374 272144 99380 272156
rect 99432 272144 99438 272196
rect 58618 272076 58624 272128
rect 58676 272116 58682 272128
rect 100754 272116 100760 272128
rect 58676 272088 100760 272116
rect 58676 272076 58682 272088
rect 100754 272076 100760 272088
rect 100812 272076 100818 272128
rect 356882 272076 356888 272128
rect 356940 272116 356946 272128
rect 358814 272116 358820 272128
rect 356940 272088 358820 272116
rect 356940 272076 356946 272088
rect 358814 272076 358820 272088
rect 358872 272076 358878 272128
rect 47946 272008 47952 272060
rect 48004 272048 48010 272060
rect 52822 272048 52828 272060
rect 48004 272020 52828 272048
rect 48004 272008 48010 272020
rect 52822 272008 52828 272020
rect 52880 272048 52886 272060
rect 96614 272048 96620 272060
rect 52880 272020 96620 272048
rect 52880 272008 52886 272020
rect 96614 272008 96620 272020
rect 96672 272008 96678 272060
rect 85758 271940 85764 271992
rect 85816 271980 85822 271992
rect 106550 271980 106556 271992
rect 85816 271952 106556 271980
rect 85816 271940 85822 271952
rect 106550 271940 106556 271952
rect 106608 271940 106614 271992
rect 427078 271940 427084 271992
rect 427136 271980 427142 271992
rect 436094 271980 436100 271992
rect 427136 271952 436100 271980
rect 427136 271940 427142 271952
rect 436094 271940 436100 271952
rect 436152 271940 436158 271992
rect 60826 271872 60832 271924
rect 60884 271912 60890 271924
rect 106274 271912 106280 271924
rect 60884 271884 106280 271912
rect 60884 271872 60890 271884
rect 106274 271872 106280 271884
rect 106332 271872 106338 271924
rect 112346 271872 112352 271924
rect 112404 271912 112410 271924
rect 196618 271912 196624 271924
rect 112404 271884 196624 271912
rect 112404 271872 112410 271884
rect 196618 271872 196624 271884
rect 196676 271872 196682 271924
rect 396718 271872 396724 271924
rect 396776 271912 396782 271924
rect 415854 271912 415860 271924
rect 396776 271884 415860 271912
rect 396776 271872 396782 271884
rect 415854 271872 415860 271884
rect 415912 271872 415918 271924
rect 425698 271872 425704 271924
rect 425756 271912 425762 271924
rect 427814 271912 427820 271924
rect 425756 271884 427820 271912
rect 425756 271872 425762 271884
rect 427814 271872 427820 271884
rect 427872 271872 427878 271924
rect 42426 271804 42432 271856
rect 42484 271844 42490 271856
rect 123110 271844 123116 271856
rect 42484 271816 123116 271844
rect 42484 271804 42490 271816
rect 123110 271804 123116 271816
rect 123168 271804 123174 271856
rect 154482 271804 154488 271856
rect 154540 271844 154546 271856
rect 201770 271844 201776 271856
rect 154540 271816 201776 271844
rect 154540 271804 154546 271816
rect 201770 271804 201776 271816
rect 201828 271804 201834 271856
rect 213178 271804 213184 271856
rect 213236 271844 213242 271856
rect 313274 271844 313280 271856
rect 213236 271816 313280 271844
rect 213236 271804 213242 271816
rect 313274 271804 313280 271816
rect 313332 271804 313338 271856
rect 358354 271804 358360 271856
rect 358412 271844 358418 271856
rect 455782 271844 455788 271856
rect 358412 271816 455788 271844
rect 358412 271804 358418 271816
rect 455782 271804 455788 271816
rect 455840 271804 455846 271856
rect 517698 271804 517704 271856
rect 517756 271844 517762 271856
rect 517882 271844 517888 271856
rect 517756 271816 517888 271844
rect 517756 271804 517762 271816
rect 517882 271804 517888 271816
rect 517940 271804 517946 271856
rect 57146 271736 57152 271788
rect 57204 271776 57210 271788
rect 128354 271776 128360 271788
rect 57204 271748 128360 271776
rect 57204 271736 57210 271748
rect 128354 271736 128360 271748
rect 128412 271736 128418 271788
rect 151354 271736 151360 271788
rect 151412 271776 151418 271788
rect 198918 271776 198924 271788
rect 151412 271748 198924 271776
rect 151412 271736 151418 271748
rect 198918 271736 198924 271748
rect 198976 271736 198982 271788
rect 212166 271736 212172 271788
rect 212224 271776 212230 271788
rect 307754 271776 307760 271788
rect 212224 271748 307760 271776
rect 212224 271736 212230 271748
rect 307754 271736 307760 271748
rect 307812 271736 307818 271788
rect 368014 271736 368020 271788
rect 368072 271776 368078 271788
rect 458174 271776 458180 271788
rect 368072 271748 458180 271776
rect 368072 271736 368078 271748
rect 458174 271736 458180 271748
rect 458232 271736 458238 271788
rect 54478 271668 54484 271720
rect 54536 271708 54542 271720
rect 125594 271708 125600 271720
rect 54536 271680 125600 271708
rect 54536 271668 54542 271680
rect 125594 271668 125600 271680
rect 125652 271668 125658 271720
rect 157242 271668 157248 271720
rect 157300 271708 157306 271720
rect 203058 271708 203064 271720
rect 157300 271680 203064 271708
rect 157300 271668 157306 271680
rect 203058 271668 203064 271680
rect 203116 271668 203122 271720
rect 206462 271668 206468 271720
rect 206520 271708 206526 271720
rect 280246 271708 280252 271720
rect 206520 271680 280252 271708
rect 206520 271668 206526 271680
rect 280246 271668 280252 271680
rect 280304 271668 280310 271720
rect 365346 271668 365352 271720
rect 365404 271708 365410 271720
rect 447134 271708 447140 271720
rect 365404 271680 447140 271708
rect 365404 271668 365410 271680
rect 447134 271668 447140 271680
rect 447192 271668 447198 271720
rect 54570 271600 54576 271652
rect 54628 271640 54634 271652
rect 120074 271640 120080 271652
rect 54628 271612 120080 271640
rect 54628 271600 54634 271612
rect 120074 271600 120080 271612
rect 120132 271600 120138 271652
rect 158622 271600 158628 271652
rect 158680 271640 158686 271652
rect 198366 271640 198372 271652
rect 158680 271612 198372 271640
rect 158680 271600 158686 271612
rect 198366 271600 198372 271612
rect 198424 271600 198430 271652
rect 202322 271600 202328 271652
rect 202380 271640 202386 271652
rect 270494 271640 270500 271652
rect 202380 271612 270500 271640
rect 202380 271600 202386 271612
rect 270494 271600 270500 271612
rect 270552 271600 270558 271652
rect 370682 271600 370688 271652
rect 370740 271640 370746 271652
rect 449894 271640 449900 271652
rect 370740 271612 449900 271640
rect 370740 271600 370746 271612
rect 449894 271600 449900 271612
rect 449952 271600 449958 271652
rect 54662 271532 54668 271584
rect 54720 271572 54726 271584
rect 117314 271572 117320 271584
rect 54720 271544 117320 271572
rect 54720 271532 54726 271544
rect 117314 271532 117320 271544
rect 117372 271532 117378 271584
rect 161290 271532 161296 271584
rect 161348 271572 161354 271584
rect 204806 271572 204812 271584
rect 161348 271544 204812 271572
rect 161348 271532 161354 271544
rect 204806 271532 204812 271544
rect 204864 271532 204870 271584
rect 216122 271532 216128 271584
rect 216180 271572 216186 271584
rect 276014 271572 276020 271584
rect 216180 271544 276020 271572
rect 216180 271532 216186 271544
rect 276014 271532 276020 271544
rect 276072 271532 276078 271584
rect 364150 271532 364156 271584
rect 364208 271572 364214 271584
rect 442994 271572 443000 271584
rect 364208 271544 443000 271572
rect 364208 271532 364214 271544
rect 442994 271532 443000 271544
rect 443052 271532 443058 271584
rect 53190 271464 53196 271516
rect 53248 271504 53254 271516
rect 115934 271504 115940 271516
rect 53248 271476 115940 271504
rect 53248 271464 53254 271476
rect 115934 271464 115940 271476
rect 115992 271464 115998 271516
rect 164142 271464 164148 271516
rect 164200 271504 164206 271516
rect 197722 271504 197728 271516
rect 164200 271476 197728 271504
rect 164200 271464 164206 271476
rect 197722 271464 197728 271476
rect 197780 271464 197786 271516
rect 204990 271464 204996 271516
rect 205048 271504 205054 271516
rect 263594 271504 263600 271516
rect 205048 271476 263600 271504
rect 205048 271464 205054 271476
rect 263594 271464 263600 271476
rect 263652 271464 263658 271516
rect 362678 271464 362684 271516
rect 362736 271504 362742 271516
rect 437474 271504 437480 271516
rect 362736 271476 437480 271504
rect 362736 271464 362742 271476
rect 437474 271464 437480 271476
rect 437532 271464 437538 271516
rect 53098 271396 53104 271448
rect 53156 271436 53162 271448
rect 53156 271408 108344 271436
rect 53156 271396 53162 271408
rect 52914 271328 52920 271380
rect 52972 271368 52978 271380
rect 52972 271340 106872 271368
rect 52972 271328 52978 271340
rect 53006 271260 53012 271312
rect 53064 271300 53070 271312
rect 53064 271272 105952 271300
rect 53064 271260 53070 271272
rect 51626 271192 51632 271244
rect 51684 271232 51690 271244
rect 104894 271232 104900 271244
rect 51684 271204 104900 271232
rect 51684 271192 51690 271204
rect 104894 271192 104900 271204
rect 104952 271192 104958 271244
rect 51810 271124 51816 271176
rect 51868 271164 51874 271176
rect 103514 271164 103520 271176
rect 51868 271136 103520 271164
rect 51868 271124 51874 271136
rect 103514 271124 103520 271136
rect 103572 271124 103578 271176
rect 50246 271056 50252 271108
rect 50304 271096 50310 271108
rect 100754 271096 100760 271108
rect 50304 271068 100760 271096
rect 50304 271056 50310 271068
rect 100754 271056 100760 271068
rect 100812 271056 100818 271108
rect 105924 271096 105952 271272
rect 106844 271164 106872 271340
rect 108316 271232 108344 271408
rect 197354 271396 197360 271448
rect 197412 271436 197418 271448
rect 197630 271436 197636 271448
rect 197412 271408 197636 271436
rect 197412 271396 197418 271408
rect 197630 271396 197636 271408
rect 197688 271396 197694 271448
rect 219066 271396 219072 271448
rect 219124 271436 219130 271448
rect 277946 271436 277952 271448
rect 219124 271408 277952 271436
rect 219124 271396 219130 271408
rect 277946 271396 277952 271408
rect 278004 271396 278010 271448
rect 343542 271396 343548 271448
rect 343600 271436 343606 271448
rect 356882 271436 356888 271448
rect 343600 271408 356888 271436
rect 343600 271396 343606 271408
rect 356882 271396 356888 271408
rect 356940 271396 356946 271448
rect 372154 271396 372160 271448
rect 372212 271436 372218 271448
rect 445754 271436 445760 271448
rect 372212 271408 445760 271436
rect 372212 271396 372218 271408
rect 445754 271396 445760 271408
rect 445812 271396 445818 271448
rect 210878 271328 210884 271380
rect 210936 271368 210942 271380
rect 268010 271368 268016 271380
rect 210936 271340 268016 271368
rect 210936 271328 210942 271340
rect 268010 271328 268016 271340
rect 268068 271328 268074 271380
rect 361114 271328 361120 271380
rect 361172 271368 361178 271380
rect 433334 271368 433340 271380
rect 361172 271340 433340 271368
rect 361172 271328 361178 271340
rect 433334 271328 433340 271340
rect 433392 271328 433398 271380
rect 183462 271260 183468 271312
rect 183520 271300 183526 271312
rect 197354 271300 197360 271312
rect 183520 271272 197360 271300
rect 183520 271260 183526 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 209222 271260 209228 271312
rect 209280 271300 209286 271312
rect 264974 271300 264980 271312
rect 209280 271272 264980 271300
rect 209280 271260 209286 271272
rect 264974 271260 264980 271272
rect 265032 271260 265038 271312
rect 343450 271260 343456 271312
rect 343508 271300 343514 271312
rect 360194 271300 360200 271312
rect 343508 271272 360200 271300
rect 343508 271260 343514 271272
rect 360194 271260 360200 271272
rect 360252 271260 360258 271312
rect 368198 271260 368204 271312
rect 368256 271300 368262 271312
rect 440234 271300 440240 271312
rect 368256 271272 440240 271300
rect 368256 271260 368262 271272
rect 440234 271260 440240 271272
rect 440292 271260 440298 271312
rect 503622 271260 503628 271312
rect 503680 271300 503686 271312
rect 517606 271300 517612 271312
rect 503680 271272 517612 271300
rect 503680 271260 503686 271272
rect 517606 271260 517612 271272
rect 517664 271260 517670 271312
rect 113174 271232 113180 271244
rect 108316 271204 113180 271232
rect 113174 271192 113180 271204
rect 113232 271192 113238 271244
rect 207842 271192 207848 271244
rect 207900 271232 207906 271244
rect 260834 271232 260840 271244
rect 207900 271204 260840 271232
rect 207900 271192 207906 271204
rect 260834 271192 260840 271204
rect 260892 271192 260898 271244
rect 280062 271192 280068 271244
rect 280120 271232 280126 271244
rect 357434 271232 357440 271244
rect 280120 271204 357440 271232
rect 280120 271192 280126 271204
rect 357434 271192 357440 271204
rect 357492 271192 357498 271244
rect 366634 271192 366640 271244
rect 366692 271232 366698 271244
rect 434714 271232 434720 271244
rect 366692 271204 434720 271232
rect 366692 271192 366698 271204
rect 434714 271192 434720 271204
rect 434772 271192 434778 271244
rect 110414 271164 110420 271176
rect 106844 271136 110420 271164
rect 110414 271124 110420 271136
rect 110472 271124 110478 271176
rect 183462 271124 183468 271176
rect 183520 271164 183526 271176
rect 201586 271164 201592 271176
rect 183520 271136 201592 271164
rect 183520 271124 183526 271136
rect 201586 271124 201592 271136
rect 201644 271124 201650 271176
rect 206370 271124 206376 271176
rect 206428 271164 206434 271176
rect 258258 271164 258264 271176
rect 206428 271136 258264 271164
rect 206428 271124 206434 271136
rect 258258 271124 258264 271136
rect 258316 271124 258322 271176
rect 277210 271124 277216 271176
rect 277268 271164 277274 271176
rect 356606 271164 356612 271176
rect 277268 271136 356612 271164
rect 277268 271124 277274 271136
rect 356606 271124 356612 271136
rect 356664 271124 356670 271176
rect 369578 271124 369584 271176
rect 369636 271164 369642 271176
rect 416038 271164 416044 271176
rect 369636 271136 416044 271164
rect 369636 271124 369642 271136
rect 416038 271124 416044 271136
rect 416096 271124 416102 271176
rect 503530 271124 503536 271176
rect 503588 271164 503594 271176
rect 517882 271164 517888 271176
rect 503588 271136 517888 271164
rect 503588 271124 503594 271136
rect 517882 271124 517888 271136
rect 517940 271124 517946 271176
rect 107654 271096 107660 271108
rect 105924 271068 107660 271096
rect 107654 271056 107660 271068
rect 107712 271056 107718 271108
rect 202138 271056 202144 271108
rect 202196 271096 202202 271108
rect 252554 271096 252560 271108
rect 202196 271068 252560 271096
rect 202196 271056 202202 271068
rect 252554 271056 252560 271068
rect 252612 271056 252618 271108
rect 379054 271056 379060 271108
rect 379112 271096 379118 271108
rect 418154 271096 418160 271108
rect 379112 271068 418160 271096
rect 379112 271056 379118 271068
rect 418154 271056 418160 271068
rect 418212 271056 418218 271108
rect 54846 270988 54852 271040
rect 54904 271028 54910 271040
rect 88334 271028 88340 271040
rect 54904 271000 88340 271028
rect 54904 270988 54910 271000
rect 88334 270988 88340 271000
rect 88392 270988 88398 271040
rect 106918 270988 106924 271040
rect 106976 271028 106982 271040
rect 113266 271028 113272 271040
rect 106976 271000 113272 271028
rect 106976 270988 106982 271000
rect 113266 270988 113272 271000
rect 113324 270988 113330 271040
rect 206554 270988 206560 271040
rect 206612 271028 206618 271040
rect 255314 271028 255320 271040
rect 206612 271000 255320 271028
rect 206612 270988 206618 271000
rect 255314 270988 255320 271000
rect 255372 270988 255378 271040
rect 376202 270988 376208 271040
rect 376260 271028 376266 271040
rect 412726 271028 412732 271040
rect 376260 271000 412732 271028
rect 376260 270988 376266 271000
rect 412726 270988 412732 271000
rect 412784 270988 412790 271040
rect 46106 270920 46112 270972
rect 46164 270960 46170 270972
rect 77294 270960 77300 270972
rect 46164 270932 77300 270960
rect 46164 270920 46170 270932
rect 77294 270920 77300 270932
rect 77352 270920 77358 270972
rect 214834 270920 214840 270972
rect 214892 270960 214898 270972
rect 247034 270960 247040 270972
rect 214892 270932 247040 270960
rect 214892 270920 214898 270932
rect 247034 270920 247040 270932
rect 247092 270920 247098 270972
rect 374914 270920 374920 270972
rect 374972 270960 374978 270972
rect 409874 270960 409880 270972
rect 374972 270932 409880 270960
rect 374972 270920 374978 270932
rect 409874 270920 409880 270932
rect 409932 270920 409938 270972
rect 43438 270444 43444 270496
rect 43496 270484 43502 270496
rect 129734 270484 129740 270496
rect 43496 270456 129740 270484
rect 43496 270444 43502 270456
rect 129734 270444 129740 270456
rect 129792 270444 129798 270496
rect 196710 270444 196716 270496
rect 196768 270484 196774 270496
rect 197814 270484 197820 270496
rect 196768 270456 197820 270484
rect 196768 270444 196774 270456
rect 197814 270444 197820 270456
rect 197872 270444 197878 270496
rect 211706 270444 211712 270496
rect 211764 270484 211770 270496
rect 212350 270484 212356 270496
rect 211764 270456 212356 270484
rect 211764 270444 211770 270456
rect 212350 270444 212356 270456
rect 212408 270444 212414 270496
rect 213086 270444 213092 270496
rect 213144 270484 213150 270496
rect 213546 270484 213552 270496
rect 213144 270456 213552 270484
rect 213144 270444 213150 270456
rect 213546 270444 213552 270456
rect 213604 270444 213610 270496
rect 220538 270444 220544 270496
rect 220596 270484 220602 270496
rect 248506 270484 248512 270496
rect 220596 270456 248512 270484
rect 220596 270444 220602 270456
rect 248506 270444 248512 270456
rect 248564 270444 248570 270496
rect 411254 270484 411260 270496
rect 379624 270456 411260 270484
rect 50522 270376 50528 270428
rect 50580 270416 50586 270428
rect 84194 270416 84200 270428
rect 50580 270388 84200 270416
rect 50580 270376 50586 270388
rect 84194 270376 84200 270388
rect 84252 270376 84258 270428
rect 220722 270376 220728 270428
rect 220780 270416 220786 270428
rect 247034 270416 247040 270428
rect 220780 270388 247040 270416
rect 220780 270376 220786 270388
rect 247034 270376 247040 270388
rect 247092 270376 247098 270428
rect 377030 270376 377036 270428
rect 377088 270416 377094 270428
rect 378042 270416 378048 270428
rect 377088 270388 378048 270416
rect 377088 270376 377094 270388
rect 378042 270376 378048 270388
rect 378100 270416 378106 270428
rect 379624 270416 379652 270456
rect 411254 270444 411260 270456
rect 411312 270444 411318 270496
rect 378100 270388 379652 270416
rect 378100 270376 378106 270388
rect 380526 270376 380532 270428
rect 380584 270416 380590 270428
rect 411346 270416 411352 270428
rect 380584 270388 411352 270416
rect 380584 270376 380590 270388
rect 411346 270376 411352 270388
rect 411404 270376 411410 270428
rect 81434 270308 81440 270360
rect 81492 270348 81498 270360
rect 107654 270348 107660 270360
rect 81492 270320 107660 270348
rect 81492 270308 81498 270320
rect 107654 270308 107660 270320
rect 107712 270308 107718 270360
rect 218606 270308 218612 270360
rect 218664 270348 218670 270360
rect 219342 270348 219348 270360
rect 218664 270320 219348 270348
rect 218664 270308 218670 270320
rect 219342 270308 219348 270320
rect 219400 270348 219406 270360
rect 252554 270348 252560 270360
rect 219400 270320 252560 270348
rect 219400 270308 219406 270320
rect 252554 270308 252560 270320
rect 252612 270308 252618 270360
rect 370958 270308 370964 270360
rect 371016 270348 371022 270360
rect 401686 270348 401692 270360
rect 371016 270320 401692 270348
rect 371016 270308 371022 270320
rect 401686 270308 401692 270320
rect 401744 270308 401750 270360
rect 80054 270240 80060 270292
rect 80112 270280 80118 270292
rect 109218 270280 109224 270292
rect 80112 270252 109224 270280
rect 80112 270240 80118 270252
rect 109218 270240 109224 270252
rect 109276 270240 109282 270292
rect 212350 270240 212356 270292
rect 212408 270280 212414 270292
rect 245654 270280 245660 270292
rect 212408 270252 245660 270280
rect 212408 270240 212414 270252
rect 245654 270240 245660 270252
rect 245712 270240 245718 270292
rect 379238 270240 379244 270292
rect 379296 270280 379302 270292
rect 379422 270280 379428 270292
rect 379296 270252 379428 270280
rect 379296 270240 379302 270252
rect 379422 270240 379428 270252
rect 379480 270240 379486 270292
rect 404354 270280 404360 270292
rect 379808 270252 404360 270280
rect 63494 270172 63500 270224
rect 63552 270212 63558 270224
rect 92474 270212 92480 270224
rect 63552 270184 92480 270212
rect 63552 270172 63558 270184
rect 92474 270172 92480 270184
rect 92532 270172 92538 270224
rect 219158 270172 219164 270224
rect 219216 270212 219222 270224
rect 251174 270212 251180 270224
rect 219216 270184 251180 270212
rect 219216 270172 219222 270184
rect 251174 270172 251180 270184
rect 251232 270172 251238 270224
rect 376662 270172 376668 270224
rect 376720 270212 376726 270224
rect 379808 270212 379836 270252
rect 404354 270240 404360 270252
rect 404412 270240 404418 270292
rect 376720 270184 379836 270212
rect 376720 270172 376726 270184
rect 379882 270172 379888 270224
rect 379940 270212 379946 270224
rect 405734 270212 405740 270224
rect 379940 270184 405740 270212
rect 379940 270172 379946 270184
rect 405734 270172 405740 270184
rect 405792 270172 405798 270224
rect 51718 270104 51724 270156
rect 51776 270144 51782 270156
rect 54570 270144 54576 270156
rect 51776 270116 54576 270144
rect 51776 270104 51782 270116
rect 54570 270104 54576 270116
rect 54628 270144 54634 270156
rect 84654 270144 84660 270156
rect 54628 270116 84660 270144
rect 54628 270104 54634 270116
rect 84654 270104 84660 270116
rect 84712 270104 84718 270156
rect 216766 270104 216772 270156
rect 216824 270144 216830 270156
rect 219250 270144 219256 270156
rect 216824 270116 219256 270144
rect 216824 270104 216830 270116
rect 219250 270104 219256 270116
rect 219308 270144 219314 270156
rect 251266 270144 251272 270156
rect 219308 270116 251272 270144
rect 219308 270104 219314 270116
rect 251266 270104 251272 270116
rect 251324 270104 251330 270156
rect 373166 270104 373172 270156
rect 373224 270144 373230 270156
rect 398834 270144 398840 270156
rect 373224 270116 398840 270144
rect 373224 270104 373230 270116
rect 398834 270104 398840 270116
rect 398892 270104 398898 270156
rect 57974 270036 57980 270088
rect 58032 270076 58038 270088
rect 91094 270076 91100 270088
rect 58032 270048 91100 270076
rect 58032 270036 58038 270048
rect 91094 270036 91100 270048
rect 91152 270036 91158 270088
rect 213546 270036 213552 270088
rect 213604 270076 213610 270088
rect 244274 270076 244280 270088
rect 213604 270048 244280 270076
rect 213604 270036 213610 270048
rect 244274 270036 244280 270048
rect 244332 270036 244338 270088
rect 373902 270036 373908 270088
rect 373960 270076 373966 270088
rect 374454 270076 374460 270088
rect 373960 270048 374460 270076
rect 373960 270036 373966 270048
rect 374454 270036 374460 270048
rect 374512 270036 374518 270088
rect 375098 270036 375104 270088
rect 375156 270076 375162 270088
rect 400214 270076 400220 270088
rect 375156 270048 400220 270076
rect 375156 270036 375162 270048
rect 400214 270036 400220 270048
rect 400272 270036 400278 270088
rect 53190 269968 53196 270020
rect 53248 270008 53254 270020
rect 58618 270008 58624 270020
rect 53248 269980 58624 270008
rect 53248 269968 53254 269980
rect 58618 269968 58624 269980
rect 58676 269968 58682 270020
rect 77386 269968 77392 270020
rect 77444 270008 77450 270020
rect 110414 270008 110420 270020
rect 77444 269980 110420 270008
rect 77444 269968 77450 269980
rect 110414 269968 110420 269980
rect 110472 269968 110478 270020
rect 220354 269968 220360 270020
rect 220412 270008 220418 270020
rect 249794 270008 249800 270020
rect 220412 269980 249800 270008
rect 220412 269968 220418 269980
rect 249794 269968 249800 269980
rect 249852 269968 249858 270020
rect 370406 269968 370412 270020
rect 370464 270008 370470 270020
rect 373718 270008 373724 270020
rect 370464 269980 373724 270008
rect 370464 269968 370470 269980
rect 373718 269968 373724 269980
rect 373776 270008 373782 270020
rect 397454 270008 397460 270020
rect 373776 269980 397460 270008
rect 373776 269968 373782 269980
rect 397454 269968 397460 269980
rect 397512 269968 397518 270020
rect 55950 269900 55956 269952
rect 56008 269940 56014 269952
rect 88334 269940 88340 269952
rect 56008 269912 88340 269940
rect 56008 269900 56014 269912
rect 88334 269900 88340 269912
rect 88392 269900 88398 269952
rect 220630 269900 220636 269952
rect 220688 269940 220694 269952
rect 262214 269940 262220 269952
rect 220688 269912 262220 269940
rect 220688 269900 220694 269912
rect 262214 269900 262220 269912
rect 262272 269900 262278 269952
rect 371786 269900 371792 269952
rect 371844 269940 371850 269952
rect 373626 269940 373632 269952
rect 371844 269912 373632 269940
rect 371844 269900 371850 269912
rect 373626 269900 373632 269912
rect 373684 269940 373690 269952
rect 403342 269940 403348 269952
rect 373684 269912 403348 269940
rect 373684 269900 373690 269912
rect 403342 269900 403348 269912
rect 403400 269900 403406 269952
rect 57146 269832 57152 269884
rect 57204 269872 57210 269884
rect 89714 269872 89720 269884
rect 57204 269844 89720 269872
rect 57204 269832 57210 269844
rect 89714 269832 89720 269844
rect 89772 269832 89778 269884
rect 115842 269832 115848 269884
rect 115900 269872 115906 269884
rect 197722 269872 197728 269884
rect 115900 269844 197728 269872
rect 115900 269832 115906 269844
rect 197722 269832 197728 269844
rect 197780 269872 197786 269884
rect 201494 269872 201500 269884
rect 197780 269844 201500 269872
rect 197780 269832 197786 269844
rect 201494 269832 201500 269844
rect 201552 269832 201558 269884
rect 220722 269832 220728 269884
rect 220780 269872 220786 269884
rect 265158 269872 265164 269884
rect 220780 269844 265164 269872
rect 220780 269832 220786 269844
rect 265158 269832 265164 269844
rect 265216 269832 265222 269884
rect 374454 269832 374460 269884
rect 374512 269872 374518 269884
rect 407114 269872 407120 269884
rect 374512 269844 407120 269872
rect 374512 269832 374518 269844
rect 407114 269832 407120 269844
rect 407172 269832 407178 269884
rect 51718 269764 51724 269816
rect 51776 269804 51782 269816
rect 85574 269804 85580 269816
rect 51776 269776 85580 269804
rect 51776 269764 51782 269776
rect 85574 269764 85580 269776
rect 85632 269764 85638 269816
rect 113358 269764 113364 269816
rect 113416 269804 113422 269816
rect 196710 269804 196716 269816
rect 113416 269776 196716 269804
rect 113416 269764 113422 269776
rect 196710 269764 196716 269776
rect 196768 269764 196774 269816
rect 217134 269764 217140 269816
rect 217192 269804 217198 269816
rect 218606 269804 218612 269816
rect 217192 269776 218612 269804
rect 217192 269764 217198 269776
rect 218606 269764 218612 269776
rect 218664 269804 218670 269816
rect 266354 269804 266360 269816
rect 218664 269776 266360 269804
rect 218664 269764 218670 269776
rect 266354 269764 266360 269776
rect 266412 269764 266418 269816
rect 372246 269764 372252 269816
rect 372304 269804 372310 269816
rect 375098 269804 375104 269816
rect 372304 269776 375104 269804
rect 372304 269764 372310 269776
rect 375098 269764 375104 269776
rect 375156 269764 375162 269816
rect 379514 269764 379520 269816
rect 379572 269804 379578 269816
rect 413002 269804 413008 269816
rect 379572 269776 413008 269804
rect 379572 269764 379578 269776
rect 413002 269764 413008 269776
rect 413060 269764 413066 269816
rect 205266 269696 205272 269748
rect 205324 269736 205330 269748
rect 209498 269736 209504 269748
rect 205324 269708 209504 269736
rect 205324 269696 205330 269708
rect 209498 269696 209504 269708
rect 209556 269736 209562 269748
rect 237374 269736 237380 269748
rect 209556 269708 237380 269736
rect 209556 269696 209562 269708
rect 237374 269696 237380 269708
rect 237432 269696 237438 269748
rect 376478 269696 376484 269748
rect 376536 269736 376542 269748
rect 377122 269736 377128 269748
rect 376536 269708 377128 269736
rect 376536 269696 376542 269708
rect 377122 269696 377128 269708
rect 377180 269736 377186 269748
rect 391934 269736 391940 269748
rect 377180 269708 391940 269736
rect 377180 269696 377186 269708
rect 391934 269696 391940 269708
rect 391992 269696 391998 269748
rect 212258 269628 212264 269680
rect 212316 269668 212322 269680
rect 271874 269668 271880 269680
rect 212316 269640 271880 269668
rect 212316 269628 212322 269640
rect 271874 269628 271880 269640
rect 271932 269628 271938 269680
rect 375098 269628 375104 269680
rect 375156 269668 375162 269680
rect 380158 269668 380164 269680
rect 375156 269640 380164 269668
rect 375156 269628 375162 269640
rect 380158 269628 380164 269640
rect 380216 269628 380222 269680
rect 216674 269560 216680 269612
rect 216732 269600 216738 269612
rect 217962 269600 217968 269612
rect 216732 269572 217968 269600
rect 216732 269560 216738 269572
rect 217962 269560 217968 269572
rect 218020 269600 218026 269612
rect 263594 269600 263600 269612
rect 218020 269572 263600 269600
rect 218020 269560 218026 269572
rect 263594 269560 263600 269572
rect 263652 269560 263658 269612
rect 378410 269560 378416 269612
rect 378468 269600 378474 269612
rect 379606 269600 379612 269612
rect 378468 269572 379612 269600
rect 378468 269560 378474 269572
rect 379606 269560 379612 269572
rect 379664 269600 379670 269612
rect 380526 269600 380532 269612
rect 379664 269572 380532 269600
rect 379664 269560 379670 269572
rect 380526 269560 380532 269572
rect 380584 269560 380590 269612
rect 214374 269492 214380 269544
rect 214432 269532 214438 269544
rect 219526 269532 219532 269544
rect 214432 269504 219532 269532
rect 214432 269492 214438 269504
rect 219526 269492 219532 269504
rect 219584 269532 219590 269544
rect 220538 269532 220544 269544
rect 219584 269504 220544 269532
rect 219584 269492 219590 269504
rect 220538 269492 220544 269504
rect 220596 269492 220602 269544
rect 378594 269492 378600 269544
rect 378652 269532 378658 269544
rect 379882 269532 379888 269544
rect 378652 269504 379888 269532
rect 378652 269492 378658 269504
rect 379882 269492 379888 269504
rect 379940 269492 379946 269544
rect 215846 269424 215852 269476
rect 215904 269464 215910 269476
rect 219710 269464 219716 269476
rect 215904 269436 219716 269464
rect 215904 269424 215910 269436
rect 219710 269424 219716 269436
rect 219768 269464 219774 269476
rect 220354 269464 220360 269476
rect 219768 269436 220360 269464
rect 219768 269424 219774 269436
rect 220354 269424 220360 269436
rect 220412 269424 220418 269476
rect 218514 269356 218520 269408
rect 218572 269396 218578 269408
rect 219618 269396 219624 269408
rect 218572 269368 219624 269396
rect 218572 269356 218578 269368
rect 219618 269356 219624 269368
rect 219676 269396 219682 269408
rect 220722 269396 220728 269408
rect 219676 269368 220728 269396
rect 219676 269356 219682 269368
rect 220722 269356 220728 269368
rect 220780 269356 220786 269408
rect 217226 269220 217232 269272
rect 217284 269260 217290 269272
rect 219434 269260 219440 269272
rect 217284 269232 219440 269260
rect 217284 269220 217290 269232
rect 219434 269220 219440 269232
rect 219492 269260 219498 269272
rect 220630 269260 220636 269272
rect 219492 269232 220636 269260
rect 219492 269220 219498 269232
rect 220630 269220 220636 269232
rect 220688 269220 220694 269272
rect 370774 269084 370780 269136
rect 370832 269124 370838 269136
rect 373166 269124 373172 269136
rect 370832 269096 373172 269124
rect 370832 269084 370838 269096
rect 373166 269084 373172 269096
rect 373224 269084 373230 269136
rect 46750 269016 46756 269068
rect 46808 269056 46814 269068
rect 51718 269056 51724 269068
rect 46808 269028 51724 269056
rect 46808 269016 46814 269028
rect 51718 269016 51724 269028
rect 51776 269016 51782 269068
rect 210326 269016 210332 269068
rect 210384 269056 210390 269068
rect 210878 269056 210884 269068
rect 210384 269028 210884 269056
rect 210384 269016 210390 269028
rect 210878 269016 210884 269028
rect 210936 269016 210942 269068
rect 213270 269016 213276 269068
rect 213328 269056 213334 269068
rect 216122 269056 216128 269068
rect 213328 269028 216128 269056
rect 213328 269016 213334 269028
rect 216122 269016 216128 269028
rect 216180 269016 216186 269068
rect 216398 269016 216404 269068
rect 216456 269056 216462 269068
rect 219066 269056 219072 269068
rect 216456 269028 219072 269056
rect 216456 269016 216462 269028
rect 219066 269016 219072 269028
rect 219124 269016 219130 269068
rect 267918 269056 267924 269068
rect 219406 269028 267924 269056
rect 43714 268948 43720 269000
rect 43772 268988 43778 269000
rect 57974 268988 57980 269000
rect 43772 268960 57980 268988
rect 43772 268948 43778 268960
rect 57974 268948 57980 268960
rect 58032 268948 58038 269000
rect 215754 268948 215760 269000
rect 215812 268988 215818 269000
rect 218514 268988 218520 269000
rect 215812 268960 218520 268988
rect 215812 268948 215818 268960
rect 218514 268948 218520 268960
rect 218572 268948 218578 269000
rect 45462 268880 45468 268932
rect 45520 268920 45526 268932
rect 57146 268920 57152 268932
rect 45520 268892 57152 268920
rect 45520 268880 45526 268892
rect 57146 268880 57152 268892
rect 57204 268880 57210 268932
rect 215018 268880 215024 268932
rect 215076 268920 215082 268932
rect 217134 268920 217140 268932
rect 215076 268892 217140 268920
rect 215076 268880 215082 268892
rect 217134 268880 217140 268892
rect 217192 268880 217198 268932
rect 48222 268812 48228 268864
rect 48280 268852 48286 268864
rect 55950 268852 55956 268864
rect 48280 268824 55956 268852
rect 48280 268812 48286 268824
rect 55950 268812 55956 268824
rect 56008 268812 56014 268864
rect 210878 268812 210884 268864
rect 210936 268852 210942 268864
rect 219406 268852 219434 269028
rect 267918 269016 267924 269028
rect 267976 269016 267982 269068
rect 374362 269016 374368 269068
rect 374420 269056 374426 269068
rect 375926 269056 375932 269068
rect 374420 269028 375932 269056
rect 374420 269016 374426 269028
rect 375926 269016 375932 269028
rect 375984 269056 375990 269068
rect 416774 269056 416780 269068
rect 375984 269028 416780 269056
rect 375984 269016 375990 269028
rect 416774 269016 416780 269028
rect 416832 269016 416838 269068
rect 219802 268948 219808 269000
rect 219860 268988 219866 269000
rect 253934 268988 253940 269000
rect 219860 268960 253940 268988
rect 219860 268948 219866 268960
rect 253934 268948 253940 268960
rect 253992 268948 253998 269000
rect 379974 268948 379980 269000
rect 380032 268988 380038 269000
rect 414014 268988 414020 269000
rect 380032 268960 414020 268988
rect 380032 268948 380038 268960
rect 414014 268948 414020 268960
rect 414072 268948 414078 269000
rect 232498 268880 232504 268932
rect 232556 268920 232562 268932
rect 259454 268920 259460 268932
rect 232556 268892 259460 268920
rect 232556 268880 232562 268892
rect 259454 268880 259460 268892
rect 259512 268880 259518 268932
rect 387886 268880 387892 268932
rect 387944 268920 387950 268932
rect 420914 268920 420920 268932
rect 387944 268892 420920 268920
rect 387944 268880 387950 268892
rect 420914 268880 420920 268892
rect 420972 268880 420978 268932
rect 210936 268824 219434 268852
rect 210936 268812 210942 268824
rect 231118 268812 231124 268864
rect 231176 268852 231182 268864
rect 259546 268852 259552 268864
rect 231176 268824 259552 268852
rect 231176 268812 231182 268824
rect 259546 268812 259552 268824
rect 259604 268812 259610 268864
rect 377490 268812 377496 268864
rect 377548 268852 377554 268864
rect 377950 268852 377956 268864
rect 377548 268824 377956 268852
rect 377548 268812 377554 268824
rect 377950 268812 377956 268824
rect 378008 268852 378014 268864
rect 408494 268852 408500 268864
rect 378008 268824 408500 268852
rect 378008 268812 378014 268824
rect 408494 268812 408500 268824
rect 408552 268812 408558 268864
rect 45278 268744 45284 268796
rect 45336 268784 45342 268796
rect 147674 268784 147680 268796
rect 45336 268756 147680 268784
rect 45336 268744 45342 268756
rect 147674 268744 147680 268756
rect 147732 268744 147738 268796
rect 216490 268744 216496 268796
rect 216548 268784 216554 268796
rect 229094 268784 229100 268796
rect 216548 268756 229100 268784
rect 216548 268744 216554 268756
rect 229094 268744 229100 268756
rect 229152 268784 229158 268796
rect 260834 268784 260840 268796
rect 229152 268756 260840 268784
rect 229152 268744 229158 268756
rect 260834 268744 260840 268756
rect 260892 268744 260898 268796
rect 379146 268744 379152 268796
rect 379204 268784 379210 268796
rect 379330 268784 379336 268796
rect 379204 268756 379336 268784
rect 379204 268744 379210 268756
rect 379330 268744 379336 268756
rect 379388 268784 379394 268796
rect 409874 268784 409880 268796
rect 379388 268756 409880 268784
rect 379388 268744 379394 268756
rect 409874 268744 409880 268756
rect 409932 268744 409938 268796
rect 216122 268676 216128 268728
rect 216180 268716 216186 268728
rect 255314 268716 255320 268728
rect 216180 268688 255320 268716
rect 216180 268676 216186 268688
rect 255314 268676 255320 268688
rect 255372 268676 255378 268728
rect 390554 268676 390560 268728
rect 390612 268716 390618 268728
rect 419534 268716 419540 268728
rect 390612 268688 419540 268716
rect 390612 268676 390618 268688
rect 419534 268676 419540 268688
rect 419592 268676 419598 268728
rect 49234 268608 49240 268660
rect 49292 268648 49298 268660
rect 63494 268648 63500 268660
rect 49292 268620 63500 268648
rect 49292 268608 49298 268620
rect 63494 268608 63500 268620
rect 63552 268608 63558 268660
rect 213730 268608 213736 268660
rect 213788 268648 213794 268660
rect 216490 268648 216496 268660
rect 213788 268620 216496 268648
rect 213788 268608 213794 268620
rect 216490 268608 216496 268620
rect 216548 268608 216554 268660
rect 217134 268608 217140 268660
rect 217192 268648 217198 268660
rect 256694 268648 256700 268660
rect 217192 268620 256700 268648
rect 217192 268608 217198 268620
rect 256694 268608 256700 268620
rect 256752 268608 256758 268660
rect 391934 268608 391940 268660
rect 391992 268648 391998 268660
rect 418154 268648 418160 268660
rect 391992 268620 418160 268648
rect 391992 268608 391998 268620
rect 418154 268608 418160 268620
rect 418212 268608 418218 268660
rect 49050 268540 49056 268592
rect 49108 268580 49114 268592
rect 80054 268580 80060 268592
rect 49108 268552 80060 268580
rect 49108 268540 49114 268552
rect 80054 268540 80060 268552
rect 80112 268540 80118 268592
rect 218514 268540 218520 268592
rect 218572 268580 218578 268592
rect 258074 268580 258080 268592
rect 218572 268552 258080 268580
rect 218572 268540 218578 268552
rect 258074 268540 258080 268552
rect 258132 268540 258138 268592
rect 42334 268472 42340 268524
rect 42392 268512 42398 268524
rect 46658 268512 46664 268524
rect 42392 268484 46664 268512
rect 42392 268472 42398 268484
rect 46658 268472 46664 268484
rect 46716 268512 46722 268524
rect 81434 268512 81440 268524
rect 46716 268484 81440 268512
rect 46716 268472 46722 268484
rect 81434 268472 81440 268484
rect 81492 268472 81498 268524
rect 208210 268472 208216 268524
rect 208268 268512 208274 268524
rect 213638 268512 213644 268524
rect 208268 268484 213644 268512
rect 208268 268472 208274 268484
rect 213638 268472 213644 268484
rect 213696 268512 213702 268524
rect 269114 268512 269120 268524
rect 213696 268484 269120 268512
rect 213696 268472 213702 268484
rect 269114 268472 269120 268484
rect 269172 268472 269178 268524
rect 43806 268404 43812 268456
rect 43864 268444 43870 268456
rect 49234 268444 49240 268456
rect 43864 268416 49240 268444
rect 43864 268404 43870 268416
rect 49234 268404 49240 268416
rect 49292 268404 49298 268456
rect 58710 268404 58716 268456
rect 58768 268444 58774 268456
rect 104894 268444 104900 268456
rect 58768 268416 104900 268444
rect 58768 268404 58774 268416
rect 104894 268404 104900 268416
rect 104952 268404 104958 268456
rect 209590 268404 209596 268456
rect 209648 268444 209654 268456
rect 212166 268444 212172 268456
rect 209648 268416 212172 268444
rect 209648 268404 209654 268416
rect 212166 268404 212172 268416
rect 212224 268444 212230 268456
rect 270494 268444 270500 268456
rect 212224 268416 270500 268444
rect 212224 268404 212230 268416
rect 270494 268404 270500 268416
rect 270552 268404 270558 268456
rect 43530 268336 43536 268388
rect 43588 268376 43594 268388
rect 49050 268376 49056 268388
rect 43588 268348 49056 268376
rect 43588 268336 43594 268348
rect 49050 268336 49056 268348
rect 49108 268336 49114 268388
rect 50430 268336 50436 268388
rect 50488 268376 50494 268388
rect 98086 268376 98092 268388
rect 50488 268348 98092 268376
rect 50488 268336 50494 268348
rect 98086 268336 98092 268348
rect 98144 268336 98150 268388
rect 206830 268336 206836 268388
rect 206888 268376 206894 268388
rect 213454 268376 213460 268388
rect 206888 268348 213460 268376
rect 206888 268336 206894 268348
rect 213454 268336 213460 268348
rect 213512 268376 213518 268388
rect 273162 268376 273168 268388
rect 213512 268348 273168 268376
rect 213512 268336 213518 268348
rect 273162 268336 273168 268348
rect 273220 268336 273226 268388
rect 374546 268336 374552 268388
rect 374604 268376 374610 268388
rect 376570 268376 376576 268388
rect 374604 268348 376576 268376
rect 374604 268336 374610 268348
rect 376570 268336 376576 268348
rect 376628 268376 376634 268388
rect 402974 268376 402980 268388
rect 376628 268348 402980 268376
rect 376628 268336 376634 268348
rect 402974 268336 402980 268348
rect 403032 268336 403038 268388
rect 216490 268268 216496 268320
rect 216548 268308 216554 268320
rect 242894 268308 242900 268320
rect 216548 268280 242900 268308
rect 216548 268268 216554 268280
rect 242894 268268 242900 268280
rect 242952 268268 242958 268320
rect 219066 268200 219072 268252
rect 219124 268240 219130 268252
rect 244366 268240 244372 268252
rect 219124 268212 244372 268240
rect 219124 268200 219130 268212
rect 244366 268200 244372 268212
rect 244424 268200 244430 268252
rect 45370 267656 45376 267708
rect 45428 267696 45434 267708
rect 58066 267696 58072 267708
rect 45428 267668 58072 267696
rect 45428 267656 45434 267668
rect 58066 267656 58072 267668
rect 58124 267656 58130 267708
rect 213362 267656 213368 267708
rect 213420 267696 213426 267708
rect 274634 267696 274640 267708
rect 213420 267668 274640 267696
rect 213420 267656 213426 267668
rect 274634 267656 274640 267668
rect 274692 267656 274698 267708
rect 377674 267656 377680 267708
rect 377732 267696 377738 267708
rect 437474 267696 437480 267708
rect 377732 267668 437480 267696
rect 377732 267656 377738 267668
rect 437474 267656 437480 267668
rect 437532 267656 437538 267708
rect 216306 267588 216312 267640
rect 216364 267628 216370 267640
rect 277394 267628 277400 267640
rect 216364 267600 277400 267628
rect 216364 267588 216370 267600
rect 277394 267588 277400 267600
rect 277452 267588 277458 267640
rect 380066 267588 380072 267640
rect 380124 267628 380130 267640
rect 438854 267628 438860 267640
rect 380124 267600 438860 267628
rect 380124 267588 380130 267600
rect 438854 267588 438860 267600
rect 438912 267588 438918 267640
rect 375282 267520 375288 267572
rect 375340 267560 375346 267572
rect 433334 267560 433340 267572
rect 375340 267532 433340 267560
rect 375340 267520 375346 267532
rect 433334 267520 433340 267532
rect 433392 267520 433398 267572
rect 58066 267180 58072 267232
rect 58124 267220 58130 267232
rect 58710 267220 58716 267232
rect 58124 267192 58716 267220
rect 58124 267180 58130 267192
rect 58710 267180 58716 267192
rect 58768 267180 58774 267232
rect 379054 266364 379060 266416
rect 379112 266404 379118 266416
rect 380066 266404 380072 266416
rect 379112 266376 380072 266404
rect 379112 266364 379118 266376
rect 380066 266364 380072 266376
rect 380124 266364 380130 266416
rect 356974 253960 356980 253972
rect 356440 253932 356980 253960
rect 191742 253852 191748 253904
rect 191800 253892 191806 253904
rect 201402 253892 201408 253904
rect 191800 253864 201408 253892
rect 191800 253852 191806 253864
rect 201402 253852 201408 253864
rect 201460 253892 201466 253904
rect 202874 253892 202880 253904
rect 201460 253864 202880 253892
rect 201460 253852 201466 253864
rect 202874 253852 202880 253864
rect 202932 253852 202938 253904
rect 339402 253852 339408 253904
rect 339460 253892 339466 253904
rect 356440 253892 356468 253932
rect 356974 253920 356980 253932
rect 357032 253960 357038 253972
rect 357802 253960 357808 253972
rect 357032 253932 357808 253960
rect 357032 253920 357038 253932
rect 357802 253920 357808 253932
rect 357860 253920 357866 253972
rect 339460 253864 356468 253892
rect 339460 253852 339466 253864
rect 500862 253308 500868 253360
rect 500920 253348 500926 253360
rect 517698 253348 517704 253360
rect 500920 253320 517704 253348
rect 500920 253308 500926 253320
rect 517698 253308 517704 253320
rect 517756 253308 517762 253360
rect 180518 253240 180524 253292
rect 180576 253280 180582 253292
rect 197538 253280 197544 253292
rect 180576 253252 197544 253280
rect 180576 253240 180582 253252
rect 197538 253240 197544 253252
rect 197596 253240 197602 253292
rect 340782 253240 340788 253292
rect 340840 253280 340846 253292
rect 357526 253280 357532 253292
rect 340840 253252 357532 253280
rect 340840 253240 340846 253252
rect 357526 253240 357532 253252
rect 357584 253280 357590 253292
rect 357710 253280 357716 253292
rect 357584 253252 357716 253280
rect 357584 253240 357590 253252
rect 357710 253240 357716 253252
rect 357768 253240 357774 253292
rect 499206 253240 499212 253292
rect 499264 253280 499270 253292
rect 517790 253280 517796 253292
rect 499264 253252 517796 253280
rect 499264 253240 499270 253252
rect 517790 253240 517796 253252
rect 517848 253240 517854 253292
rect 179322 253172 179328 253224
rect 179380 253212 179386 253224
rect 197446 253212 197452 253224
rect 179380 253184 197452 253212
rect 179380 253172 179386 253184
rect 197446 253172 197452 253184
rect 197504 253212 197510 253224
rect 197630 253212 197636 253224
rect 197504 253184 197636 253212
rect 197504 253172 197510 253184
rect 197630 253172 197636 253184
rect 197688 253172 197694 253224
rect 351822 253172 351828 253224
rect 351880 253212 351886 253224
rect 358078 253212 358084 253224
rect 351880 253184 358084 253212
rect 351880 253172 351886 253184
rect 358078 253172 358084 253184
rect 358136 253172 358142 253224
rect 517698 253172 517704 253224
rect 517756 253212 517762 253224
rect 517974 253212 517980 253224
rect 517756 253184 517980 253212
rect 517756 253172 517762 253184
rect 517974 253172 517980 253184
rect 518032 253172 518038 253224
rect 510890 252560 510896 252612
rect 510948 252600 510954 252612
rect 517514 252600 517520 252612
rect 510948 252572 517520 252600
rect 510948 252560 510954 252572
rect 517514 252560 517520 252572
rect 517572 252560 517578 252612
rect 214466 252492 214472 252544
rect 214524 252532 214530 252544
rect 231118 252532 231124 252544
rect 214524 252504 231124 252532
rect 214524 252492 214530 252504
rect 231118 252492 231124 252504
rect 231176 252492 231182 252544
rect 375190 252492 375196 252544
rect 375248 252532 375254 252544
rect 377674 252532 377680 252544
rect 375248 252504 377680 252532
rect 375248 252492 375254 252504
rect 377674 252492 377680 252504
rect 377732 252532 377738 252544
rect 396718 252532 396724 252544
rect 377732 252504 396724 252532
rect 377732 252492 377738 252504
rect 396718 252492 396724 252504
rect 396776 252492 396782 252544
rect 217962 252424 217968 252476
rect 218020 252464 218026 252476
rect 232498 252464 232504 252476
rect 218020 252436 232504 252464
rect 218020 252424 218026 252436
rect 232498 252424 232504 252436
rect 232556 252424 232562 252476
rect 368382 252424 368388 252476
rect 368440 252464 368446 252476
rect 376202 252464 376208 252476
rect 368440 252436 376208 252464
rect 368440 252424 368446 252436
rect 376202 252424 376208 252436
rect 376260 252424 376266 252476
rect 58618 252084 58624 252136
rect 58676 252124 58682 252136
rect 60826 252124 60832 252136
rect 58676 252096 60832 252124
rect 58676 252084 58682 252096
rect 60826 252084 60832 252096
rect 60884 252084 60890 252136
rect 375926 252016 375932 252068
rect 375984 252056 375990 252068
rect 376202 252056 376208 252068
rect 375984 252028 376208 252056
rect 375984 252016 375990 252028
rect 376202 252016 376208 252028
rect 376260 252056 376266 252068
rect 427078 252056 427084 252068
rect 376260 252028 427084 252056
rect 376260 252016 376266 252028
rect 427078 252016 427084 252028
rect 427136 252016 427142 252068
rect 54386 251948 54392 252000
rect 54444 251988 54450 252000
rect 60918 251988 60924 252000
rect 54444 251960 60924 251988
rect 54444 251948 54450 251960
rect 60918 251948 60924 251960
rect 60976 251948 60982 252000
rect 369670 251948 369676 252000
rect 369728 251988 369734 252000
rect 372522 251988 372528 252000
rect 369728 251960 372528 251988
rect 369728 251948 369734 251960
rect 372522 251948 372528 251960
rect 372580 251988 372586 252000
rect 425698 251988 425704 252000
rect 372580 251960 425704 251988
rect 372580 251948 372586 251960
rect 425698 251948 425704 251960
rect 425756 251948 425762 252000
rect 54478 251880 54484 251932
rect 54536 251920 54542 251932
rect 61102 251920 61108 251932
rect 54536 251892 61108 251920
rect 54536 251880 54542 251892
rect 61102 251880 61108 251892
rect 61160 251880 61166 251932
rect 372338 251880 372344 251932
rect 372396 251920 372402 251932
rect 373534 251920 373540 251932
rect 372396 251892 373540 251920
rect 372396 251880 372402 251892
rect 373534 251880 373540 251892
rect 373592 251920 373598 251932
rect 429194 251920 429200 251932
rect 373592 251892 429200 251920
rect 373592 251880 373598 251892
rect 429194 251880 429200 251892
rect 429252 251880 429258 251932
rect 52454 251812 52460 251864
rect 52512 251852 52518 251864
rect 106918 251852 106924 251864
rect 52512 251824 106924 251852
rect 52512 251812 52518 251824
rect 106918 251812 106924 251824
rect 106976 251812 106982 251864
rect 214834 251812 214840 251864
rect 214892 251852 214898 251864
rect 229094 251852 229100 251864
rect 214892 251824 229100 251852
rect 214892 251812 214898 251824
rect 229094 251812 229100 251824
rect 229152 251812 229158 251864
rect 375190 251812 375196 251864
rect 375248 251852 375254 251864
rect 431954 251852 431960 251864
rect 375248 251824 431960 251852
rect 375248 251812 375254 251824
rect 431954 251812 431960 251824
rect 432012 251812 432018 251864
rect 58710 251744 58716 251796
rect 58768 251784 58774 251796
rect 61010 251784 61016 251796
rect 58768 251756 61016 251784
rect 58768 251744 58774 251756
rect 61010 251744 61016 251756
rect 61068 251744 61074 251796
rect 56962 251336 56968 251388
rect 57020 251376 57026 251388
rect 62114 251376 62120 251388
rect 57020 251348 62120 251376
rect 57020 251336 57026 251348
rect 62114 251336 62120 251348
rect 62172 251336 62178 251388
rect 46842 251132 46848 251184
rect 46900 251172 46906 251184
rect 52454 251172 52460 251184
rect 46900 251144 52460 251172
rect 46900 251132 46906 251144
rect 52454 251132 52460 251144
rect 52512 251172 52518 251184
rect 53006 251172 53012 251184
rect 52512 251144 53012 251172
rect 52512 251132 52518 251144
rect 53006 251132 53012 251144
rect 53064 251132 53070 251184
rect 372430 251132 372436 251184
rect 372488 251172 372494 251184
rect 374546 251172 374552 251184
rect 372488 251144 374552 251172
rect 372488 251132 372494 251144
rect 374546 251132 374552 251144
rect 374604 251172 374610 251184
rect 375190 251172 375196 251184
rect 374604 251144 375196 251172
rect 374604 251132 374610 251144
rect 375190 251132 375196 251144
rect 375248 251132 375254 251184
rect 519078 183540 519084 183592
rect 519136 183580 519142 183592
rect 520182 183580 520188 183592
rect 519136 183552 520188 183580
rect 519136 183540 519142 183552
rect 520182 183540 520188 183552
rect 520240 183580 520246 183592
rect 580258 183580 580264 183592
rect 520240 183552 580264 183580
rect 520240 183540 520246 183552
rect 580258 183540 580264 183552
rect 580316 183540 580322 183592
rect 520090 183472 520096 183524
rect 520148 183512 520154 183524
rect 580350 183512 580356 183524
rect 520148 183484 580356 183512
rect 520148 183472 520154 183484
rect 580350 183472 580356 183484
rect 580408 183472 580414 183524
rect 216858 178168 216864 178220
rect 216916 178168 216922 178220
rect 216876 178016 216904 178168
rect 204898 177964 204904 178016
rect 204956 178004 204962 178016
rect 216766 178004 216772 178016
rect 204956 177976 216772 178004
rect 204956 177964 204962 177976
rect 216766 177964 216772 177976
rect 216824 177964 216830 178016
rect 216858 177964 216864 178016
rect 216916 177964 216922 178016
rect 365254 177964 365260 178016
rect 365312 178004 365318 178016
rect 376938 178004 376944 178016
rect 365312 177976 376944 178004
rect 365312 177964 365318 177976
rect 376938 177964 376944 177976
rect 376996 177964 377002 178016
rect 202874 176604 202880 176656
rect 202932 176644 202938 176656
rect 216674 176644 216680 176656
rect 202932 176616 216680 176644
rect 202932 176604 202938 176616
rect 216674 176604 216680 176616
rect 216732 176604 216738 176656
rect 202138 176128 202144 176180
rect 202196 176168 202202 176180
rect 202874 176168 202880 176180
rect 202196 176140 202880 176168
rect 202196 176128 202202 176140
rect 202874 176128 202880 176140
rect 202932 176128 202938 176180
rect 358078 175924 358084 175976
rect 358136 175964 358142 175976
rect 376938 175964 376944 175976
rect 358136 175936 376944 175964
rect 358136 175924 358142 175936
rect 376938 175924 376944 175936
rect 376996 175924 377002 175976
rect 43990 175176 43996 175228
rect 44048 175216 44054 175228
rect 57054 175216 57060 175228
rect 44048 175188 57060 175216
rect 44048 175176 44054 175188
rect 57054 175176 57060 175188
rect 57112 175176 57118 175228
rect 207750 175176 207756 175228
rect 207808 175216 207814 175228
rect 217042 175216 217048 175228
rect 207808 175188 217048 175216
rect 207808 175176 207814 175188
rect 217042 175176 217048 175188
rect 217100 175176 217106 175228
rect 365070 175176 365076 175228
rect 365128 175216 365134 175228
rect 376938 175216 376944 175228
rect 365128 175188 376944 175216
rect 365128 175176 365134 175188
rect 376938 175176 376944 175188
rect 376996 175176 377002 175228
rect 216766 175108 216772 175160
rect 216824 175148 216830 175160
rect 216950 175148 216956 175160
rect 216824 175120 216956 175148
rect 216824 175108 216830 175120
rect 216950 175108 216956 175120
rect 217008 175108 217014 175160
rect 49418 166948 49424 167000
rect 49476 166988 49482 167000
rect 98454 166988 98460 167000
rect 49476 166960 98460 166988
rect 49476 166948 49482 166960
rect 98454 166948 98460 166960
rect 98512 166948 98518 167000
rect 197446 166948 197452 167000
rect 197504 166988 197510 167000
rect 201586 166988 201592 167000
rect 197504 166960 201592 166988
rect 197504 166948 197510 166960
rect 201586 166948 201592 166960
rect 201644 166948 201650 167000
rect 373258 166948 373264 167000
rect 373316 166988 373322 167000
rect 421006 166988 421012 167000
rect 373316 166960 421012 166988
rect 373316 166948 373322 166960
rect 421006 166948 421012 166960
rect 421064 166948 421070 167000
rect 50798 166880 50804 166932
rect 50856 166920 50862 166932
rect 101030 166920 101036 166932
rect 50856 166892 101036 166920
rect 50856 166880 50862 166892
rect 101030 166880 101036 166892
rect 101088 166880 101094 166932
rect 362402 166880 362408 166932
rect 362460 166920 362466 166932
rect 423398 166920 423404 166932
rect 362460 166892 423404 166920
rect 362460 166880 362466 166892
rect 423398 166880 423404 166892
rect 423456 166880 423462 166932
rect 51994 166812 52000 166864
rect 52052 166852 52058 166864
rect 105814 166852 105820 166864
rect 52052 166824 105820 166852
rect 52052 166812 52058 166824
rect 105814 166812 105820 166824
rect 105872 166812 105878 166864
rect 358262 166812 358268 166864
rect 358320 166852 358326 166864
rect 418430 166852 418436 166864
rect 358320 166824 418436 166852
rect 358320 166812 358326 166824
rect 418430 166812 418436 166824
rect 418488 166812 418494 166864
rect 53558 166744 53564 166796
rect 53616 166784 53622 166796
rect 108206 166784 108212 166796
rect 53616 166756 108212 166784
rect 53616 166744 53622 166756
rect 108206 166744 108212 166756
rect 108264 166744 108270 166796
rect 210878 166744 210884 166796
rect 210936 166784 210942 166796
rect 220814 166784 220820 166796
rect 210936 166756 220820 166784
rect 210936 166744 210942 166756
rect 220814 166744 220820 166756
rect 220872 166744 220878 166796
rect 363966 166744 363972 166796
rect 364024 166784 364030 166796
rect 428182 166784 428188 166796
rect 364024 166756 428188 166784
rect 364024 166744 364030 166756
rect 428182 166744 428188 166756
rect 428240 166744 428246 166796
rect 56410 166676 56416 166728
rect 56468 166716 56474 166728
rect 138474 166716 138480 166728
rect 56468 166688 138480 166716
rect 56468 166676 56474 166688
rect 138474 166676 138480 166688
rect 138532 166676 138538 166728
rect 214650 166676 214656 166728
rect 214708 166716 214714 166728
rect 260926 166716 260932 166728
rect 214708 166688 260932 166716
rect 214708 166676 214714 166688
rect 260926 166676 260932 166688
rect 260984 166676 260990 166728
rect 356790 166676 356796 166728
rect 356848 166716 356854 166728
rect 445846 166716 445852 166728
rect 356848 166688 445852 166716
rect 356848 166676 356854 166688
rect 445846 166676 445852 166688
rect 445904 166676 445910 166728
rect 58986 166608 58992 166660
rect 59044 166648 59050 166660
rect 140866 166648 140872 166660
rect 59044 166620 140872 166648
rect 59044 166608 59050 166620
rect 140866 166608 140872 166620
rect 140924 166608 140930 166660
rect 203610 166608 203616 166660
rect 203668 166648 203674 166660
rect 265894 166648 265900 166660
rect 203668 166620 265900 166648
rect 203668 166608 203674 166620
rect 265894 166608 265900 166620
rect 265952 166608 265958 166660
rect 372062 166608 372068 166660
rect 372120 166648 372126 166660
rect 470962 166648 470968 166660
rect 372120 166620 470968 166648
rect 372120 166608 372126 166620
rect 470962 166608 470968 166620
rect 471020 166608 471026 166660
rect 59998 166540 60004 166592
rect 60056 166580 60062 166592
rect 145926 166580 145932 166592
rect 60056 166552 145932 166580
rect 60056 166540 60062 166552
rect 145926 166540 145932 166552
rect 145984 166540 145990 166592
rect 210602 166540 210608 166592
rect 210660 166580 210666 166592
rect 293402 166580 293408 166592
rect 210660 166552 293408 166580
rect 210660 166540 210666 166552
rect 293402 166540 293408 166552
rect 293460 166540 293466 166592
rect 373442 166540 373448 166592
rect 373500 166580 373506 166592
rect 475838 166580 475844 166592
rect 373500 166552 475844 166580
rect 373500 166540 373506 166552
rect 475838 166540 475844 166552
rect 475896 166540 475902 166592
rect 59078 166472 59084 166524
rect 59136 166512 59142 166524
rect 148502 166512 148508 166524
rect 59136 166484 148508 166512
rect 59136 166472 59142 166484
rect 148502 166472 148508 166484
rect 148560 166472 148566 166524
rect 203518 166472 203524 166524
rect 203576 166512 203582 166524
rect 285950 166512 285956 166524
rect 203576 166484 285956 166512
rect 203576 166472 203582 166484
rect 285950 166472 285956 166484
rect 286008 166472 286014 166524
rect 367922 166472 367928 166524
rect 367980 166512 367986 166524
rect 478414 166512 478420 166524
rect 367980 166484 478420 166512
rect 367980 166472 367986 166484
rect 478414 166472 478420 166484
rect 478472 166472 478478 166524
rect 58894 166404 58900 166456
rect 58952 166444 58958 166456
rect 153286 166444 153292 166456
rect 58952 166416 153292 166444
rect 58952 166404 58958 166416
rect 153286 166404 153292 166416
rect 153344 166404 153350 166456
rect 203702 166404 203708 166456
rect 203760 166444 203766 166456
rect 288250 166444 288256 166456
rect 203760 166416 288256 166444
rect 203760 166404 203766 166416
rect 288250 166404 288256 166416
rect 288308 166404 288314 166456
rect 365162 166404 365168 166456
rect 365220 166444 365226 166456
rect 480898 166444 480904 166456
rect 365220 166416 480904 166444
rect 365220 166404 365226 166416
rect 480898 166404 480904 166416
rect 480956 166404 480962 166456
rect 43898 166336 43904 166388
rect 43956 166376 43962 166388
rect 163314 166376 163320 166388
rect 43956 166348 163320 166376
rect 43956 166336 43962 166348
rect 163314 166336 163320 166348
rect 163372 166336 163378 166388
rect 209130 166336 209136 166388
rect 209188 166376 209194 166388
rect 295886 166376 295892 166388
rect 209188 166348 295892 166376
rect 209188 166336 209194 166348
rect 295886 166336 295892 166348
rect 295944 166336 295950 166388
rect 369302 166336 369308 166388
rect 369360 166376 369366 166388
rect 485958 166376 485964 166388
rect 369360 166348 485964 166376
rect 369360 166336 369366 166348
rect 485958 166336 485964 166348
rect 486016 166336 486022 166388
rect 42518 166268 42524 166320
rect 42576 166308 42582 166320
rect 165890 166308 165896 166320
rect 42576 166280 165896 166308
rect 42576 166268 42582 166280
rect 165890 166268 165896 166280
rect 165948 166268 165954 166320
rect 202230 166268 202236 166320
rect 202288 166308 202294 166320
rect 303522 166308 303528 166320
rect 202288 166280 303528 166308
rect 202288 166268 202294 166280
rect 303522 166268 303528 166280
rect 303580 166268 303586 166320
rect 366542 166268 366548 166320
rect 366600 166308 366606 166320
rect 483382 166308 483388 166320
rect 366600 166280 483388 166308
rect 366600 166268 366606 166280
rect 483382 166268 483388 166280
rect 483440 166268 483446 166320
rect 50614 166200 50620 166252
rect 50672 166240 50678 166252
rect 96062 166240 96068 166252
rect 50672 166212 96068 166240
rect 50672 166200 50678 166212
rect 96062 166200 96068 166212
rect 96120 166200 96126 166252
rect 517606 165860 517612 165912
rect 517664 165900 517670 165912
rect 517974 165900 517980 165912
rect 517664 165872 517980 165900
rect 517664 165860 517670 165872
rect 517974 165860 517980 165872
rect 518032 165860 518038 165912
rect 53006 165656 53012 165708
rect 53064 165696 53070 165708
rect 114370 165696 114376 165708
rect 53064 165668 114376 165696
rect 53064 165656 53070 165668
rect 114370 165656 114376 165668
rect 114428 165656 114434 165708
rect 54018 165588 54024 165640
rect 54076 165628 54082 165640
rect 54386 165628 54392 165640
rect 54076 165600 54392 165628
rect 54076 165588 54082 165600
rect 54386 165588 54392 165600
rect 54444 165628 54450 165640
rect 116946 165628 116952 165640
rect 54444 165600 116952 165628
rect 54444 165588 54450 165600
rect 116946 165588 116952 165600
rect 117004 165588 117010 165640
rect 357434 165588 357440 165640
rect 357492 165628 357498 165640
rect 360194 165628 360200 165640
rect 357492 165600 360200 165628
rect 357492 165588 357498 165600
rect 360194 165588 360200 165600
rect 360252 165588 360258 165640
rect 375834 165588 375840 165640
rect 375892 165628 375898 165640
rect 436094 165628 436100 165640
rect 375892 165600 436100 165628
rect 375892 165588 375898 165600
rect 436094 165588 436100 165600
rect 436152 165588 436158 165640
rect 56502 165520 56508 165572
rect 56560 165560 56566 165572
rect 132494 165560 132500 165572
rect 56560 165532 132500 165560
rect 56560 165520 56566 165532
rect 132494 165520 132500 165532
rect 132552 165520 132558 165572
rect 214742 165520 214748 165572
rect 214800 165560 214806 165572
rect 300854 165560 300860 165572
rect 214800 165532 300860 165560
rect 214800 165520 214806 165532
rect 300854 165520 300860 165532
rect 300912 165520 300918 165572
rect 362494 165520 362500 165572
rect 362552 165560 362558 165572
rect 455414 165560 455420 165572
rect 362552 165532 455420 165560
rect 362552 165520 362558 165532
rect 455414 165520 455420 165532
rect 455472 165520 455478 165572
rect 517606 165520 517612 165572
rect 517664 165560 517670 165572
rect 517882 165560 517888 165572
rect 517664 165532 517888 165560
rect 517664 165520 517670 165532
rect 517882 165520 517888 165532
rect 517940 165520 517946 165572
rect 55030 165452 55036 165504
rect 55088 165492 55094 165504
rect 129734 165492 129740 165504
rect 55088 165464 129740 165492
rect 55088 165452 55094 165464
rect 129734 165452 129740 165464
rect 129792 165452 129798 165504
rect 214558 165452 214564 165504
rect 214616 165492 214622 165504
rect 280246 165492 280252 165504
rect 214616 165464 280252 165492
rect 214616 165452 214622 165464
rect 280246 165452 280252 165464
rect 280304 165452 280310 165504
rect 369210 165452 369216 165504
rect 369268 165492 369274 165504
rect 458358 165492 458364 165504
rect 369268 165464 458364 165492
rect 369268 165452 369274 165464
rect 458358 165452 458364 165464
rect 458416 165452 458422 165504
rect 56318 165384 56324 165436
rect 56376 165424 56382 165436
rect 128354 165424 128360 165436
rect 56376 165396 128360 165424
rect 56376 165384 56382 165396
rect 128354 165384 128360 165396
rect 128412 165384 128418 165436
rect 211890 165384 211896 165436
rect 211948 165424 211954 165436
rect 277394 165424 277400 165436
rect 211948 165396 277400 165424
rect 211948 165384 211954 165396
rect 277394 165384 277400 165396
rect 277452 165384 277458 165436
rect 360930 165384 360936 165436
rect 360988 165424 360994 165436
rect 442994 165424 443000 165436
rect 360988 165396 443000 165424
rect 360988 165384 360994 165396
rect 442994 165384 443000 165396
rect 443052 165384 443058 165436
rect 55122 165316 55128 165368
rect 55180 165356 55186 165368
rect 125870 165356 125876 165368
rect 55180 165328 125876 165356
rect 55180 165316 55186 165328
rect 125870 165316 125876 165328
rect 125928 165316 125934 165368
rect 218790 165316 218796 165368
rect 218848 165356 218854 165368
rect 283374 165356 283380 165368
rect 218848 165328 283380 165356
rect 218848 165316 218854 165328
rect 283374 165316 283380 165328
rect 283432 165316 283438 165368
rect 370590 165316 370596 165368
rect 370648 165356 370654 165368
rect 452654 165356 452660 165368
rect 370648 165328 452660 165356
rect 370648 165316 370654 165328
rect 452654 165316 452660 165328
rect 452712 165316 452718 165368
rect 53466 165248 53472 165300
rect 53524 165288 53530 165300
rect 120902 165288 120908 165300
rect 53524 165260 120908 165288
rect 53524 165248 53530 165260
rect 120902 165248 120908 165260
rect 120960 165248 120966 165300
rect 207658 165248 207664 165300
rect 207716 165288 207722 165300
rect 267734 165288 267740 165300
rect 207716 165260 267740 165288
rect 207716 165248 207722 165260
rect 267734 165248 267740 165260
rect 267792 165248 267798 165300
rect 371970 165248 371976 165300
rect 372028 165288 372034 165300
rect 449894 165288 449900 165300
rect 372028 165260 449900 165288
rect 372028 165248 372034 165260
rect 449894 165248 449900 165260
rect 449952 165248 449958 165300
rect 56226 165180 56232 165232
rect 56284 165220 56290 165232
rect 123478 165220 123484 165232
rect 56284 165192 123484 165220
rect 56284 165180 56290 165192
rect 123478 165180 123484 165192
rect 123536 165180 123542 165232
rect 183278 165180 183284 165232
rect 183336 165220 183342 165232
rect 197354 165220 197360 165232
rect 183336 165192 197360 165220
rect 183336 165180 183342 165192
rect 197354 165180 197360 165192
rect 197412 165180 197418 165232
rect 216030 165180 216036 165232
rect 216088 165220 216094 165232
rect 273438 165220 273444 165232
rect 216088 165192 273444 165220
rect 216088 165180 216094 165192
rect 273438 165180 273444 165192
rect 273496 165180 273502 165232
rect 373350 165180 373356 165232
rect 373408 165220 373414 165232
rect 447318 165220 447324 165232
rect 373408 165192 447324 165220
rect 373408 165180 373414 165192
rect 447318 165180 447324 165192
rect 447376 165180 447382 165232
rect 54938 165112 54944 165164
rect 54996 165152 55002 165164
rect 118326 165152 118332 165164
rect 54996 165124 118332 165152
rect 54996 165112 55002 165124
rect 118326 165112 118332 165124
rect 118384 165112 118390 165164
rect 218974 165112 218980 165164
rect 219032 165152 219038 165164
rect 276198 165152 276204 165164
rect 219032 165124 276204 165152
rect 219032 165112 219038 165124
rect 276198 165112 276204 165124
rect 276256 165112 276262 165164
rect 370498 165112 370504 165164
rect 370556 165152 370562 165164
rect 438026 165152 438032 165164
rect 370556 165124 438032 165152
rect 370556 165112 370562 165124
rect 438026 165112 438032 165124
rect 438084 165112 438090 165164
rect 53374 165044 53380 165096
rect 53432 165084 53438 165096
rect 113542 165084 113548 165096
rect 53432 165056 113548 165084
rect 53432 165044 53438 165056
rect 113542 165044 113548 165056
rect 113600 165044 113606 165096
rect 183370 165044 183376 165096
rect 183428 165084 183434 165096
rect 197446 165084 197452 165096
rect 183428 165056 197452 165084
rect 183428 165044 183434 165056
rect 197446 165044 197452 165056
rect 197504 165044 197510 165096
rect 215938 165044 215944 165096
rect 215996 165084 216002 165096
rect 258074 165084 258080 165096
rect 215996 165056 258080 165084
rect 215996 165044 216002 165056
rect 258074 165044 258080 165056
rect 258132 165044 258138 165096
rect 367830 165044 367836 165096
rect 367888 165084 367894 165096
rect 419258 165084 419264 165096
rect 367888 165056 419264 165084
rect 367888 165044 367894 165056
rect 419258 165044 419264 165056
rect 419316 165044 419322 165096
rect 503254 165044 503260 165096
rect 503312 165084 503318 165096
rect 517974 165084 517980 165096
rect 503312 165056 517980 165084
rect 503312 165044 503318 165056
rect 517974 165044 517980 165056
rect 518032 165044 518038 165096
rect 56134 164976 56140 165028
rect 56192 165016 56198 165028
rect 115934 165016 115940 165028
rect 56192 164988 115940 165016
rect 56192 164976 56198 164988
rect 115934 164976 115940 164988
rect 115992 164976 115998 165028
rect 211798 164976 211804 165028
rect 211856 165016 211862 165028
rect 252554 165016 252560 165028
rect 211856 164988 252560 165016
rect 211856 164976 211862 164988
rect 252554 164976 252560 164988
rect 252612 164976 252618 165028
rect 343450 164976 343456 165028
rect 343508 165016 343514 165028
rect 356882 165016 356888 165028
rect 343508 164988 356888 165016
rect 343508 164976 343514 164988
rect 356882 164976 356888 164988
rect 356940 164976 356946 165028
rect 374822 164976 374828 165028
rect 374880 165016 374886 165028
rect 440326 165016 440332 165028
rect 374880 164988 440332 165016
rect 374880 164976 374886 164988
rect 440326 164976 440332 164988
rect 440384 164976 440390 165028
rect 52086 164908 52092 164960
rect 52144 164948 52150 164960
rect 103514 164948 103520 164960
rect 52144 164920 103520 164948
rect 52144 164908 52150 164920
rect 103514 164908 103520 164920
rect 103572 164908 103578 164960
rect 114554 164908 114560 164960
rect 114612 164948 114618 164960
rect 196710 164948 196716 164960
rect 114612 164920 196716 164948
rect 114612 164908 114618 164920
rect 196710 164908 196716 164920
rect 196768 164908 196774 164960
rect 210510 164908 210516 164960
rect 210568 164948 210574 164960
rect 249794 164948 249800 164960
rect 210568 164920 249800 164948
rect 210568 164908 210574 164920
rect 249794 164908 249800 164920
rect 249852 164908 249858 164960
rect 369394 164908 369400 164960
rect 369452 164948 369458 164960
rect 434714 164948 434720 164960
rect 369452 164920 434720 164948
rect 369452 164908 369458 164920
rect 434714 164908 434720 164920
rect 434772 164908 434778 164960
rect 503346 164908 503352 164960
rect 503404 164948 503410 164960
rect 503404 164920 509234 164948
rect 503404 164908 503410 164920
rect 50706 164840 50712 164892
rect 50764 164880 50770 164892
rect 89990 164880 89996 164892
rect 50764 164852 89996 164880
rect 50764 164840 50770 164852
rect 89990 164840 89996 164852
rect 90048 164840 90054 164892
rect 113174 164840 113180 164892
rect 113232 164880 113238 164892
rect 196618 164880 196624 164892
rect 113232 164852 196624 164880
rect 113232 164840 113238 164852
rect 196618 164840 196624 164852
rect 196676 164840 196682 164892
rect 218882 164840 218888 164892
rect 218940 164880 218946 164892
rect 247678 164880 247684 164892
rect 218940 164852 247684 164880
rect 218940 164840 218946 164852
rect 247678 164840 247684 164852
rect 247736 164840 247742 164892
rect 343542 164840 343548 164892
rect 343600 164880 343606 164892
rect 357434 164880 357440 164892
rect 343600 164852 357440 164880
rect 343600 164840 343606 164852
rect 357434 164840 357440 164852
rect 357492 164880 357498 164892
rect 357618 164880 357624 164892
rect 357492 164852 357624 164880
rect 357492 164840 357498 164852
rect 357618 164840 357624 164852
rect 357676 164840 357682 164892
rect 363874 164840 363880 164892
rect 363932 164880 363938 164892
rect 409874 164880 409880 164892
rect 363932 164852 409880 164880
rect 363932 164840 363938 164852
rect 409874 164840 409880 164852
rect 409932 164840 409938 164892
rect 419258 164840 419264 164892
rect 419316 164880 419322 164892
rect 433334 164880 433340 164892
rect 419316 164852 433340 164880
rect 419316 164840 419322 164852
rect 433334 164840 433340 164852
rect 433392 164840 433398 164892
rect 509206 164880 509234 164920
rect 510522 164908 510528 164960
rect 510580 164948 510586 164960
rect 517514 164948 517520 164960
rect 510580 164920 517520 164948
rect 510580 164908 510586 164920
rect 517514 164908 517520 164920
rect 517572 164908 517578 164960
rect 517606 164880 517612 164892
rect 509206 164852 517612 164880
rect 517606 164840 517612 164852
rect 517664 164840 517670 164892
rect 52178 164772 52184 164824
rect 52236 164812 52242 164824
rect 88334 164812 88340 164824
rect 52236 164784 88340 164812
rect 52236 164772 52242 164784
rect 88334 164772 88340 164784
rect 88392 164772 88398 164824
rect 115934 164772 115940 164824
rect 115992 164812 115998 164824
rect 197722 164812 197728 164824
rect 115992 164784 197728 164812
rect 115992 164772 115998 164784
rect 197722 164772 197728 164784
rect 197780 164772 197786 164824
rect 366450 164772 366456 164824
rect 366508 164812 366514 164824
rect 407114 164812 407120 164824
rect 366508 164784 407120 164812
rect 366508 164772 366514 164784
rect 407114 164772 407120 164784
rect 407172 164772 407178 164824
rect 428918 164772 428924 164824
rect 428976 164812 428982 164824
rect 433426 164812 433432 164824
rect 428976 164784 433432 164812
rect 428976 164772 428982 164784
rect 433426 164772 433432 164784
rect 433484 164772 433490 164824
rect 374730 164704 374736 164756
rect 374788 164744 374794 164756
rect 412634 164744 412640 164756
rect 374788 164716 412640 164744
rect 374788 164704 374794 164716
rect 412634 164704 412640 164716
rect 412692 164704 412698 164756
rect 378870 164636 378876 164688
rect 378928 164676 378934 164688
rect 416038 164676 416044 164688
rect 378928 164648 416044 164676
rect 378928 164636 378934 164648
rect 416038 164636 416044 164648
rect 416096 164636 416102 164688
rect 98638 164432 98644 164484
rect 98696 164472 98702 164484
rect 100754 164472 100760 164484
rect 98696 164444 100760 164472
rect 98696 164432 98702 164444
rect 100754 164432 100760 164444
rect 100812 164432 100818 164484
rect 83458 164364 83464 164416
rect 83516 164404 83522 164416
rect 107654 164404 107660 164416
rect 83516 164376 107660 164404
rect 83516 164364 83522 164376
rect 107654 164364 107660 164376
rect 107712 164364 107718 164416
rect 87598 164296 87604 164348
rect 87656 164336 87662 164348
rect 106274 164336 106280 164348
rect 87656 164308 106280 164336
rect 87656 164296 87662 164308
rect 106274 164296 106280 164308
rect 106332 164296 106338 164348
rect 49050 164160 49056 164212
rect 49108 164200 49114 164212
rect 50890 164200 50896 164212
rect 49108 164172 50896 164200
rect 49108 164160 49114 164172
rect 50890 164160 50896 164172
rect 50948 164160 50954 164212
rect 58618 164160 58624 164212
rect 58676 164200 58682 164212
rect 59998 164200 60004 164212
rect 58676 164172 60004 164200
rect 58676 164160 58682 164172
rect 59998 164160 60004 164172
rect 60056 164160 60062 164212
rect 117958 164200 117964 164212
rect 62684 164172 117964 164200
rect 46382 164092 46388 164144
rect 46440 164132 46446 164144
rect 50798 164132 50804 164144
rect 46440 164104 50804 164132
rect 46440 164092 46446 164104
rect 50798 164092 50804 164104
rect 50856 164092 50862 164144
rect 58158 164024 58164 164076
rect 58216 164064 58222 164076
rect 62684 164064 62712 164172
rect 117958 164160 117964 164172
rect 118016 164160 118022 164212
rect 211982 164160 211988 164212
rect 212040 164200 212046 164212
rect 323302 164200 323308 164212
rect 212040 164172 323308 164200
rect 212040 164160 212046 164172
rect 323302 164160 323308 164172
rect 323360 164160 323366 164212
rect 361022 164160 361028 164212
rect 361080 164200 361086 164212
rect 430574 164200 430580 164212
rect 361080 164172 430580 164200
rect 361080 164160 361086 164172
rect 430574 164160 430580 164172
rect 430632 164160 430638 164212
rect 110874 164132 110880 164144
rect 58216 164036 62712 164064
rect 64846 164104 110880 164132
rect 58216 164024 58222 164036
rect 56962 163956 56968 164008
rect 57020 163996 57026 164008
rect 59354 163996 59360 164008
rect 57020 163968 59360 163996
rect 57020 163956 57026 163968
rect 59354 163956 59360 163968
rect 59412 163956 59418 164008
rect 53650 163888 53656 163940
rect 53708 163928 53714 163940
rect 64846 163928 64874 164104
rect 110874 164092 110880 164104
rect 110932 164092 110938 164144
rect 219618 164092 219624 164144
rect 219676 164132 219682 164144
rect 264974 164132 264980 164144
rect 219676 164104 264980 164132
rect 219676 164092 219682 164104
rect 264974 164092 264980 164104
rect 265032 164092 265038 164144
rect 374270 164092 374276 164144
rect 374328 164132 374334 164144
rect 374914 164132 374920 164144
rect 374328 164104 374920 164132
rect 374328 164092 374334 164104
rect 374914 164092 374920 164104
rect 374972 164132 374978 164144
rect 434806 164132 434812 164144
rect 374972 164104 434812 164132
rect 374972 164092 374978 164104
rect 434806 164092 434812 164104
rect 434864 164092 434870 164144
rect 213178 164024 213184 164076
rect 213236 164064 213242 164076
rect 235994 164064 236000 164076
rect 213236 164036 236000 164064
rect 213236 164024 213242 164036
rect 235994 164024 236000 164036
rect 236052 164024 236058 164076
rect 374546 164024 374552 164076
rect 374604 164064 374610 164076
rect 431954 164064 431960 164076
rect 374604 164036 431960 164064
rect 374604 164024 374610 164036
rect 431954 164024 431960 164036
rect 432012 164024 432018 164076
rect 216214 163956 216220 164008
rect 216272 163996 216278 164008
rect 236086 163996 236092 164008
rect 216272 163968 236092 163996
rect 216272 163956 216278 163968
rect 236086 163956 236092 163968
rect 236144 163956 236150 164008
rect 379698 163956 379704 164008
rect 379756 163996 379762 164008
rect 426526 163996 426532 164008
rect 379756 163968 426532 163996
rect 379756 163956 379762 163968
rect 426526 163956 426532 163968
rect 426584 163956 426590 164008
rect 53708 163900 64874 163928
rect 53708 163888 53714 163900
rect 375006 163888 375012 163940
rect 375064 163928 375070 163940
rect 396166 163928 396172 163940
rect 375064 163900 396172 163928
rect 375064 163888 375070 163900
rect 396166 163888 396172 163900
rect 396224 163888 396230 163940
rect 51534 163820 51540 163872
rect 51592 163860 51598 163872
rect 56870 163860 56876 163872
rect 51592 163832 56876 163860
rect 51592 163820 51598 163832
rect 56870 163820 56876 163832
rect 56928 163860 56934 163872
rect 95234 163860 95240 163872
rect 56928 163832 95240 163860
rect 56928 163820 56934 163832
rect 95234 163820 95240 163832
rect 95292 163820 95298 163872
rect 375742 163820 375748 163872
rect 375800 163860 375806 163872
rect 396074 163860 396080 163872
rect 375800 163832 396080 163860
rect 375800 163820 375806 163832
rect 396074 163820 396080 163832
rect 396132 163820 396138 163872
rect 52914 163752 52920 163804
rect 52972 163792 52978 163804
rect 56502 163792 56508 163804
rect 52972 163764 56508 163792
rect 52972 163752 52978 163764
rect 56502 163752 56508 163764
rect 56560 163792 56566 163804
rect 96614 163792 96620 163804
rect 56560 163764 96620 163792
rect 56560 163752 56566 163764
rect 96614 163752 96620 163764
rect 96672 163752 96678 163804
rect 59998 163684 60004 163736
rect 60056 163724 60062 163736
rect 106366 163724 106372 163736
rect 60056 163696 106372 163724
rect 60056 163684 60062 163696
rect 106366 163684 106372 163696
rect 106424 163684 106430 163736
rect 50890 163616 50896 163668
rect 50948 163656 50954 163668
rect 109494 163656 109500 163668
rect 50948 163628 109500 163656
rect 50948 163616 50954 163628
rect 109494 163616 109500 163628
rect 109552 163616 109558 163668
rect 59354 163548 59360 163600
rect 59412 163588 59418 163600
rect 118970 163588 118976 163600
rect 59412 163560 118976 163588
rect 59412 163548 59418 163560
rect 118970 163548 118976 163560
rect 119028 163548 119034 163600
rect 373534 163548 373540 163600
rect 373592 163588 373598 163600
rect 375190 163588 375196 163600
rect 373592 163560 375196 163588
rect 373592 163548 373598 163560
rect 375190 163548 375196 163560
rect 375248 163588 375254 163600
rect 429286 163588 429292 163600
rect 375248 163560 429292 163588
rect 375248 163548 375254 163560
rect 429286 163548 429292 163560
rect 429344 163548 429350 163600
rect 50798 163480 50804 163532
rect 50856 163520 50862 163532
rect 111150 163520 111156 163532
rect 50856 163492 111156 163520
rect 50856 163480 50862 163492
rect 111150 163480 111156 163492
rect 111208 163480 111214 163532
rect 216674 163480 216680 163532
rect 216732 163520 216738 163532
rect 218974 163520 218980 163532
rect 216732 163492 218980 163520
rect 216732 163480 216738 163492
rect 218974 163480 218980 163492
rect 219032 163520 219038 163532
rect 263778 163520 263784 163532
rect 219032 163492 263784 163520
rect 219032 163480 219038 163492
rect 263778 163480 263784 163492
rect 263836 163480 263842 163532
rect 373074 163480 373080 163532
rect 373132 163520 373138 163532
rect 375098 163520 375104 163532
rect 373132 163492 375104 163520
rect 373132 163480 373138 163492
rect 375098 163480 375104 163492
rect 375156 163520 375162 163532
rect 430666 163520 430672 163532
rect 375156 163492 430672 163520
rect 375156 163480 375162 163492
rect 430666 163480 430672 163492
rect 430724 163480 430730 163532
rect 57146 162800 57152 162852
rect 57204 162840 57210 162852
rect 59078 162840 59084 162852
rect 57204 162812 59084 162840
rect 57204 162800 57210 162812
rect 59078 162800 59084 162812
rect 59136 162800 59142 162852
rect 214282 162800 214288 162852
rect 214340 162840 214346 162852
rect 214466 162840 214472 162852
rect 214340 162812 214472 162840
rect 214340 162800 214346 162812
rect 214466 162800 214472 162812
rect 214524 162800 214530 162852
rect 214834 162800 214840 162852
rect 214892 162840 214898 162852
rect 260834 162840 260840 162852
rect 214892 162812 260840 162840
rect 214892 162800 214898 162812
rect 260834 162800 260840 162812
rect 260892 162800 260898 162852
rect 376478 162800 376484 162852
rect 376536 162840 376542 162852
rect 379606 162840 379612 162852
rect 376536 162812 379612 162840
rect 376536 162800 376542 162812
rect 379606 162800 379612 162812
rect 379664 162800 379670 162852
rect 379974 162800 379980 162852
rect 380032 162840 380038 162852
rect 428918 162840 428924 162852
rect 380032 162812 428924 162840
rect 380032 162800 380038 162812
rect 428918 162800 428924 162812
rect 428976 162800 428982 162852
rect 214484 162772 214512 162800
rect 259546 162772 259552 162784
rect 214484 162744 259552 162772
rect 259546 162732 259552 162744
rect 259604 162732 259610 162784
rect 376754 162732 376760 162784
rect 376812 162772 376818 162784
rect 420914 162772 420920 162784
rect 376812 162744 420920 162772
rect 376812 162732 376818 162744
rect 420914 162732 420920 162744
rect 420972 162732 420978 162784
rect 217962 162664 217968 162716
rect 218020 162704 218026 162716
rect 259454 162704 259460 162716
rect 218020 162676 259460 162704
rect 218020 162664 218026 162676
rect 259454 162664 259460 162676
rect 259512 162664 259518 162716
rect 376202 162664 376208 162716
rect 376260 162704 376266 162716
rect 418522 162704 418528 162716
rect 376260 162676 418528 162704
rect 376260 162664 376266 162676
rect 418522 162664 418528 162676
rect 418580 162664 418586 162716
rect 218514 162596 218520 162648
rect 218572 162636 218578 162648
rect 218882 162636 218888 162648
rect 218572 162608 218888 162636
rect 218572 162596 218578 162608
rect 218882 162596 218888 162608
rect 218940 162636 218946 162648
rect 258074 162636 258080 162648
rect 218940 162608 258080 162636
rect 218940 162596 218946 162608
rect 258074 162596 258080 162608
rect 258132 162596 258138 162648
rect 375742 162596 375748 162648
rect 375800 162636 375806 162648
rect 378686 162636 378692 162648
rect 375800 162608 378692 162636
rect 375800 162596 375806 162608
rect 378686 162596 378692 162608
rect 378744 162636 378750 162648
rect 419534 162636 419540 162648
rect 378744 162608 419540 162636
rect 378744 162596 378750 162608
rect 419534 162596 419540 162608
rect 419592 162596 419598 162648
rect 375282 162528 375288 162580
rect 375340 162568 375346 162580
rect 379974 162568 379980 162580
rect 375340 162540 379980 162568
rect 375340 162528 375346 162540
rect 379974 162528 379980 162540
rect 380032 162528 380038 162580
rect 374362 162460 374368 162512
rect 374420 162500 374426 162512
rect 378962 162500 378968 162512
rect 374420 162472 378968 162500
rect 374420 162460 374426 162472
rect 378962 162460 378968 162472
rect 379020 162460 379026 162512
rect 59078 162120 59084 162172
rect 59136 162160 59142 162172
rect 89898 162160 89904 162172
rect 59136 162132 89904 162160
rect 59136 162120 59142 162132
rect 89898 162120 89904 162132
rect 89956 162120 89962 162172
rect 218606 162120 218612 162172
rect 218664 162160 218670 162172
rect 219526 162160 219532 162172
rect 218664 162132 219532 162160
rect 218664 162120 218670 162132
rect 219526 162120 219532 162132
rect 219584 162160 219590 162172
rect 266354 162160 266360 162172
rect 219584 162132 266360 162160
rect 219584 162120 219590 162132
rect 266354 162120 266360 162132
rect 266412 162120 266418 162172
rect 379606 162120 379612 162172
rect 379664 162160 379670 162172
rect 418154 162160 418160 162172
rect 379664 162132 418160 162160
rect 379664 162120 379670 162132
rect 418154 162120 418160 162132
rect 418212 162120 418218 162172
rect 376294 161848 376300 161900
rect 376352 161888 376358 161900
rect 376754 161888 376760 161900
rect 376352 161860 376760 161888
rect 376352 161848 376358 161860
rect 376754 161848 376760 161860
rect 376812 161848 376818 161900
rect 216122 161576 216128 161628
rect 216180 161616 216186 161628
rect 216180 161588 219434 161616
rect 216180 161576 216186 161588
rect 219406 161548 219434 161588
rect 235258 161548 235264 161560
rect 219406 161520 235264 161548
rect 235258 161508 235264 161520
rect 235316 161508 235322 161560
rect 217134 161440 217140 161492
rect 217192 161480 217198 161492
rect 236638 161480 236644 161492
rect 217192 161452 236644 161480
rect 217192 161440 217198 161452
rect 236638 161440 236644 161452
rect 236696 161440 236702 161492
rect 378962 161440 378968 161492
rect 379020 161480 379026 161492
rect 396718 161480 396724 161492
rect 379020 161452 396724 161480
rect 379020 161440 379026 161452
rect 396718 161440 396724 161452
rect 396776 161440 396782 161492
rect 58066 148996 58072 149048
rect 58124 149036 58130 149048
rect 106274 149036 106280 149048
rect 58124 149008 106280 149036
rect 58124 148996 58130 149008
rect 106274 148996 106280 149008
rect 106332 148996 106338 149048
rect 213270 148996 213276 149048
rect 213328 149036 213334 149048
rect 276106 149036 276112 149048
rect 213328 149008 276112 149036
rect 213328 148996 213334 149008
rect 276106 148996 276112 149008
rect 276164 148996 276170 149048
rect 379054 148996 379060 149048
rect 379112 149036 379118 149048
rect 440234 149036 440240 149048
rect 379112 149008 440240 149036
rect 379112 148996 379118 149008
rect 440234 148996 440240 149008
rect 440292 148996 440298 149048
rect 58710 148928 58716 148980
rect 58768 148968 58774 148980
rect 103514 148968 103520 148980
rect 58768 148940 103520 148968
rect 58768 148928 58774 148940
rect 103514 148928 103520 148940
rect 103572 148928 103578 148980
rect 213454 148928 213460 148980
rect 213512 148968 213518 148980
rect 274726 148968 274732 148980
rect 213512 148940 274732 148968
rect 213512 148928 213518 148940
rect 274726 148928 274732 148940
rect 274784 148928 274790 148980
rect 373810 148928 373816 148980
rect 373868 148968 373874 148980
rect 434714 148968 434720 148980
rect 373868 148940 434720 148968
rect 373868 148928 373874 148940
rect 434714 148928 434720 148940
rect 434772 148928 434778 148980
rect 216306 148860 216312 148912
rect 216364 148900 216370 148912
rect 277394 148900 277400 148912
rect 216364 148872 277400 148900
rect 216364 148860 216370 148872
rect 277394 148860 277400 148872
rect 277452 148860 277458 148912
rect 379790 148860 379796 148912
rect 379848 148900 379854 148912
rect 427814 148900 427820 148912
rect 379848 148872 427820 148900
rect 379848 148860 379854 148872
rect 427814 148860 427820 148872
rect 427872 148860 427878 148912
rect 46658 148792 46664 148844
rect 46716 148832 46722 148844
rect 59906 148832 59912 148844
rect 46716 148804 59912 148832
rect 46716 148792 46722 148804
rect 59906 148792 59912 148804
rect 59964 148832 59970 148844
rect 83458 148832 83464 148844
rect 59964 148804 83464 148832
rect 59964 148792 59970 148804
rect 83458 148792 83464 148804
rect 83516 148792 83522 148844
rect 214926 148792 214932 148844
rect 214984 148832 214990 148844
rect 274634 148832 274640 148844
rect 214984 148804 274640 148832
rect 214984 148792 214990 148804
rect 274634 148792 274640 148804
rect 274692 148792 274698 148844
rect 373718 148792 373724 148844
rect 373776 148832 373782 148844
rect 397454 148832 397460 148844
rect 373776 148804 397460 148832
rect 373776 148792 373782 148804
rect 397454 148792 397460 148804
rect 397512 148792 397518 148844
rect 48038 148724 48044 148776
rect 48096 148764 48102 148776
rect 55030 148764 55036 148776
rect 48096 148736 55036 148764
rect 48096 148724 48102 148736
rect 55030 148724 55036 148736
rect 55088 148764 55094 148776
rect 80054 148764 80060 148776
rect 55088 148736 80060 148764
rect 55088 148724 55094 148736
rect 80054 148724 80060 148736
rect 80112 148724 80118 148776
rect 213546 148724 213552 148776
rect 213604 148764 213610 148776
rect 241514 148764 241520 148776
rect 213604 148736 241520 148764
rect 213604 148724 213610 148736
rect 241514 148724 241520 148736
rect 241572 148724 241578 148776
rect 46474 148656 46480 148708
rect 46532 148696 46538 148708
rect 58986 148696 58992 148708
rect 46532 148668 58992 148696
rect 46532 148656 46538 148668
rect 58986 148656 58992 148668
rect 59044 148696 59050 148708
rect 87598 148696 87604 148708
rect 59044 148668 87604 148696
rect 59044 148656 59050 148668
rect 87598 148656 87604 148668
rect 87656 148656 87662 148708
rect 49142 148588 49148 148640
rect 49200 148628 49206 148640
rect 52178 148628 52184 148640
rect 49200 148600 52184 148628
rect 49200 148588 49206 148600
rect 52178 148588 52184 148600
rect 52236 148628 52242 148640
rect 81434 148628 81440 148640
rect 52236 148600 81440 148628
rect 52236 148588 52242 148600
rect 81434 148588 81440 148600
rect 81492 148588 81498 148640
rect 54478 148520 54484 148572
rect 54536 148560 54542 148572
rect 56226 148560 56232 148572
rect 54536 148532 56232 148560
rect 54536 148520 54542 148532
rect 56226 148520 56232 148532
rect 56284 148560 56290 148572
rect 102134 148560 102140 148572
rect 56284 148532 102140 148560
rect 56284 148520 56290 148532
rect 102134 148520 102140 148532
rect 102192 148520 102198 148572
rect 213730 148520 213736 148572
rect 213788 148560 213794 148572
rect 238754 148560 238760 148572
rect 213788 148532 238760 148560
rect 213788 148520 213794 148532
rect 238754 148520 238760 148532
rect 238812 148520 238818 148572
rect 372246 148520 372252 148572
rect 372304 148560 372310 148572
rect 374730 148560 374736 148572
rect 372304 148532 374736 148560
rect 372304 148520 372310 148532
rect 374730 148520 374736 148532
rect 374788 148560 374794 148572
rect 400214 148560 400220 148572
rect 374788 148532 400220 148560
rect 374788 148520 374794 148532
rect 400214 148520 400220 148532
rect 400272 148520 400278 148572
rect 53466 148452 53472 148504
rect 53524 148492 53530 148504
rect 113174 148492 113180 148504
rect 53524 148464 113180 148492
rect 53524 148452 53530 148464
rect 113174 148452 113180 148464
rect 113232 148452 113238 148504
rect 215018 148452 215024 148504
rect 215076 148492 215082 148504
rect 240134 148492 240140 148504
rect 215076 148464 240140 148492
rect 215076 148452 215082 148464
rect 240134 148452 240140 148464
rect 240192 148452 240198 148504
rect 370774 148452 370780 148504
rect 370832 148492 370838 148504
rect 373258 148492 373264 148504
rect 370832 148464 373264 148492
rect 370832 148452 370838 148464
rect 373258 148452 373264 148464
rect 373316 148492 373322 148504
rect 398834 148492 398840 148504
rect 373316 148464 398840 148492
rect 373316 148452 373322 148464
rect 398834 148452 398840 148464
rect 398892 148452 398898 148504
rect 53558 148384 53564 148436
rect 53616 148424 53622 148436
rect 114554 148424 114560 148436
rect 53616 148396 114560 148424
rect 53616 148384 53622 148396
rect 114554 148384 114560 148396
rect 114612 148384 114618 148436
rect 212166 148384 212172 148436
rect 212224 148424 212230 148436
rect 214650 148424 214656 148436
rect 212224 148396 214656 148424
rect 212224 148384 212230 148396
rect 214650 148384 214656 148396
rect 214708 148424 214714 148436
rect 270494 148424 270500 148436
rect 214708 148396 270500 148424
rect 214708 148384 214714 148396
rect 270494 148384 270500 148396
rect 270552 148384 270558 148436
rect 370958 148384 370964 148436
rect 371016 148424 371022 148436
rect 373350 148424 373356 148436
rect 371016 148396 373356 148424
rect 371016 148384 371022 148396
rect 373350 148384 373356 148396
rect 373408 148424 373414 148436
rect 401594 148424 401600 148436
rect 373408 148396 401600 148424
rect 373408 148384 373414 148396
rect 401594 148384 401600 148396
rect 401652 148384 401658 148436
rect 53374 148316 53380 148368
rect 53432 148356 53438 148368
rect 115934 148356 115940 148368
rect 53432 148328 115940 148356
rect 53432 148316 53438 148328
rect 115934 148316 115940 148328
rect 115992 148316 115998 148368
rect 215754 148316 215760 148368
rect 215812 148356 215818 148368
rect 271874 148356 271880 148368
rect 215812 148328 271880 148356
rect 215812 148316 215818 148328
rect 271874 148316 271880 148328
rect 271932 148316 271938 148368
rect 372522 148316 372528 148368
rect 372580 148356 372586 148368
rect 379974 148356 379980 148368
rect 372580 148328 379980 148356
rect 372580 148316 372586 148328
rect 379974 148316 379980 148328
rect 380032 148356 380038 148368
rect 429194 148356 429200 148368
rect 380032 148328 429200 148356
rect 380032 148316 380038 148328
rect 429194 148316 429200 148328
rect 429252 148316 429258 148368
rect 56318 147636 56324 147688
rect 56376 147676 56382 147688
rect 58710 147676 58716 147688
rect 56376 147648 58716 147676
rect 56376 147636 56382 147648
rect 58710 147636 58716 147648
rect 58768 147636 58774 147688
rect 213362 147636 213368 147688
rect 213420 147676 213426 147688
rect 214926 147676 214932 147688
rect 213420 147648 214932 147676
rect 213420 147636 213426 147648
rect 214926 147636 214932 147648
rect 214984 147636 214990 147688
rect 379330 147636 379336 147688
rect 379388 147676 379394 147688
rect 379790 147676 379796 147688
rect 379388 147648 379796 147676
rect 379388 147636 379394 147648
rect 379790 147636 379796 147648
rect 379848 147636 379854 147688
rect 206738 147568 206744 147620
rect 206796 147608 206802 147620
rect 213178 147608 213184 147620
rect 206796 147580 213184 147608
rect 206796 147568 206802 147580
rect 213178 147568 213184 147580
rect 213236 147608 213242 147620
rect 213730 147608 213736 147620
rect 213236 147580 213736 147608
rect 213236 147568 213242 147580
rect 213730 147568 213736 147580
rect 213788 147568 213794 147620
rect 212258 147500 212264 147552
rect 212316 147540 212322 147552
rect 215754 147540 215760 147552
rect 212316 147512 215760 147540
rect 212316 147500 212322 147512
rect 215754 147500 215760 147512
rect 215812 147540 215818 147552
rect 215938 147540 215944 147552
rect 215812 147512 215944 147540
rect 215812 147500 215818 147512
rect 215938 147500 215944 147512
rect 215996 147500 216002 147552
rect 213270 147432 213276 147484
rect 213328 147472 213334 147484
rect 213730 147472 213736 147484
rect 213328 147444 213736 147472
rect 213328 147432 213334 147444
rect 213730 147432 213736 147444
rect 213788 147432 213794 147484
rect 210970 147364 210976 147416
rect 211028 147404 211034 147416
rect 214558 147404 214564 147416
rect 211028 147376 214564 147404
rect 211028 147364 211034 147376
rect 214558 147364 214564 147376
rect 214616 147404 214622 147416
rect 215018 147404 215024 147416
rect 214616 147376 215024 147404
rect 214616 147364 214622 147376
rect 215018 147364 215024 147376
rect 215076 147364 215082 147416
rect 215018 146276 215024 146328
rect 215076 146316 215082 146328
rect 276014 146316 276020 146328
rect 215076 146288 276020 146316
rect 215076 146276 215082 146288
rect 276014 146276 276020 146288
rect 276072 146316 276078 146328
rect 276072 146288 277394 146316
rect 276072 146276 276078 146288
rect 46290 146208 46296 146260
rect 46348 146248 46354 146260
rect 52086 146248 52092 146260
rect 46348 146220 52092 146248
rect 46348 146208 46354 146220
rect 52086 146208 52092 146220
rect 52144 146208 52150 146260
rect 57054 146208 57060 146260
rect 57112 146248 57118 146260
rect 57974 146248 57980 146260
rect 57112 146220 57980 146248
rect 57112 146208 57118 146220
rect 57974 146208 57980 146220
rect 58032 146208 58038 146260
rect 59814 146208 59820 146260
rect 59872 146248 59878 146260
rect 93854 146248 93860 146260
rect 59872 146220 93860 146248
rect 59872 146208 59878 146220
rect 93854 146208 93860 146220
rect 93912 146208 93918 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197630 146248 197636 146260
rect 179104 146220 197636 146248
rect 179104 146208 179110 146220
rect 197630 146208 197636 146220
rect 197688 146208 197694 146260
rect 236638 146208 236644 146260
rect 236696 146248 236702 146260
rect 256694 146248 256700 146260
rect 236696 146220 256700 146248
rect 236696 146208 236702 146220
rect 256694 146208 256700 146220
rect 256752 146208 256758 146260
rect 277366 146248 277394 146288
rect 356606 146248 356612 146260
rect 277366 146220 356612 146248
rect 356606 146208 356612 146220
rect 356664 146208 356670 146260
rect 375926 146208 375932 146260
rect 375984 146248 375990 146260
rect 377950 146248 377956 146260
rect 375984 146220 377956 146248
rect 375984 146208 375990 146220
rect 377950 146208 377956 146220
rect 378008 146208 378014 146260
rect 378594 146208 378600 146260
rect 378652 146248 378658 146260
rect 379238 146248 379244 146260
rect 378652 146220 379244 146248
rect 378652 146208 378658 146220
rect 379238 146208 379244 146220
rect 379296 146208 379302 146260
rect 379882 146208 379888 146260
rect 379940 146248 379946 146260
rect 414014 146248 414020 146260
rect 379940 146220 414020 146248
rect 379940 146208 379946 146220
rect 414014 146208 414020 146220
rect 414072 146208 414078 146260
rect 57992 146180 58020 146208
rect 91186 146180 91192 146192
rect 57992 146152 91192 146180
rect 91186 146140 91192 146152
rect 91244 146140 91250 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197538 146180 197544 146192
rect 179748 146152 197544 146180
rect 179748 146140 179754 146152
rect 197538 146140 197544 146152
rect 197596 146140 197602 146192
rect 235258 146140 235264 146192
rect 235316 146180 235322 146192
rect 255314 146180 255320 146192
rect 235316 146152 255320 146180
rect 235316 146140 235322 146152
rect 255314 146140 255320 146152
rect 255372 146140 255378 146192
rect 338482 146140 338488 146192
rect 338540 146180 338546 146192
rect 357802 146180 357808 146192
rect 338540 146152 357808 146180
rect 338540 146140 338546 146152
rect 357802 146140 357808 146152
rect 357860 146140 357866 146192
rect 378410 146140 378416 146192
rect 378468 146180 378474 146192
rect 379422 146180 379428 146192
rect 378468 146152 379428 146180
rect 378468 146140 378474 146152
rect 379422 146140 379428 146152
rect 379480 146140 379486 146192
rect 396718 146140 396724 146192
rect 396776 146180 396782 146192
rect 416774 146180 416780 146192
rect 396776 146152 416780 146180
rect 396776 146140 396782 146152
rect 416774 146140 416780 146152
rect 416832 146140 416838 146192
rect 500218 146140 500224 146192
rect 500276 146180 500282 146192
rect 517698 146180 517704 146192
rect 500276 146152 517704 146180
rect 500276 146140 500282 146152
rect 517698 146140 517704 146152
rect 517756 146140 517762 146192
rect 55950 146072 55956 146124
rect 56008 146112 56014 146124
rect 88426 146112 88432 146124
rect 56008 146084 88432 146112
rect 56008 146072 56014 146084
rect 88426 146072 88432 146084
rect 88484 146072 88490 146124
rect 215846 146072 215852 146124
rect 215904 146072 215910 146124
rect 219342 146072 219348 146124
rect 219400 146112 219406 146124
rect 252554 146112 252560 146124
rect 219400 146084 252560 146112
rect 219400 146072 219406 146084
rect 252554 146072 252560 146084
rect 252612 146072 252618 146124
rect 340230 146072 340236 146124
rect 340288 146112 340294 146124
rect 357710 146112 357716 146124
rect 340288 146084 357716 146112
rect 340288 146072 340294 146084
rect 357710 146072 357716 146084
rect 357768 146072 357774 146124
rect 379054 146072 379060 146124
rect 379112 146112 379118 146124
rect 379514 146112 379520 146124
rect 379112 146084 379520 146112
rect 379112 146072 379118 146084
rect 379514 146072 379520 146084
rect 379572 146112 379578 146124
rect 412726 146112 412732 146124
rect 379572 146084 412732 146112
rect 379572 146072 379578 146084
rect 412726 146072 412732 146084
rect 412784 146072 412790 146124
rect 498654 146072 498660 146124
rect 498712 146112 498718 146124
rect 517514 146112 517520 146124
rect 498712 146084 517520 146112
rect 498712 146072 498718 146084
rect 517514 146072 517520 146084
rect 517572 146112 517578 146124
rect 517790 146112 517796 146124
rect 517572 146084 517796 146112
rect 517572 146072 517578 146084
rect 517790 146072 517796 146084
rect 517848 146072 517854 146124
rect 53650 146004 53656 146056
rect 53708 146044 53714 146056
rect 54110 146044 54116 146056
rect 53708 146016 54116 146044
rect 53708 146004 53714 146016
rect 54110 146004 54116 146016
rect 54168 146044 54174 146056
rect 86954 146044 86960 146056
rect 54168 146016 86960 146044
rect 54168 146004 54174 146016
rect 86954 146004 86960 146016
rect 87012 146004 87018 146056
rect 215864 146044 215892 146072
rect 216490 146044 216496 146056
rect 215864 146016 216496 146044
rect 216490 146004 216496 146016
rect 216548 146044 216554 146056
rect 249794 146044 249800 146056
rect 216548 146016 249800 146044
rect 216548 146004 216554 146016
rect 249794 146004 249800 146016
rect 249852 146004 249858 146056
rect 379422 146004 379428 146056
rect 379480 146044 379486 146056
rect 411346 146044 411352 146056
rect 379480 146016 411352 146044
rect 379480 146004 379486 146016
rect 411346 146004 411352 146016
rect 411404 146004 411410 146056
rect 54294 145936 54300 145988
rect 54352 145976 54358 145988
rect 54846 145976 54852 145988
rect 54352 145948 54852 145976
rect 54352 145936 54358 145948
rect 54846 145936 54852 145948
rect 54904 145976 54910 145988
rect 82814 145976 82820 145988
rect 54904 145948 82820 145976
rect 54904 145936 54910 145948
rect 82814 145936 82820 145948
rect 82872 145936 82878 145988
rect 219158 145936 219164 145988
rect 219216 145976 219222 145988
rect 251174 145976 251180 145988
rect 219216 145948 251180 145976
rect 219216 145936 219222 145948
rect 251174 145936 251180 145948
rect 251232 145936 251238 145988
rect 377306 145936 377312 145988
rect 377364 145976 377370 145988
rect 379146 145976 379152 145988
rect 377364 145948 379152 145976
rect 377364 145936 377370 145948
rect 379146 145936 379152 145948
rect 379204 145976 379210 145988
rect 409874 145976 409880 145988
rect 379204 145948 409880 145976
rect 379204 145936 379210 145948
rect 409874 145936 409880 145948
rect 409932 145936 409938 145988
rect 58802 145868 58808 145920
rect 58860 145908 58866 145920
rect 84194 145908 84200 145920
rect 58860 145880 84200 145908
rect 58860 145868 58866 145880
rect 84194 145868 84200 145880
rect 84252 145868 84258 145920
rect 216122 145868 216128 145920
rect 216180 145908 216186 145920
rect 217318 145908 217324 145920
rect 216180 145880 217324 145908
rect 216180 145868 216186 145880
rect 217318 145868 217324 145880
rect 217376 145908 217382 145920
rect 247034 145908 247040 145920
rect 217376 145880 247040 145908
rect 217376 145868 217382 145880
rect 247034 145868 247040 145880
rect 247092 145868 247098 145920
rect 377950 145868 377956 145920
rect 378008 145908 378014 145920
rect 408494 145908 408500 145920
rect 378008 145880 408500 145908
rect 378008 145868 378014 145880
rect 408494 145868 408500 145880
rect 408552 145868 408558 145920
rect 47854 145800 47860 145852
rect 47912 145840 47918 145852
rect 53098 145840 53104 145852
rect 47912 145812 53104 145840
rect 47912 145800 47918 145812
rect 53098 145800 53104 145812
rect 53156 145840 53162 145852
rect 78674 145840 78680 145852
rect 53156 145812 78680 145840
rect 53156 145800 53162 145812
rect 78674 145800 78680 145812
rect 78732 145800 78738 145852
rect 216398 145800 216404 145852
rect 216456 145840 216462 145852
rect 242894 145840 242900 145852
rect 216456 145812 242900 145840
rect 216456 145800 216462 145812
rect 242894 145800 242900 145812
rect 242952 145800 242958 145852
rect 375834 145800 375840 145852
rect 375892 145840 375898 145852
rect 376570 145840 376576 145852
rect 375892 145812 376576 145840
rect 375892 145800 375898 145812
rect 376570 145800 376576 145812
rect 376628 145800 376634 145852
rect 376662 145800 376668 145852
rect 376720 145840 376726 145852
rect 404354 145840 404360 145852
rect 376720 145812 404360 145840
rect 376720 145800 376726 145812
rect 404354 145800 404360 145812
rect 404412 145800 404418 145852
rect 56410 145732 56416 145784
rect 56468 145772 56474 145784
rect 84286 145772 84292 145784
rect 56468 145744 84292 145772
rect 56468 145732 56474 145744
rect 84286 145732 84292 145744
rect 84344 145732 84350 145784
rect 214926 145732 214932 145784
rect 214984 145772 214990 145784
rect 219066 145772 219072 145784
rect 214984 145744 219072 145772
rect 214984 145732 214990 145744
rect 219066 145732 219072 145744
rect 219124 145772 219130 145784
rect 244366 145772 244372 145784
rect 219124 145744 244372 145772
rect 219124 145732 219130 145744
rect 244366 145732 244372 145744
rect 244424 145732 244430 145784
rect 376588 145772 376616 145800
rect 403066 145772 403072 145784
rect 376588 145744 403072 145772
rect 403066 145732 403072 145744
rect 403124 145732 403130 145784
rect 53834 145664 53840 145716
rect 53892 145704 53898 145716
rect 85574 145704 85580 145716
rect 53892 145676 85580 145704
rect 53892 145664 53898 145676
rect 85574 145664 85580 145676
rect 85632 145664 85638 145716
rect 218054 145664 218060 145716
rect 218112 145704 218118 145716
rect 245654 145704 245660 145716
rect 218112 145676 245660 145704
rect 218112 145664 218118 145676
rect 245654 145664 245660 145676
rect 245712 145664 245718 145716
rect 375006 145664 375012 145716
rect 375064 145704 375070 145716
rect 402974 145704 402980 145716
rect 375064 145676 402980 145704
rect 375064 145664 375070 145676
rect 402974 145664 402980 145676
rect 403032 145664 403038 145716
rect 58618 145596 58624 145648
rect 58676 145636 58682 145648
rect 91094 145636 91100 145648
rect 58676 145608 91100 145636
rect 58676 145596 58682 145608
rect 91094 145596 91100 145608
rect 91152 145596 91158 145648
rect 216030 145596 216036 145648
rect 216088 145636 216094 145648
rect 244274 145636 244280 145648
rect 216088 145608 244280 145636
rect 216088 145596 216094 145608
rect 244274 145596 244280 145608
rect 244332 145596 244338 145648
rect 280062 145596 280068 145648
rect 280120 145636 280126 145648
rect 356606 145636 356612 145648
rect 280120 145608 356612 145636
rect 280120 145596 280126 145608
rect 356606 145596 356612 145608
rect 356664 145636 356670 145648
rect 357526 145636 357532 145648
rect 356664 145608 357532 145636
rect 356664 145596 356670 145608
rect 357526 145596 357532 145608
rect 357584 145596 357590 145648
rect 376110 145596 376116 145648
rect 376168 145636 376174 145648
rect 407206 145636 407212 145648
rect 376168 145608 407212 145636
rect 376168 145596 376174 145608
rect 407206 145596 407212 145608
rect 407264 145596 407270 145648
rect 517514 145596 517520 145648
rect 517572 145636 517578 145648
rect 580350 145636 580356 145648
rect 517572 145608 580356 145636
rect 517572 145596 517578 145608
rect 580350 145596 580356 145608
rect 580408 145596 580414 145648
rect 53926 145528 53932 145580
rect 53984 145568 53990 145580
rect 97994 145568 98000 145580
rect 53984 145540 98000 145568
rect 53984 145528 53990 145540
rect 97994 145528 98000 145540
rect 98052 145528 98058 145580
rect 191282 145528 191288 145580
rect 191340 145568 191346 145580
rect 202138 145568 202144 145580
rect 191340 145540 202144 145568
rect 191340 145528 191346 145540
rect 202138 145528 202144 145540
rect 202196 145568 202202 145580
rect 204898 145568 204904 145580
rect 202196 145540 204904 145568
rect 202196 145528 202202 145540
rect 204898 145528 204904 145540
rect 204956 145528 204962 145580
rect 217042 145528 217048 145580
rect 217100 145568 217106 145580
rect 248414 145568 248420 145580
rect 217100 145540 248420 145568
rect 217100 145528 217106 145540
rect 248414 145528 248420 145540
rect 248472 145528 248478 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358078 145568 358084 145580
rect 351696 145540 358084 145568
rect 351696 145528 351702 145540
rect 358078 145528 358084 145540
rect 358136 145568 358142 145580
rect 358722 145568 358728 145580
rect 358136 145540 358728 145568
rect 358136 145528 358142 145540
rect 358722 145528 358728 145540
rect 358780 145568 358786 145580
rect 510522 145568 510528 145580
rect 358780 145540 510528 145568
rect 358780 145528 358786 145540
rect 510522 145528 510528 145540
rect 510580 145528 510586 145580
rect 517698 145528 517704 145580
rect 517756 145568 517762 145580
rect 580258 145568 580264 145580
rect 517756 145540 580264 145568
rect 517756 145528 517762 145540
rect 580258 145528 580264 145540
rect 580316 145528 580322 145580
rect 52086 145460 52092 145512
rect 52144 145500 52150 145512
rect 77294 145500 77300 145512
rect 52144 145472 77300 145500
rect 52144 145460 52150 145472
rect 77294 145460 77300 145472
rect 77352 145460 77358 145512
rect 218514 145460 218520 145512
rect 218572 145500 218578 145512
rect 236086 145500 236092 145512
rect 218572 145472 236092 145500
rect 218572 145460 218578 145472
rect 236086 145460 236092 145472
rect 236144 145460 236150 145512
rect 379238 145460 379244 145512
rect 379296 145500 379302 145512
rect 405734 145500 405740 145512
rect 379296 145472 405740 145500
rect 379296 145460 379302 145472
rect 405734 145460 405740 145472
rect 405792 145460 405798 145512
rect 47946 145392 47952 145444
rect 48004 145432 48010 145444
rect 54386 145432 54392 145444
rect 48004 145404 54392 145432
rect 48004 145392 48010 145404
rect 54386 145392 54392 145404
rect 54444 145432 54450 145444
rect 76006 145432 76012 145444
rect 54444 145404 76012 145432
rect 54444 145392 54450 145404
rect 76006 145392 76012 145404
rect 76064 145392 76070 145444
rect 218606 145392 218612 145444
rect 218664 145432 218670 145444
rect 235994 145432 236000 145444
rect 218664 145404 236000 145432
rect 218664 145392 218670 145404
rect 235994 145392 236000 145404
rect 236052 145392 236058 145444
rect 378686 145392 378692 145444
rect 378744 145432 378750 145444
rect 396166 145432 396172 145444
rect 378744 145404 396172 145432
rect 378744 145392 378750 145404
rect 396166 145392 396172 145404
rect 396224 145392 396230 145444
rect 46566 145324 46572 145376
rect 46624 145364 46630 145376
rect 54938 145364 54944 145376
rect 46624 145336 54944 145364
rect 46624 145324 46630 145336
rect 54938 145324 54944 145336
rect 54996 145364 55002 145376
rect 75914 145364 75920 145376
rect 54996 145336 75920 145364
rect 54996 145324 55002 145336
rect 75914 145324 75920 145336
rect 75972 145324 75978 145376
rect 219802 145324 219808 145376
rect 219860 145364 219866 145376
rect 253934 145364 253940 145376
rect 219860 145336 253940 145364
rect 219860 145324 219866 145336
rect 253934 145324 253940 145336
rect 253992 145324 253998 145376
rect 378778 145324 378784 145376
rect 378836 145364 378842 145376
rect 396074 145364 396080 145376
rect 378836 145336 396080 145364
rect 378836 145324 378842 145336
rect 396074 145324 396080 145336
rect 396132 145324 396138 145376
rect 216766 145256 216772 145308
rect 216824 145296 216830 145308
rect 217226 145296 217232 145308
rect 216824 145268 217232 145296
rect 216824 145256 216830 145268
rect 217226 145256 217232 145268
rect 217284 145296 217290 145308
rect 251266 145296 251272 145308
rect 217284 145268 251272 145296
rect 217284 145256 217290 145268
rect 251266 145256 251272 145268
rect 251324 145256 251330 145308
rect 378042 145256 378048 145308
rect 378100 145296 378106 145308
rect 411254 145296 411260 145308
rect 378100 145268 411260 145296
rect 378100 145256 378106 145268
rect 411254 145256 411260 145268
rect 411312 145256 411318 145308
rect 51718 144848 51724 144900
rect 51776 144888 51782 144900
rect 53834 144888 53840 144900
rect 51776 144860 53840 144888
rect 51776 144848 51782 144860
rect 53834 144848 53840 144860
rect 53892 144888 53898 144900
rect 54478 144888 54484 144900
rect 53892 144860 54484 144888
rect 53892 144848 53898 144860
rect 54478 144848 54484 144860
rect 54536 144848 54542 144900
rect 54570 144848 54576 144900
rect 54628 144888 54634 144900
rect 58802 144888 58808 144900
rect 54628 144860 58808 144888
rect 54628 144848 54634 144860
rect 58802 144848 58808 144860
rect 58860 144848 58866 144900
rect 209498 144848 209504 144900
rect 209556 144888 209562 144900
rect 213270 144888 213276 144900
rect 209556 144860 213276 144888
rect 209556 144848 209562 144860
rect 213270 144848 213276 144860
rect 213328 144848 213334 144900
rect 214374 144848 214380 144900
rect 214432 144888 214438 144900
rect 217042 144888 217048 144900
rect 214432 144860 217048 144888
rect 214432 144848 214438 144860
rect 217042 144848 217048 144860
rect 217100 144848 217106 144900
rect 373626 144848 373632 144900
rect 373684 144888 373690 144900
rect 374822 144888 374828 144900
rect 373684 144860 374828 144888
rect 373684 144848 373690 144860
rect 374822 144848 374828 144860
rect 374880 144888 374886 144900
rect 375006 144888 375012 144900
rect 374880 144860 375012 144888
rect 374880 144848 374886 144860
rect 375006 144848 375012 144860
rect 375064 144848 375070 144900
rect 51810 144780 51816 144832
rect 51868 144820 51874 144832
rect 58618 144820 58624 144832
rect 51868 144792 58624 144820
rect 51868 144780 51874 144792
rect 58618 144780 58624 144792
rect 58676 144780 58682 144832
rect 213638 144780 213644 144832
rect 213696 144820 213702 144832
rect 214466 144820 214472 144832
rect 213696 144792 214472 144820
rect 213696 144780 213702 144792
rect 214466 144780 214472 144792
rect 214524 144780 214530 144832
rect 374454 144780 374460 144832
rect 374512 144820 374518 144832
rect 376110 144820 376116 144832
rect 374512 144792 376116 144820
rect 374512 144780 374518 144792
rect 376110 144780 376116 144792
rect 376168 144780 376174 144832
rect 50430 144712 50436 144764
rect 50488 144752 50494 144764
rect 53926 144752 53932 144764
rect 50488 144724 53932 144752
rect 50488 144712 50494 144724
rect 53926 144712 53932 144724
rect 53984 144752 53990 144764
rect 54662 144752 54668 144764
rect 53984 144724 54668 144752
rect 53984 144712 53990 144724
rect 54662 144712 54668 144724
rect 54720 144712 54726 144764
rect 213086 144712 213092 144764
rect 213144 144752 213150 144764
rect 216030 144752 216036 144764
rect 213144 144724 216036 144752
rect 213144 144712 213150 144724
rect 216030 144712 216036 144724
rect 216088 144712 216094 144764
rect 50522 144644 50528 144696
rect 50580 144684 50586 144696
rect 55858 144684 55864 144696
rect 50580 144656 55864 144684
rect 50580 144644 50586 144656
rect 55858 144644 55864 144656
rect 55916 144684 55922 144696
rect 56410 144684 56416 144696
rect 55916 144656 56416 144684
rect 55916 144644 55922 144656
rect 56410 144644 56416 144656
rect 56468 144644 56474 144696
rect 212350 144644 212356 144696
rect 212408 144684 212414 144696
rect 218054 144684 218060 144696
rect 212408 144656 218060 144684
rect 212408 144644 212414 144656
rect 218054 144644 218060 144656
rect 218112 144684 218118 144696
rect 218790 144684 218796 144696
rect 218112 144656 218796 144684
rect 218112 144644 218118 144656
rect 218790 144644 218796 144656
rect 218848 144644 218854 144696
rect 49234 144576 49240 144628
rect 49292 144616 49298 144628
rect 58710 144616 58716 144628
rect 49292 144588 58716 144616
rect 49292 144576 49298 144588
rect 58710 144576 58716 144588
rect 58768 144576 58774 144628
rect 53190 144508 53196 144560
rect 53248 144548 53254 144560
rect 58894 144548 58900 144560
rect 53248 144520 58900 144548
rect 53248 144508 53254 144520
rect 58894 144508 58900 144520
rect 58952 144508 58958 144560
rect 55950 144372 55956 144424
rect 56008 144412 56014 144424
rect 56318 144412 56324 144424
rect 56008 144384 56324 144412
rect 56008 144372 56014 144384
rect 56318 144372 56324 144384
rect 56376 144372 56382 144424
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 42610 70320 42616 70372
rect 42668 70360 42674 70372
rect 57606 70360 57612 70372
rect 42668 70332 57612 70360
rect 42668 70320 42674 70332
rect 57606 70320 57612 70332
rect 57664 70320 57670 70372
rect 209038 70320 209044 70372
rect 209096 70360 209102 70372
rect 216674 70360 216680 70372
rect 209096 70332 216680 70360
rect 209096 70320 209102 70332
rect 216674 70320 216680 70332
rect 216732 70320 216738 70372
rect 362310 70320 362316 70372
rect 362368 70360 362374 70372
rect 376938 70360 376944 70372
rect 362368 70332 376944 70360
rect 362368 70320 362374 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 358722 68280 358728 68332
rect 358780 68320 358786 68332
rect 376938 68320 376944 68332
rect 358780 68292 376944 68320
rect 358780 68280 358786 68292
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 358078 68144 358084 68196
rect 358136 68184 358142 68196
rect 358722 68184 358728 68196
rect 358136 68156 358728 68184
rect 358136 68144 358142 68156
rect 358722 68144 358728 68156
rect 358780 68144 358786 68196
rect 204898 67600 204904 67652
rect 204956 67640 204962 67652
rect 216674 67640 216680 67652
rect 204956 67612 216680 67640
rect 204956 67600 204962 67612
rect 216674 67600 216680 67612
rect 216732 67600 216738 67652
rect 218606 61208 218612 61260
rect 218664 61248 218670 61260
rect 219066 61248 219072 61260
rect 218664 61220 219072 61248
rect 218664 61208 218670 61220
rect 219066 61208 219072 61220
rect 219124 61208 219130 61260
rect 54386 59644 54392 59696
rect 54444 59684 54450 59696
rect 77110 59684 77116 59696
rect 54444 59656 77116 59684
rect 54444 59644 54450 59656
rect 77110 59644 77116 59656
rect 77168 59644 77174 59696
rect 218514 59644 218520 59696
rect 218572 59684 218578 59696
rect 237098 59684 237104 59696
rect 218572 59656 237104 59684
rect 218572 59644 218578 59656
rect 237098 59644 237104 59656
rect 237156 59644 237162 59696
rect 378778 59644 378784 59696
rect 378836 59684 378842 59696
rect 396074 59684 396080 59696
rect 378836 59656 396080 59684
rect 378836 59644 378842 59656
rect 396074 59644 396080 59656
rect 396132 59644 396138 59696
rect 54846 59576 54852 59628
rect 54904 59616 54910 59628
rect 83090 59616 83096 59628
rect 54904 59588 83096 59616
rect 54904 59576 54910 59588
rect 83090 59576 83096 59588
rect 83148 59576 83154 59628
rect 216950 59576 216956 59628
rect 217008 59616 217014 59628
rect 256970 59616 256976 59628
rect 217008 59588 256976 59616
rect 217008 59576 217014 59588
rect 256970 59576 256976 59588
rect 257028 59576 257034 59628
rect 378686 59576 378692 59628
rect 378744 59616 378750 59628
rect 397086 59616 397092 59628
rect 378744 59588 397092 59616
rect 378744 59576 378750 59588
rect 397086 59576 397092 59588
rect 397144 59576 397150 59628
rect 58894 59508 58900 59560
rect 58952 59548 58958 59560
rect 100754 59548 100760 59560
rect 58952 59520 100760 59548
rect 58952 59508 58958 59520
rect 100754 59508 100760 59520
rect 100812 59508 100818 59560
rect 216214 59508 216220 59560
rect 216272 59548 216278 59560
rect 255866 59548 255872 59560
rect 216272 59520 255872 59548
rect 216272 59508 216278 59520
rect 255866 59508 255872 59520
rect 255924 59508 255930 59560
rect 378962 59508 378968 59560
rect 379020 59548 379026 59560
rect 416958 59548 416964 59560
rect 379020 59520 416964 59548
rect 379020 59508 379026 59520
rect 416958 59508 416964 59520
rect 417016 59508 417022 59560
rect 54754 59440 54760 59492
rect 54812 59480 54818 59492
rect 101766 59480 101772 59492
rect 54812 59452 101772 59480
rect 54812 59440 54818 59452
rect 101766 59440 101772 59452
rect 101824 59440 101830 59492
rect 218974 59440 218980 59492
rect 219032 59480 219038 59492
rect 263870 59480 263876 59492
rect 219032 59452 263876 59480
rect 219032 59440 219038 59452
rect 263870 59440 263876 59452
rect 263928 59440 263934 59492
rect 377490 59440 377496 59492
rect 377548 59480 377554 59492
rect 423950 59480 423956 59492
rect 377548 59452 423956 59480
rect 377548 59440 377554 59452
rect 423950 59440 423956 59452
rect 424008 59440 424014 59492
rect 49510 59372 49516 59424
rect 49568 59412 49574 59424
rect 113542 59412 113548 59424
rect 49568 59384 113548 59412
rect 49568 59372 49574 59384
rect 113542 59372 113548 59384
rect 113600 59372 113606 59424
rect 215846 59372 215852 59424
rect 215904 59412 215910 59424
rect 262858 59412 262864 59424
rect 215904 59384 262864 59412
rect 215904 59372 215910 59384
rect 262858 59372 262864 59384
rect 262916 59372 262922 59424
rect 358170 59372 358176 59424
rect 358228 59412 358234 59424
rect 423490 59412 423496 59424
rect 358228 59384 423496 59412
rect 358228 59372 358234 59384
rect 423490 59372 423496 59384
rect 423548 59372 423554 59424
rect 55858 59304 55864 59356
rect 55916 59344 55922 59356
rect 84194 59344 84200 59356
rect 55916 59316 84200 59344
rect 55916 59304 55922 59316
rect 84194 59304 84200 59316
rect 84252 59304 84258 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 358078 59344 358084 59356
rect 218020 59316 358084 59344
rect 218020 59304 218026 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 379606 59304 379612 59356
rect 379664 59344 379670 59356
rect 418154 59344 418160 59356
rect 379664 59316 418160 59344
rect 379664 59304 379670 59316
rect 418154 59304 418160 59316
rect 418212 59304 418218 59356
rect 59078 59236 59084 59288
rect 59136 59276 59142 59288
rect 89990 59276 89996 59288
rect 59136 59248 89996 59276
rect 59136 59236 59142 59248
rect 89990 59236 89996 59248
rect 90048 59236 90054 59288
rect 218882 59236 218888 59288
rect 218940 59276 218946 59288
rect 258074 59276 258080 59288
rect 218940 59248 258080 59276
rect 218940 59236 218946 59248
rect 258074 59236 258080 59248
rect 258132 59236 258138 59288
rect 371878 59236 371884 59288
rect 371936 59276 371942 59288
rect 410702 59276 410708 59288
rect 371936 59248 410708 59276
rect 371936 59236 371942 59248
rect 410702 59236 410708 59248
rect 410760 59236 410766 59288
rect 59814 59168 59820 59220
rect 59872 59208 59878 59220
rect 94498 59208 94504 59220
rect 59872 59180 94504 59208
rect 59872 59168 59878 59180
rect 94498 59168 94504 59180
rect 94556 59168 94562 59220
rect 214282 59168 214288 59220
rect 214340 59208 214346 59220
rect 260650 59208 260656 59220
rect 214340 59180 260656 59208
rect 214340 59168 214346 59180
rect 260650 59168 260656 59180
rect 260708 59168 260714 59220
rect 376202 59168 376208 59220
rect 376260 59208 376266 59220
rect 419442 59208 419448 59220
rect 376260 59180 419448 59208
rect 376260 59168 376266 59180
rect 419442 59168 419448 59180
rect 419500 59168 419506 59220
rect 56870 59100 56876 59152
rect 56928 59140 56934 59152
rect 95878 59140 95884 59152
rect 56928 59112 95884 59140
rect 56928 59100 56934 59112
rect 95878 59100 95884 59112
rect 95936 59100 95942 59152
rect 214742 59100 214748 59152
rect 214800 59140 214806 59152
rect 261754 59140 261760 59152
rect 214800 59112 261760 59140
rect 214800 59100 214806 59112
rect 261754 59100 261760 59112
rect 261812 59100 261818 59152
rect 279234 59100 279240 59152
rect 279292 59140 279298 59152
rect 356606 59140 356612 59152
rect 279292 59112 356612 59140
rect 279292 59100 279298 59112
rect 356606 59100 356612 59112
rect 356664 59100 356670 59152
rect 375742 59100 375748 59152
rect 375800 59140 375806 59152
rect 420638 59140 420644 59152
rect 375800 59112 420644 59140
rect 375800 59100 375806 59112
rect 420638 59100 420644 59112
rect 420696 59100 420702 59152
rect 56502 59032 56508 59084
rect 56560 59072 56566 59084
rect 96982 59072 96988 59084
rect 56560 59044 96988 59072
rect 56560 59032 56566 59044
rect 96982 59032 96988 59044
rect 97040 59032 97046 59084
rect 205174 59032 205180 59084
rect 205232 59072 205238 59084
rect 290918 59072 290924 59084
rect 205232 59044 290924 59072
rect 205232 59032 205238 59044
rect 290918 59032 290924 59044
rect 290976 59032 290982 59084
rect 376294 59032 376300 59084
rect 376352 59072 376358 59084
rect 421742 59072 421748 59084
rect 376352 59044 421748 59072
rect 376352 59032 376358 59044
rect 421742 59032 421748 59044
rect 421800 59032 421806 59084
rect 54662 58964 54668 59016
rect 54720 59004 54726 59016
rect 98086 59004 98092 59016
rect 54720 58976 98092 59004
rect 54720 58964 54726 58976
rect 98086 58964 98092 58976
rect 98144 58964 98150 59016
rect 213822 58964 213828 59016
rect 213880 59004 213886 59016
rect 300854 59004 300860 59016
rect 213880 58976 300860 59004
rect 213880 58964 213886 58976
rect 300854 58964 300860 58976
rect 300912 58964 300918 59016
rect 360838 58964 360844 59016
rect 360896 59004 360902 59016
rect 416038 59004 416044 59016
rect 360896 58976 416044 59004
rect 360896 58964 360902 58976
rect 416038 58964 416044 58976
rect 416096 58964 416102 59016
rect 56226 58896 56232 58948
rect 56284 58936 56290 58948
rect 102778 58936 102784 58948
rect 56284 58908 102784 58936
rect 56284 58896 56290 58908
rect 102778 58896 102784 58908
rect 102836 58896 102842 58948
rect 212442 58896 212448 58948
rect 212500 58936 212506 58948
rect 315850 58936 315856 58948
rect 212500 58908 315856 58936
rect 212500 58896 212506 58908
rect 315850 58896 315856 58908
rect 315908 58896 315914 58948
rect 356698 58896 356704 58948
rect 356756 58936 356762 58948
rect 425974 58936 425980 58948
rect 356756 58908 425980 58936
rect 356756 58896 356762 58908
rect 425974 58896 425980 58908
rect 426032 58896 426038 58948
rect 58986 58828 58992 58880
rect 59044 58868 59050 58880
rect 107562 58868 107568 58880
rect 59044 58840 107568 58868
rect 59044 58828 59050 58840
rect 107562 58828 107568 58840
rect 107620 58828 107626 58880
rect 202782 58828 202788 58880
rect 202840 58868 202846 58880
rect 308490 58868 308496 58880
rect 202840 58840 308496 58868
rect 202840 58828 202846 58840
rect 308490 58828 308496 58840
rect 308548 58828 308554 58880
rect 369118 58828 369124 58880
rect 369176 58868 369182 58880
rect 458450 58868 458456 58880
rect 369176 58840 458456 58868
rect 369176 58828 369182 58840
rect 458450 58828 458456 58840
rect 458508 58828 458514 58880
rect 48774 58760 48780 58812
rect 48832 58800 48838 58812
rect 110966 58800 110972 58812
rect 48832 58772 110972 58800
rect 48832 58760 48838 58772
rect 110966 58760 110972 58772
rect 111024 58760 111030 58812
rect 206922 58760 206928 58812
rect 206980 58800 206986 58812
rect 320910 58800 320916 58812
rect 206980 58772 320916 58800
rect 206980 58760 206986 58772
rect 320910 58760 320916 58772
rect 320968 58760 320974 58812
rect 362218 58760 362224 58812
rect 362276 58800 362282 58812
rect 453390 58800 453396 58812
rect 362276 58772 453396 58800
rect 362276 58760 362282 58772
rect 453390 58760 453396 58772
rect 453448 58760 453454 58812
rect 53282 58692 53288 58744
rect 53340 58732 53346 58744
rect 148502 58732 148508 58744
rect 53340 58704 148508 58732
rect 53340 58692 53346 58704
rect 148502 58692 148508 58704
rect 148560 58692 148566 58744
rect 205358 58692 205364 58744
rect 205416 58732 205422 58744
rect 325878 58732 325884 58744
rect 205416 58704 325884 58732
rect 205416 58692 205422 58704
rect 325878 58692 325884 58704
rect 325936 58692 325942 58744
rect 364978 58692 364984 58744
rect 365036 58732 365042 58744
rect 475838 58732 475844 58744
rect 365036 58704 475844 58732
rect 365036 58692 365042 58704
rect 475838 58692 475844 58704
rect 475896 58692 475902 58744
rect 50982 58624 50988 58676
rect 51040 58664 51046 58676
rect 150894 58664 150900 58676
rect 51040 58636 150900 58664
rect 51040 58624 51046 58636
rect 150894 58624 150900 58636
rect 150952 58624 150958 58676
rect 219250 58624 219256 58676
rect 219308 58664 219314 58676
rect 428182 58664 428188 58676
rect 219308 58636 428188 58664
rect 219308 58624 219314 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 374822 58556 374828 58608
rect 374880 58596 374886 58608
rect 404170 58596 404176 58608
rect 374880 58568 404176 58596
rect 374880 58556 374886 58568
rect 404170 58556 404176 58568
rect 404228 58556 404234 58608
rect 375834 58420 375840 58472
rect 375892 58460 375898 58472
rect 403066 58460 403072 58472
rect 375892 58432 403072 58460
rect 375892 58420 375898 58432
rect 403066 58420 403072 58432
rect 403124 58420 403130 58472
rect 57882 57876 57888 57928
rect 57940 57916 57946 57928
rect 204898 57916 204904 57928
rect 57940 57888 204904 57916
rect 57940 57876 57946 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 210234 57876 210240 57928
rect 210292 57916 210298 57928
rect 323302 57916 323308 57928
rect 210292 57888 323308 57916
rect 210292 57876 210298 57888
rect 323302 57876 323308 57888
rect 323360 57876 323366 57928
rect 343174 57876 343180 57928
rect 343232 57916 343238 57928
rect 357618 57916 357624 57928
rect 343232 57888 357624 57916
rect 343232 57876 343238 57888
rect 357618 57876 357624 57888
rect 357676 57876 357682 57928
rect 376662 57876 376668 57928
rect 376720 57916 376726 57928
rect 485958 57916 485964 57928
rect 376720 57888 485964 57916
rect 376720 57876 376726 57888
rect 485958 57876 485964 57888
rect 486016 57876 486022 57928
rect 503346 57876 503352 57928
rect 503404 57916 503410 57928
rect 517606 57916 517612 57928
rect 503404 57888 517612 57916
rect 503404 57876 503410 57888
rect 517606 57876 517612 57888
rect 517664 57876 517670 57928
rect 52362 57808 52368 57860
rect 52420 57848 52426 57860
rect 145558 57848 145564 57860
rect 52420 57820 145564 57848
rect 52420 57808 52426 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183462 57808 183468 57860
rect 183520 57848 183526 57860
rect 197446 57848 197452 57860
rect 183520 57820 197452 57848
rect 183520 57808 183526 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 208302 57808 208308 57860
rect 208360 57848 208366 57860
rect 313366 57848 313372 57860
rect 208360 57820 313372 57848
rect 208360 57808 208366 57820
rect 313366 57808 313372 57820
rect 313424 57808 313430 57860
rect 343450 57808 343456 57860
rect 343508 57848 343514 57860
rect 356790 57848 356796 57860
rect 343508 57820 356796 57848
rect 343508 57808 343514 57820
rect 356790 57808 356796 57820
rect 356848 57808 356854 57860
rect 366358 57808 366364 57860
rect 366416 57848 366422 57860
rect 470870 57848 470876 57860
rect 366416 57820 470876 57848
rect 366416 57808 366422 57820
rect 470870 57808 470876 57820
rect 470928 57808 470934 57860
rect 503254 57808 503260 57860
rect 503312 57848 503318 57860
rect 517974 57848 517980 57860
rect 503312 57820 517980 57848
rect 503312 57808 503318 57820
rect 517974 57808 517980 57820
rect 518032 57808 518038 57860
rect 53742 57740 53748 57792
rect 53800 57780 53806 57792
rect 133414 57780 133420 57792
rect 53800 57752 133420 57780
rect 53800 57740 53806 57752
rect 133414 57740 133420 57752
rect 133472 57740 133478 57792
rect 183186 57740 183192 57792
rect 183244 57780 183250 57792
rect 197354 57780 197360 57792
rect 183244 57752 197360 57780
rect 183244 57740 183250 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 218698 57740 218704 57792
rect 218756 57780 218762 57792
rect 318242 57780 318248 57792
rect 218756 57752 318248 57780
rect 218756 57740 218762 57752
rect 318242 57740 318248 57752
rect 318300 57740 318306 57792
rect 361482 57740 361488 57792
rect 361540 57780 361546 57792
rect 465902 57780 465908 57792
rect 361540 57752 465908 57780
rect 361540 57740 361546 57752
rect 465902 57740 465908 57752
rect 465960 57740 465966 57792
rect 52270 57672 52276 57724
rect 52328 57712 52334 57724
rect 130838 57712 130844 57724
rect 52328 57684 130844 57712
rect 52328 57672 52334 57684
rect 130838 57672 130844 57684
rect 130896 57672 130902 57724
rect 215110 57672 215116 57724
rect 215168 57712 215174 57724
rect 310974 57712 310980 57724
rect 215168 57684 310980 57712
rect 215168 57672 215174 57684
rect 310974 57672 310980 57684
rect 311032 57672 311038 57724
rect 378502 57672 378508 57724
rect 378560 57712 378566 57724
rect 478414 57712 478420 57724
rect 378560 57684 478420 57712
rect 378560 57672 378566 57684
rect 478414 57672 478420 57684
rect 478472 57672 478478 57724
rect 42702 57604 42708 57656
rect 42760 57644 42766 57656
rect 115934 57644 115940 57656
rect 42760 57616 115940 57644
rect 42760 57604 42766 57616
rect 115934 57604 115940 57616
rect 115992 57604 115998 57656
rect 216582 57604 216588 57656
rect 216640 57644 216646 57656
rect 305822 57644 305828 57656
rect 216640 57616 305828 57644
rect 216640 57604 216646 57616
rect 305822 57604 305828 57616
rect 305880 57604 305886 57656
rect 371142 57604 371148 57656
rect 371200 57644 371206 57656
rect 460934 57644 460940 57656
rect 371200 57616 460940 57644
rect 371200 57604 371206 57616
rect 460934 57604 460940 57616
rect 460992 57604 460998 57656
rect 56410 57536 56416 57588
rect 56468 57576 56474 57588
rect 103790 57576 103796 57588
rect 56468 57548 103796 57576
rect 56468 57536 56474 57548
rect 103790 57536 103796 57548
rect 103848 57536 103854 57588
rect 215202 57536 215208 57588
rect 215260 57576 215266 57588
rect 303430 57576 303436 57588
rect 215260 57548 303436 57576
rect 215260 57536 215266 57548
rect 303430 57536 303436 57548
rect 303488 57536 303494 57588
rect 363782 57536 363788 57588
rect 363840 57576 363846 57588
rect 450998 57576 451004 57588
rect 363840 57548 451004 57576
rect 363840 57536 363846 57548
rect 450998 57536 451004 57548
rect 451056 57536 451062 57588
rect 56134 57468 56140 57520
rect 56192 57508 56198 57520
rect 99374 57508 99380 57520
rect 56192 57480 99380 57508
rect 56192 57468 56198 57480
rect 99374 57468 99380 57480
rect 99432 57468 99438 57520
rect 208854 57468 208860 57520
rect 208912 57508 208918 57520
rect 295886 57508 295892 57520
rect 208912 57480 295892 57508
rect 208912 57468 208918 57480
rect 295886 57468 295892 57480
rect 295944 57468 295950 57520
rect 363690 57468 363696 57520
rect 363748 57508 363754 57520
rect 445846 57508 445852 57520
rect 363748 57480 445852 57508
rect 363748 57468 363754 57480
rect 445846 57468 445852 57480
rect 445904 57468 445910 57520
rect 51442 57400 51448 57452
rect 51500 57440 51506 57452
rect 88334 57440 88340 57452
rect 51500 57412 88340 57440
rect 51500 57400 51506 57412
rect 88334 57400 88340 57412
rect 88392 57400 88398 57452
rect 218422 57400 218428 57452
rect 218480 57440 218486 57452
rect 298094 57440 298100 57452
rect 218480 57412 298100 57440
rect 218480 57400 218486 57412
rect 298094 57400 298100 57412
rect 298152 57400 298158 57452
rect 363598 57400 363604 57452
rect 363656 57440 363662 57452
rect 430942 57440 430948 57452
rect 363656 57412 430948 57440
rect 363656 57400 363662 57412
rect 430942 57400 430948 57412
rect 431000 57400 431006 57452
rect 59262 57332 59268 57384
rect 59320 57372 59326 57384
rect 93670 57372 93676 57384
rect 59320 57344 93676 57372
rect 59320 57332 59326 57344
rect 93670 57332 93676 57344
rect 93728 57332 93734 57384
rect 205542 57332 205548 57384
rect 205600 57372 205606 57384
rect 278314 57372 278320 57384
rect 205600 57344 278320 57372
rect 205600 57332 205606 57344
rect 278314 57332 278320 57344
rect 278372 57332 278378 57384
rect 367738 57332 367744 57384
rect 367796 57372 367802 57384
rect 435910 57372 435916 57384
rect 367796 57344 435916 57372
rect 367796 57332 367802 57344
rect 435910 57332 435916 57344
rect 435968 57332 435974 57384
rect 59170 57264 59176 57316
rect 59228 57304 59234 57316
rect 90726 57304 90732 57316
rect 59228 57276 90732 57304
rect 59228 57264 59234 57276
rect 90726 57264 90732 57276
rect 90784 57264 90790 57316
rect 218606 57264 218612 57316
rect 218664 57304 218670 57316
rect 258350 57304 258356 57316
rect 218664 57276 258356 57304
rect 218664 57264 218670 57276
rect 258350 57264 258356 57276
rect 258408 57264 258414 57316
rect 374638 57264 374644 57316
rect 374696 57304 374702 57316
rect 438486 57304 438492 57316
rect 374696 57276 438492 57304
rect 374696 57264 374702 57276
rect 438486 57264 438492 57276
rect 438544 57264 438550 57316
rect 52086 57196 52092 57248
rect 52144 57236 52150 57248
rect 78214 57236 78220 57248
rect 52144 57208 78220 57236
rect 52144 57196 52150 57208
rect 78214 57196 78220 57208
rect 78272 57196 78278 57248
rect 210418 57196 210424 57248
rect 210476 57236 210482 57248
rect 248230 57236 248236 57248
rect 210476 57208 248236 57236
rect 210476 57196 210482 57208
rect 248230 57196 248236 57208
rect 248288 57196 248294 57248
rect 378870 57196 378876 57248
rect 378928 57236 378934 57248
rect 415486 57236 415492 57248
rect 378928 57208 415492 57236
rect 378928 57196 378934 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 57238 57128 57244 57180
rect 57296 57168 57302 57180
rect 57882 57168 57888 57180
rect 57296 57140 57888 57168
rect 57296 57128 57302 57140
rect 57882 57128 57888 57140
rect 57940 57128 57946 57180
rect 76006 57168 76012 57180
rect 64846 57140 76012 57168
rect 54938 57060 54944 57112
rect 54996 57100 55002 57112
rect 64846 57100 64874 57140
rect 76006 57128 76012 57140
rect 76064 57128 76070 57180
rect 54996 57072 64874 57100
rect 54996 57060 55002 57072
rect 53374 56516 53380 56568
rect 53432 56556 53438 56568
rect 115750 56556 115756 56568
rect 53432 56528 115756 56556
rect 53432 56516 53438 56528
rect 115750 56516 115756 56528
rect 115808 56516 115814 56568
rect 219986 56516 219992 56568
rect 220044 56556 220050 56568
rect 408310 56556 408316 56568
rect 220044 56528 408316 56556
rect 220044 56516 220050 56528
rect 408310 56516 408316 56528
rect 408368 56516 408374 56568
rect 50798 56448 50804 56500
rect 50856 56488 50862 56500
rect 111150 56488 111156 56500
rect 50856 56460 111156 56488
rect 50856 56448 50862 56460
rect 111150 56448 111156 56460
rect 111208 56448 111214 56500
rect 215018 56448 215024 56500
rect 215076 56488 215082 56500
rect 276934 56488 276940 56500
rect 215076 56460 276940 56488
rect 215076 56448 215082 56460
rect 276934 56448 276940 56460
rect 276992 56448 276998 56500
rect 375650 56448 375656 56500
rect 375708 56488 375714 56500
rect 436278 56488 436284 56500
rect 375708 56460 436284 56488
rect 375708 56448 375714 56460
rect 436278 56448 436284 56460
rect 436336 56448 436342 56500
rect 53466 56380 53472 56432
rect 53524 56420 53530 56432
rect 112070 56420 112076 56432
rect 53524 56392 112076 56420
rect 53524 56380 53530 56392
rect 112070 56380 112076 56392
rect 112128 56380 112134 56432
rect 219066 56380 219072 56432
rect 219124 56420 219130 56432
rect 235994 56420 236000 56432
rect 219124 56392 236000 56420
rect 219124 56380 219130 56392
rect 235994 56380 236000 56392
rect 236052 56380 236058 56432
rect 375282 56380 375288 56432
rect 375340 56420 375346 56432
rect 434438 56420 434444 56432
rect 375340 56392 434444 56420
rect 375340 56380 375346 56392
rect 434438 56380 434444 56392
rect 434496 56380 434502 56432
rect 59906 56312 59912 56364
rect 59964 56352 59970 56364
rect 108206 56352 108212 56364
rect 59964 56324 108212 56352
rect 59964 56312 59970 56324
rect 108206 56312 108212 56324
rect 108264 56312 108270 56364
rect 213362 56312 213368 56364
rect 213420 56352 213426 56364
rect 273254 56352 273260 56364
rect 213420 56324 273260 56352
rect 213420 56312 213426 56324
rect 273254 56312 273260 56324
rect 273312 56312 273318 56364
rect 374546 56312 374552 56364
rect 374604 56352 374610 56364
rect 432230 56352 432236 56364
rect 374604 56324 432236 56352
rect 374604 56312 374610 56324
rect 432230 56312 432236 56324
rect 432288 56312 432294 56364
rect 58710 56244 58716 56296
rect 58768 56284 58774 56296
rect 93302 56284 93308 56296
rect 58768 56256 93308 56284
rect 58768 56244 58774 56256
rect 93302 56244 93308 56256
rect 93360 56244 93366 56296
rect 214650 56244 214656 56296
rect 214708 56284 214714 56296
rect 271046 56284 271052 56296
rect 214708 56256 271052 56284
rect 214708 56244 214714 56256
rect 271046 56244 271052 56256
rect 271104 56244 271110 56296
rect 379330 56244 379336 56296
rect 379388 56284 379394 56296
rect 427630 56284 427636 56296
rect 379388 56256 427636 56284
rect 379388 56244 379394 56256
rect 427630 56244 427636 56256
rect 427688 56244 427694 56296
rect 56318 56176 56324 56228
rect 56376 56216 56382 56228
rect 88702 56216 88708 56228
rect 56376 56188 88708 56216
rect 56376 56176 56382 56188
rect 88702 56176 88708 56188
rect 88760 56176 88766 56228
rect 219894 56176 219900 56228
rect 219952 56216 219958 56228
rect 268102 56216 268108 56228
rect 219952 56188 268108 56216
rect 219952 56176 219958 56188
rect 268102 56176 268108 56188
rect 268160 56176 268166 56228
rect 379882 56176 379888 56228
rect 379940 56216 379946 56228
rect 414566 56216 414572 56228
rect 379940 56188 414572 56216
rect 379940 56176 379946 56188
rect 414566 56176 414572 56188
rect 414624 56176 414630 56228
rect 54478 56108 54484 56160
rect 54536 56148 54542 56160
rect 86494 56148 86500 56160
rect 54536 56120 86500 56148
rect 54536 56108 54542 56120
rect 86494 56108 86500 56120
rect 86552 56108 86558 56160
rect 218238 56108 218244 56160
rect 218296 56148 218302 56160
rect 266354 56148 266360 56160
rect 218296 56120 266360 56148
rect 218296 56108 218302 56120
rect 266354 56108 266360 56120
rect 266412 56108 266418 56160
rect 379054 56108 379060 56160
rect 379112 56148 379118 56160
rect 412634 56148 412640 56160
rect 379112 56120 412640 56148
rect 379112 56108 379118 56120
rect 412634 56108 412640 56120
rect 412692 56108 412698 56160
rect 58802 56040 58808 56092
rect 58860 56080 58866 56092
rect 85390 56080 85396 56092
rect 58860 56052 85396 56080
rect 58860 56040 58866 56052
rect 85390 56040 85396 56052
rect 85448 56040 85454 56092
rect 219342 56040 219348 56092
rect 219400 56080 219406 56092
rect 253382 56080 253388 56092
rect 219400 56052 253388 56080
rect 219400 56040 219406 56052
rect 253382 56040 253388 56052
rect 253440 56040 253446 56092
rect 375926 56040 375932 56092
rect 375984 56080 375990 56092
rect 408678 56080 408684 56092
rect 375984 56052 408684 56080
rect 375984 56040 375990 56052
rect 408678 56040 408684 56052
rect 408736 56040 408742 56092
rect 55030 55972 55036 56024
rect 55088 56012 55094 56024
rect 80422 56012 80428 56024
rect 55088 55984 80428 56012
rect 55088 55972 55094 55984
rect 80422 55972 80428 55984
rect 80480 55972 80486 56024
rect 219158 55972 219164 56024
rect 219216 56012 219222 56024
rect 251174 56012 251180 56024
rect 219216 55984 251180 56012
rect 219216 55972 219222 55984
rect 251174 55972 251180 55984
rect 251232 55972 251238 56024
rect 379422 55972 379428 56024
rect 379480 56012 379486 56024
rect 411254 56012 411260 56024
rect 379480 55984 411260 56012
rect 379480 55972 379486 55984
rect 411254 55972 411260 55984
rect 411312 55972 411318 56024
rect 217134 55904 217140 55956
rect 217192 55944 217198 55956
rect 248598 55944 248604 55956
rect 217192 55916 248604 55944
rect 217192 55904 217198 55916
rect 248598 55904 248604 55916
rect 248656 55904 248662 55956
rect 373350 55904 373356 55956
rect 373408 55944 373414 55956
rect 401686 55944 401692 55956
rect 373408 55916 401692 55944
rect 373408 55904 373414 55916
rect 401686 55904 401692 55916
rect 401744 55904 401750 55956
rect 213546 55836 213552 55888
rect 213604 55876 213610 55888
rect 241606 55876 241612 55888
rect 213604 55848 241612 55876
rect 213604 55836 213610 55848
rect 241606 55836 241612 55848
rect 241664 55836 241670 55888
rect 373258 55836 373264 55888
rect 373316 55876 373322 55888
rect 399478 55876 399484 55888
rect 373316 55848 399484 55876
rect 373316 55836 373322 55848
rect 399478 55836 399484 55848
rect 399536 55836 399542 55888
rect 216030 55768 216036 55820
rect 216088 55808 216094 55820
rect 245286 55808 245292 55820
rect 216088 55780 245292 55808
rect 216088 55768 216094 55780
rect 245286 55768 245292 55780
rect 245344 55768 245350 55820
rect 213178 55700 213184 55752
rect 213236 55740 213242 55752
rect 239214 55740 239220 55752
rect 213236 55712 239220 55740
rect 213236 55700 213242 55712
rect 239214 55700 239220 55712
rect 239272 55700 239278 55752
rect 213730 55632 213736 55684
rect 213788 55672 213794 55684
rect 275094 55672 275100 55684
rect 213788 55644 275100 55672
rect 213788 55632 213794 55644
rect 275094 55632 275100 55644
rect 275152 55632 275158 55684
rect 53098 55156 53104 55208
rect 53156 55196 53162 55208
rect 78674 55196 78680 55208
rect 53156 55168 78680 55196
rect 53156 55156 53162 55168
rect 78674 55156 78680 55168
rect 78732 55156 78738 55208
rect 216398 55156 216404 55208
rect 216456 55196 216462 55208
rect 242894 55196 242900 55208
rect 216456 55168 242900 55196
rect 216456 55156 216462 55168
rect 242894 55156 242900 55168
rect 242952 55156 242958 55208
rect 379238 55156 379244 55208
rect 379296 55196 379302 55208
rect 405826 55196 405832 55208
rect 379296 55168 405832 55196
rect 379296 55156 379302 55168
rect 405826 55156 405832 55168
rect 405884 55156 405890 55208
rect 54018 55088 54024 55140
rect 54076 55128 54082 55140
rect 116118 55128 116124 55140
rect 54076 55100 116124 55128
rect 54076 55088 54082 55100
rect 116118 55088 116124 55100
rect 116176 55088 116182 55140
rect 214558 55088 214564 55140
rect 214616 55128 214622 55140
rect 240134 55128 240140 55140
rect 214616 55100 240140 55128
rect 214616 55088 214622 55100
rect 240134 55088 240140 55100
rect 240192 55088 240198 55140
rect 374730 55088 374736 55140
rect 374788 55128 374794 55140
rect 400214 55128 400220 55140
rect 374788 55100 400220 55128
rect 374788 55088 374794 55100
rect 400214 55088 400220 55100
rect 400272 55088 400278 55140
rect 53558 55020 53564 55072
rect 53616 55060 53622 55072
rect 113174 55060 113180 55072
rect 53616 55032 113180 55060
rect 53616 55020 53622 55032
rect 113174 55020 113180 55032
rect 113232 55020 113238 55072
rect 215938 55020 215944 55072
rect 215996 55060 216002 55072
rect 271874 55060 271880 55072
rect 215996 55032 271880 55060
rect 215996 55020 216002 55032
rect 271874 55020 271880 55032
rect 271932 55020 271938 55072
rect 373810 55020 373816 55072
rect 373868 55060 373874 55072
rect 433426 55060 433432 55072
rect 373868 55032 433432 55060
rect 373868 55020 373874 55032
rect 433426 55020 433432 55032
rect 433484 55020 433490 55072
rect 53006 54952 53012 55004
rect 53064 54992 53070 55004
rect 113266 54992 113272 55004
rect 53064 54964 113272 54992
rect 53064 54952 53070 54964
rect 113266 54952 113272 54964
rect 113324 54952 113330 55004
rect 219526 54952 219532 55004
rect 219584 54992 219590 55004
rect 266446 54992 266452 55004
rect 219584 54964 266452 54992
rect 219584 54952 219590 54964
rect 266446 54952 266452 54964
rect 266504 54952 266510 55004
rect 375098 54952 375104 55004
rect 375156 54992 375162 55004
rect 430574 54992 430580 55004
rect 375156 54964 430580 54992
rect 375156 54952 375162 54964
rect 430574 54952 430580 54964
rect 430632 54952 430638 55004
rect 50890 54884 50896 54936
rect 50948 54924 50954 54936
rect 109034 54924 109040 54936
rect 50948 54896 109040 54924
rect 50948 54884 50954 54896
rect 109034 54884 109040 54896
rect 109092 54884 109098 54936
rect 219618 54884 219624 54936
rect 219676 54924 219682 54936
rect 264974 54924 264980 54936
rect 219676 54896 264980 54924
rect 219676 54884 219682 54896
rect 264974 54884 264980 54896
rect 265032 54884 265038 54936
rect 375190 54884 375196 54936
rect 375248 54924 375254 54936
rect 429194 54924 429200 54936
rect 375248 54896 429200 54924
rect 375248 54884 375254 54896
rect 429194 54884 429200 54896
rect 429252 54884 429258 54936
rect 59998 54816 60004 54868
rect 60056 54856 60062 54868
rect 106274 54856 106280 54868
rect 60056 54828 106280 54856
rect 60056 54816 60062 54828
rect 106274 54816 106280 54828
rect 106332 54816 106338 54868
rect 219802 54816 219808 54868
rect 219860 54856 219866 54868
rect 253934 54856 253940 54868
rect 219860 54828 253940 54856
rect 219860 54816 219866 54828
rect 253934 54816 253940 54828
rect 253992 54816 253998 54868
rect 379974 54816 379980 54868
rect 380032 54856 380038 54868
rect 427814 54856 427820 54868
rect 380032 54828 427820 54856
rect 380032 54816 380038 54828
rect 427814 54816 427820 54828
rect 427872 54816 427878 54868
rect 57054 54748 57060 54800
rect 57112 54788 57118 54800
rect 91094 54788 91100 54800
rect 57112 54760 91100 54788
rect 57112 54748 57118 54760
rect 91094 54748 91100 54760
rect 91152 54748 91158 54800
rect 217226 54748 217232 54800
rect 217284 54788 217290 54800
rect 251358 54788 251364 54800
rect 217284 54760 251364 54788
rect 217284 54748 217290 54760
rect 251358 54748 251364 54760
rect 251416 54748 251422 54800
rect 379698 54748 379704 54800
rect 379756 54788 379762 54800
rect 426526 54788 426532 54800
rect 379756 54760 426532 54788
rect 379756 54748 379762 54760
rect 426526 54748 426532 54760
rect 426584 54748 426590 54800
rect 53650 54680 53656 54732
rect 53708 54720 53714 54732
rect 86954 54720 86960 54732
rect 53708 54692 86960 54720
rect 53708 54680 53714 54692
rect 86954 54680 86960 54692
rect 87012 54680 87018 54732
rect 216490 54680 216496 54732
rect 216548 54720 216554 54732
rect 249794 54720 249800 54732
rect 216548 54692 249800 54720
rect 216548 54680 216554 54692
rect 249794 54680 249800 54692
rect 249852 54680 249858 54732
rect 378042 54680 378048 54732
rect 378100 54720 378106 54732
rect 411346 54720 411352 54732
rect 378100 54692 411352 54720
rect 378100 54680 378106 54692
rect 411346 54680 411352 54692
rect 411404 54680 411410 54732
rect 58618 54612 58624 54664
rect 58676 54652 58682 54664
rect 91462 54652 91468 54664
rect 58676 54624 91468 54652
rect 58676 54612 58682 54624
rect 91462 54612 91468 54624
rect 91520 54612 91526 54664
rect 216122 54612 216128 54664
rect 216180 54652 216186 54664
rect 247034 54652 247040 54664
rect 216180 54624 247040 54652
rect 216180 54612 216186 54624
rect 247034 54612 247040 54624
rect 247092 54612 247098 54664
rect 377306 54612 377312 54664
rect 377364 54652 377370 54664
rect 409874 54652 409880 54664
rect 377364 54624 409880 54652
rect 377364 54612 377370 54624
rect 409874 54612 409880 54624
rect 409932 54612 409938 54664
rect 52178 54544 52184 54596
rect 52236 54584 52242 54596
rect 81434 54584 81440 54596
rect 52236 54556 81440 54584
rect 52236 54544 52242 54556
rect 81434 54544 81440 54556
rect 81492 54544 81498 54596
rect 214926 54544 214932 54596
rect 214984 54584 214990 54596
rect 244366 54584 244372 54596
rect 214984 54556 244372 54584
rect 214984 54544 214990 54556
rect 244366 54544 244372 54556
rect 244424 54544 244430 54596
rect 376110 54544 376116 54596
rect 376168 54584 376174 54596
rect 407206 54584 407212 54596
rect 376168 54556 407212 54584
rect 376168 54544 376174 54556
rect 407206 54544 407212 54556
rect 407264 54544 407270 54596
rect 44082 54476 44088 54528
rect 44140 54516 44146 54528
rect 122834 54516 122840 54528
rect 44140 54488 122840 54516
rect 44140 54476 44146 54488
rect 122834 54476 122840 54488
rect 122892 54476 122898 54528
rect 218790 54476 218796 54528
rect 218848 54516 218854 54528
rect 245654 54516 245660 54528
rect 218848 54488 245660 54516
rect 218848 54476 218854 54488
rect 245654 54476 245660 54488
rect 245712 54476 245718 54528
rect 376478 54476 376484 54528
rect 376536 54516 376542 54528
rect 404354 54516 404360 54528
rect 376536 54488 404360 54516
rect 376536 54476 376542 54488
rect 404354 54476 404360 54488
rect 404412 54476 404418 54528
rect 216306 54408 216312 54460
rect 216364 54448 216370 54460
rect 277394 54448 277400 54460
rect 216364 54420 277400 54448
rect 216364 54408 216370 54420
rect 277394 54408 277400 54420
rect 277452 54408 277458 54460
rect 375558 54408 375564 54460
rect 375616 54448 375622 54460
rect 437474 54448 437480 54460
rect 375616 54420 437480 54448
rect 375616 54408 375622 54420
rect 437474 54408 437480 54420
rect 437532 54408 437538 54460
rect 213454 54340 213460 54392
rect 213512 54380 213518 54392
rect 273346 54380 273352 54392
rect 213512 54352 273352 54380
rect 213512 54340 213518 54352
rect 273346 54340 273352 54352
rect 273404 54340 273410 54392
rect 374270 54340 374276 54392
rect 374328 54380 374334 54392
rect 434714 54380 434720 54392
rect 374328 54352 434720 54380
rect 374328 54340 374334 54352
rect 434714 54340 434720 54352
rect 434772 54340 434778 54392
rect 213270 54272 213276 54324
rect 213328 54312 213334 54324
rect 237374 54312 237380 54324
rect 213328 54284 237380 54312
rect 213328 54272 213334 54284
rect 237374 54272 237380 54284
rect 237432 54272 237438 54324
rect 373718 54272 373724 54324
rect 373776 54312 373782 54324
rect 397454 54312 397460 54324
rect 373776 54284 397460 54312
rect 373776 54272 373782 54284
rect 397454 54272 397460 54284
rect 397512 54272 397518 54324
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 10318 20652 10324 20664
rect 3476 20624 10324 20652
rect 3476 20612 3482 20624
rect 10318 20612 10324 20624
rect 10376 20612 10382 20664
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 125870 2796 125876 2848
rect 125928 2836 125934 2848
rect 365714 2836 365720 2848
rect 125928 2808 365720 2836
rect 125928 2796 125934 2808
rect 365714 2796 365720 2808
rect 365772 2796 365778 2848
<< via1 >>
rect 235172 700408 235224 700460
rect 305644 700408 305696 700460
rect 429844 700408 429896 700460
rect 434720 700408 434772 700460
rect 170312 700340 170364 700392
rect 434812 700340 434864 700392
rect 57704 700272 57756 700324
rect 543464 700272 543516 700324
rect 147220 683136 147272 683188
rect 580172 683136 580224 683188
rect 104900 647844 104952 647896
rect 434904 647844 434956 647896
rect 299480 646484 299532 646536
rect 405924 646484 405976 646536
rect 364340 645124 364392 645176
rect 428372 645124 428424 645176
rect 322572 643084 322624 643136
rect 436100 643084 436152 643136
rect 322480 642676 322532 642728
rect 346584 642676 346636 642728
rect 323676 642608 323728 642660
rect 401692 642608 401744 642660
rect 316776 642540 316828 642592
rect 342260 642540 342312 642592
rect 309784 642472 309836 642524
rect 374000 642472 374052 642524
rect 323768 642404 323820 642456
rect 369124 642404 369176 642456
rect 318156 642336 318208 642388
rect 364616 642336 364668 642388
rect 324872 642268 324924 642320
rect 378140 642268 378192 642320
rect 322296 642200 322348 642252
rect 355600 642200 355652 642252
rect 355692 642200 355744 642252
rect 414848 642200 414900 642252
rect 307024 642132 307076 642184
rect 337568 642132 337620 642184
rect 347596 642132 347648 642184
rect 410340 642132 410392 642184
rect 323952 642064 324004 642116
rect 387800 642064 387852 642116
rect 320916 641996 320968 642048
rect 392308 641996 392360 642048
rect 311164 641928 311216 641980
rect 383660 641928 383712 641980
rect 337108 641860 337160 641912
rect 351092 641860 351144 641912
rect 322388 641792 322440 641844
rect 432880 641792 432932 641844
rect 323860 641724 323912 641776
rect 328552 641724 328604 641776
rect 365628 641724 365680 641776
rect 419540 641724 419592 641776
rect 457444 641724 457496 641776
rect 319444 641180 319496 641232
rect 436192 641180 436244 641232
rect 233240 641112 233292 641164
rect 360200 641112 360252 641164
rect 147588 641044 147640 641096
rect 164516 641044 164568 641096
rect 324228 641044 324280 641096
rect 494060 641044 494112 641096
rect 131120 640976 131172 641028
rect 161572 640976 161624 641028
rect 238024 640976 238076 641028
rect 365628 640976 365680 641028
rect 145012 640908 145064 640960
rect 207664 640908 207716 640960
rect 239496 640908 239548 640960
rect 257436 640908 257488 640960
rect 323584 640908 323636 640960
rect 457628 640908 457680 640960
rect 115388 640840 115440 640892
rect 124680 640840 124732 640892
rect 148876 640840 148928 640892
rect 172888 640840 172940 640892
rect 235264 640840 235316 640892
rect 292212 640840 292264 640892
rect 322664 640840 322716 640892
rect 457720 640840 457772 640892
rect 69020 640704 69072 640756
rect 124404 640772 124456 640824
rect 140780 640772 140832 640824
rect 167092 640772 167144 640824
rect 226340 640772 226392 640824
rect 300584 640772 300636 640824
rect 314108 640772 314160 640824
rect 457812 640772 457864 640824
rect 117964 640704 118016 640756
rect 124496 640704 124548 640756
rect 148784 640704 148836 640756
rect 176108 640704 176160 640756
rect 239588 640704 239640 640756
rect 274824 640704 274876 640756
rect 316684 640704 316736 640756
rect 471612 640704 471664 640756
rect 112168 640636 112220 640688
rect 122840 640636 122892 640688
rect 149520 640636 149572 640688
rect 190552 640636 190604 640688
rect 236644 640636 236696 640688
rect 396816 640636 396868 640688
rect 60740 640568 60792 640620
rect 98000 640568 98052 640620
rect 106372 640568 106424 640620
rect 121460 640568 121512 640620
rect 142160 640568 142212 640620
rect 184480 640568 184532 640620
rect 217416 640568 217468 640620
rect 254860 640568 254912 640620
rect 314016 640568 314068 640620
rect 483204 640568 483256 640620
rect 54852 640500 54904 640552
rect 88984 640500 89036 640552
rect 103796 640500 103848 640552
rect 121552 640500 121604 640552
rect 144920 640500 144972 640552
rect 196072 640500 196124 640552
rect 231124 640500 231176 640552
rect 243544 640500 243596 640552
rect 249708 640500 249760 640552
rect 295432 640500 295484 640552
rect 319536 640500 319588 640552
rect 494796 640500 494848 640552
rect 55128 640432 55180 640484
rect 92204 640432 92256 640484
rect 94780 640432 94832 640484
rect 120908 640432 120960 640484
rect 147312 640432 147364 640484
rect 199292 640432 199344 640484
rect 237380 640432 237432 640484
rect 289636 640432 289688 640484
rect 322204 640432 322256 640484
rect 501236 640432 501288 640484
rect 55036 640364 55088 640416
rect 65800 640364 65852 640416
rect 100576 640364 100628 640416
rect 117964 640364 118016 640416
rect 56508 640296 56560 640348
rect 77392 640296 77444 640348
rect 109592 640296 109644 640348
rect 121000 640364 121052 640416
rect 149612 640364 149664 640416
rect 201868 640364 201920 640416
rect 205548 640364 205600 640416
rect 212632 640364 212684 640416
rect 238116 640364 238168 640416
rect 251640 640364 251692 640416
rect 319628 640364 319680 640416
rect 512000 640364 512052 640416
rect 118240 640296 118292 640348
rect 124588 640296 124640 640348
rect 133880 640296 133932 640348
rect 149980 640296 150032 640348
rect 243544 640296 243596 640348
rect 249064 640296 249116 640348
rect 255320 640296 255372 640348
rect 263232 640296 263284 640348
rect 316868 640296 316920 640348
rect 512184 640296 512236 640348
rect 223580 639820 223632 639872
rect 249708 639820 249760 639872
rect 222200 639752 222252 639804
rect 255320 639752 255372 639804
rect 3424 639684 3476 639736
rect 337108 639684 337160 639736
rect 3608 639616 3660 639668
rect 347596 639616 347648 639668
rect 3700 639548 3752 639600
rect 355508 639548 355560 639600
rect 238944 639208 238996 639260
rect 580356 639208 580408 639260
rect 231216 639140 231268 639192
rect 272248 639140 272300 639192
rect 316960 639140 317012 639192
rect 457536 639140 457588 639192
rect 239036 639072 239088 639124
rect 433340 639072 433392 639124
rect 149888 639004 149940 639056
rect 170312 639004 170364 639056
rect 215944 639004 215996 639056
rect 269028 639004 269080 639056
rect 317052 639004 317104 639056
rect 512092 639004 512144 639056
rect 148324 638936 148376 638988
rect 153200 638936 153252 638988
rect 3516 638188 3568 638240
rect 321008 638188 321060 638240
rect 236736 638052 236788 638104
rect 245660 638052 245712 638104
rect 126244 637984 126296 638036
rect 187700 637984 187752 638036
rect 228364 637984 228416 638036
rect 266268 637984 266320 638036
rect 59360 637916 59412 637968
rect 60740 637916 60792 637968
rect 148968 637916 149020 637968
rect 158720 637916 158772 637968
rect 216036 637916 216088 637968
rect 260380 637916 260432 637968
rect 54944 637848 54996 637900
rect 62948 637848 63000 637900
rect 136640 637848 136692 637900
rect 178684 637848 178736 637900
rect 226984 637848 227036 637900
rect 283564 637848 283616 637900
rect 56416 637780 56468 637832
rect 71228 637780 71280 637832
rect 86776 637780 86828 637832
rect 125784 637780 125836 637832
rect 140044 637780 140096 637832
rect 193496 637780 193548 637832
rect 220084 637780 220136 637832
rect 280252 637780 280304 637832
rect 56324 637712 56376 637764
rect 74632 637712 74684 637764
rect 124220 637712 124272 637764
rect 182088 637712 182140 637764
rect 214564 637712 214616 637764
rect 286140 637712 286192 637764
rect 57796 637644 57848 637696
rect 80244 637644 80296 637696
rect 83464 637644 83516 637696
rect 124312 637644 124364 637696
rect 146116 637644 146168 637696
rect 155500 637644 155552 637696
rect 217324 637644 217376 637696
rect 297732 637644 297784 637696
rect 57888 637576 57940 637628
rect 146208 637576 146260 637628
rect 238024 637576 238076 637628
rect 238208 637576 238260 637628
rect 277676 637576 277728 637628
rect 239404 637508 239456 637560
rect 242900 637508 242952 637560
rect 213920 636828 213972 636880
rect 237380 636828 237432 636880
rect 144184 635196 144236 635248
rect 147128 635196 147180 635248
rect 232504 635128 232556 635180
rect 237380 635128 237432 635180
rect 465448 634856 465500 634908
rect 580264 634788 580316 634840
rect 312544 633428 312596 633480
rect 321560 633428 321612 633480
rect 238852 629960 238904 630012
rect 239772 629960 239824 630012
rect 233332 629280 233384 629332
rect 237380 629280 237432 629332
rect 313924 629280 313976 629332
rect 321560 629280 321612 629332
rect 140872 626560 140924 626612
rect 146300 626560 146352 626612
rect 216128 626560 216180 626612
rect 237380 626560 237432 626612
rect 318064 623772 318116 623824
rect 321560 623772 321612 623824
rect 132500 622412 132552 622464
rect 146300 622412 146352 622464
rect 222844 622412 222896 622464
rect 237380 622412 237432 622464
rect 223672 619624 223724 619676
rect 237380 619624 237432 619676
rect 311256 619624 311308 619676
rect 321560 619624 321612 619676
rect 218060 616836 218112 616888
rect 237380 616836 237432 616888
rect 309876 614116 309928 614168
rect 321560 614116 321612 614168
rect 314200 609968 314252 610020
rect 321560 609968 321612 610020
rect 220176 607180 220228 607232
rect 237380 607180 237432 607232
rect 311348 605820 311400 605872
rect 321560 605820 321612 605872
rect 129004 604460 129056 604512
rect 146300 604460 146352 604512
rect 235448 604460 235500 604512
rect 237380 604460 237432 604512
rect 303160 603712 303212 603764
rect 322664 603712 322716 603764
rect 124128 603100 124180 603152
rect 145564 603100 145616 603152
rect 214656 601672 214708 601724
rect 237380 601672 237432 601724
rect 123300 600992 123352 601044
rect 123484 600992 123536 601044
rect 229744 597524 229796 597576
rect 237380 597524 237432 597576
rect 304264 596164 304316 596216
rect 321560 596164 321612 596216
rect 231860 594804 231912 594856
rect 237380 594804 237432 594856
rect 125600 592016 125652 592068
rect 146300 592016 146352 592068
rect 235356 592016 235408 592068
rect 237380 592016 237432 592068
rect 307116 590656 307168 590708
rect 321560 590656 321612 590708
rect 130384 589296 130436 589348
rect 146300 589296 146352 589348
rect 233884 589296 233936 589348
rect 237380 589296 237432 589348
rect 57704 589228 57756 589280
rect 58624 589228 58676 589280
rect 139400 586508 139452 586560
rect 146300 586508 146352 586560
rect 214748 586508 214800 586560
rect 237380 586508 237432 586560
rect 309968 586508 310020 586560
rect 321560 586508 321612 586560
rect 513288 586508 513340 586560
rect 560944 586508 560996 586560
rect 226432 583720 226484 583772
rect 237380 583720 237432 583772
rect 120724 581612 120776 581664
rect 121184 581612 121236 581664
rect 305736 581000 305788 581052
rect 321560 581000 321612 581052
rect 218152 579640 218204 579692
rect 237380 579640 237432 579692
rect 216680 576852 216732 576904
rect 237380 576852 237432 576904
rect 148416 576784 148468 576836
rect 149428 576784 149480 576836
rect 57152 575696 57204 575748
rect 59912 575696 59964 575748
rect 3792 575424 3844 575476
rect 307116 575424 307168 575476
rect 145564 575356 145616 575408
rect 214012 575356 214064 575408
rect 302884 575356 302936 575408
rect 57060 575288 57112 575340
rect 62120 575288 62172 575340
rect 106280 575288 106332 575340
rect 124680 575288 124732 575340
rect 149336 575288 149388 575340
rect 151820 575288 151872 575340
rect 289820 575288 289872 575340
rect 314016 575288 314068 575340
rect 99564 575220 99616 575272
rect 122288 575220 122340 575272
rect 149704 575220 149756 575272
rect 154764 575220 154816 575272
rect 293960 575220 294012 575272
rect 319628 575220 319680 575272
rect 98092 575152 98144 575204
rect 121000 575152 121052 575204
rect 148600 575152 148652 575204
rect 150532 575152 150584 575204
rect 288532 575152 288584 575204
rect 316960 575152 317012 575204
rect 96804 575084 96856 575136
rect 122840 575084 122892 575136
rect 288440 575084 288492 575136
rect 316868 575084 316920 575136
rect 93860 575016 93912 575068
rect 124496 575016 124548 575068
rect 147312 575016 147364 575068
rect 156052 575016 156104 575068
rect 195244 575016 195296 575068
rect 212816 575016 212868 575068
rect 287060 575016 287112 575068
rect 317052 575016 317104 575068
rect 58900 574948 58952 575000
rect 74540 574948 74592 575000
rect 86960 574948 87012 575000
rect 121460 574948 121512 575000
rect 149796 574948 149848 575000
rect 160284 574948 160336 575000
rect 164332 574948 164384 575000
rect 212632 574948 212684 575000
rect 260840 574948 260892 575000
rect 319444 574948 319496 575000
rect 54852 574880 54904 574932
rect 78680 574880 78732 574932
rect 87052 574880 87104 574932
rect 124588 574880 124640 574932
rect 126980 574880 127032 574932
rect 211804 574880 211856 574932
rect 227720 574880 227772 574932
rect 300952 574880 301004 574932
rect 58716 574812 58768 574864
rect 67640 574812 67692 574864
rect 69020 574812 69072 574864
rect 122196 574812 122248 574864
rect 148784 574812 148836 574864
rect 161480 574812 161532 574864
rect 183652 574812 183704 574864
rect 301044 574812 301096 574864
rect 63500 574744 63552 574796
rect 123576 574744 123628 574796
rect 148876 574744 148928 574796
rect 164240 574744 164292 574796
rect 179420 574744 179472 574796
rect 300860 574744 300912 574796
rect 291200 574676 291252 574728
rect 314108 574676 314160 574728
rect 119344 574608 119396 574660
rect 123392 574608 123444 574660
rect 296904 574608 296956 574660
rect 319536 574608 319588 574660
rect 57428 574268 57480 574320
rect 60740 574268 60792 574320
rect 302884 574064 302936 574116
rect 303344 574064 303396 574116
rect 111892 573588 111944 573640
rect 123024 573588 123076 573640
rect 229100 573588 229152 573640
rect 303068 573588 303120 573640
rect 59084 573520 59136 573572
rect 92572 573520 92624 573572
rect 122840 573520 122892 573572
rect 211436 573520 211488 573572
rect 245660 573520 245712 573572
rect 322572 573520 322624 573572
rect 57520 573452 57572 573504
rect 82912 573452 82964 573504
rect 84200 573452 84252 573504
rect 122104 573452 122156 573504
rect 201684 573452 201736 573504
rect 302240 573452 302292 573504
rect 65064 573384 65116 573436
rect 122012 573384 122064 573436
rect 149612 573384 149664 573436
rect 158720 573384 158772 573436
rect 179512 573384 179564 573436
rect 301596 573384 301648 573436
rect 3516 573316 3568 573368
rect 324044 573316 324096 573368
rect 147128 572704 147180 572756
rect 151084 572704 151136 572756
rect 62764 572500 62816 572552
rect 65156 572500 65208 572552
rect 161572 572432 161624 572484
rect 178040 572432 178092 572484
rect 163044 572364 163096 572416
rect 183836 572364 183888 572416
rect 235540 572364 235592 572416
rect 248420 572364 248472 572416
rect 143540 572296 143592 572348
rect 166448 572296 166500 572348
rect 169852 572296 169904 572348
rect 175464 572296 175516 572348
rect 198004 572296 198056 572348
rect 201500 572296 201552 572348
rect 220820 572296 220872 572348
rect 240048 572296 240100 572348
rect 249064 572296 249116 572348
rect 271604 572296 271656 572348
rect 154672 572228 154724 572280
rect 181260 572228 181312 572280
rect 230480 572228 230532 572280
rect 260012 572228 260064 572280
rect 70952 572160 71004 572212
rect 86224 572160 86276 572212
rect 94136 572160 94188 572212
rect 104900 572160 104952 572212
rect 158812 572160 158864 572212
rect 192852 572160 192904 572212
rect 227812 572160 227864 572212
rect 265808 572160 265860 572212
rect 273904 572160 273956 572212
rect 283196 572160 283248 572212
rect 287704 572160 287756 572212
rect 300584 572160 300636 572212
rect 74632 572092 74684 572144
rect 97356 572092 97408 572144
rect 99932 572092 99984 572144
rect 115204 572092 115256 572144
rect 129740 572092 129792 572144
rect 163872 572092 163924 572144
rect 173900 572092 173952 572144
rect 189632 572092 189684 572144
rect 193864 572092 193916 572144
rect 210240 572092 210292 572144
rect 231952 572092 232004 572144
rect 279976 572092 280028 572144
rect 280804 572092 280856 572144
rect 297364 572092 297416 572144
rect 57336 572024 57388 572076
rect 79324 572024 79376 572076
rect 85764 572024 85816 572076
rect 108304 572024 108356 572076
rect 110420 572024 110472 572076
rect 121184 572024 121236 572076
rect 132592 572024 132644 572076
rect 187056 572024 187108 572076
rect 192484 572024 192536 572076
rect 213276 572024 213328 572076
rect 219440 572024 219492 572076
rect 268384 572024 268436 572076
rect 269120 572024 269172 572076
rect 309968 572024 310020 572076
rect 60004 571956 60056 572008
rect 71044 571956 71096 572008
rect 79968 571956 80020 572008
rect 114744 571956 114796 572008
rect 133972 571956 134024 572008
rect 207020 571956 207072 572008
rect 222292 571956 222344 572008
rect 274180 571956 274232 572008
rect 280160 571956 280212 572008
rect 322480 571956 322532 572008
rect 246304 571480 246356 571532
rect 250996 571480 251048 571532
rect 116676 571412 116728 571464
rect 120540 571412 120592 571464
rect 71780 571344 71832 571396
rect 74172 571344 74224 571396
rect 116584 571344 116636 571396
rect 117320 571344 117372 571396
rect 150348 571344 150400 571396
rect 151176 571344 151228 571396
rect 191104 571344 191156 571396
rect 195428 571344 195480 571396
rect 200120 570800 200172 570852
rect 239588 570800 239640 570852
rect 58808 570732 58860 570784
rect 91100 570732 91152 570784
rect 91560 570732 91612 570784
rect 96712 570732 96764 570784
rect 121460 570732 121512 570784
rect 211160 570732 211212 570784
rect 215300 570732 215352 570784
rect 301504 570732 301556 570784
rect 66352 570664 66404 570716
rect 120724 570664 120776 570716
rect 180800 570664 180852 570716
rect 301136 570664 301188 570716
rect 10324 570596 10376 570648
rect 321560 570596 321612 570648
rect 118700 569372 118752 569424
rect 154856 569372 154908 569424
rect 191840 569372 191892 569424
rect 238852 569372 238904 569424
rect 80060 569304 80112 569356
rect 120816 569304 120868 569356
rect 157432 569304 157484 569356
rect 213184 569304 213236 569356
rect 255320 569304 255372 569356
rect 324780 569304 324832 569356
rect 58532 569236 58584 569288
rect 110512 569236 110564 569288
rect 142804 569236 142856 569288
rect 213092 569236 213144 569288
rect 240140 569236 240192 569288
rect 309784 569236 309836 569288
rect 67732 569168 67784 569220
rect 123116 569168 123168 569220
rect 147404 569168 147456 569220
rect 165620 569168 165672 569220
rect 186320 569168 186372 569220
rect 301412 569168 301464 569220
rect 176660 568012 176712 568064
rect 235448 568012 235500 568064
rect 59452 567944 59504 567996
rect 75920 567944 75972 567996
rect 128360 567944 128412 567996
rect 211344 567944 211396 567996
rect 69112 567876 69164 567928
rect 114560 567876 114612 567928
rect 125692 567876 125744 567928
rect 211252 567876 211304 567928
rect 244464 567876 244516 567928
rect 318156 567876 318208 567928
rect 70400 567808 70452 567860
rect 121828 567808 121880 567860
rect 194600 567808 194652 567860
rect 302976 567808 303028 567860
rect 267740 567196 267792 567248
rect 321560 567196 321612 567248
rect 198740 566652 198792 566704
rect 239496 566652 239548 566704
rect 269212 566652 269264 566704
rect 311348 566652 311400 566704
rect 57244 566584 57296 566636
rect 89720 566584 89772 566636
rect 123024 566584 123076 566636
rect 211712 566584 211764 566636
rect 247040 566584 247092 566636
rect 324872 566584 324924 566636
rect 85580 566516 85632 566568
rect 121736 566516 121788 566568
rect 184940 566516 184992 566568
rect 294052 566516 294104 566568
rect 63592 566448 63644 566500
rect 122932 566448 122984 566500
rect 147036 566448 147088 566500
rect 168380 566448 168432 566500
rect 187700 566448 187752 566500
rect 302332 566448 302384 566500
rect 176752 565292 176804 565344
rect 244280 565292 244332 565344
rect 129832 565224 129884 565276
rect 212724 565224 212776 565276
rect 274640 565224 274692 565276
rect 316776 565224 316828 565276
rect 88524 565156 88576 565208
rect 104992 565156 105044 565208
rect 168472 565156 168524 565208
rect 210700 565156 210752 565208
rect 211160 565156 211212 565208
rect 301320 565156 301372 565208
rect 64972 565088 65024 565140
rect 123208 565088 123260 565140
rect 195980 565088 196032 565140
rect 302516 565088 302568 565140
rect 136732 563864 136784 563916
rect 210792 563864 210844 563916
rect 263600 563864 263652 563916
rect 307024 563864 307076 563916
rect 81440 563796 81492 563848
rect 89812 563796 89864 563848
rect 152004 563796 152056 563848
rect 213000 563796 213052 563848
rect 273260 563796 273312 563848
rect 322388 563796 322440 563848
rect 59544 563728 59596 563780
rect 100760 563728 100812 563780
rect 210056 563728 210108 563780
rect 302700 563728 302752 563780
rect 78772 563660 78824 563712
rect 123484 563660 123536 563712
rect 186412 563660 186464 563712
rect 302424 563660 302476 563712
rect 204352 562436 204404 562488
rect 239404 562436 239456 562488
rect 146944 562368 146996 562420
rect 212540 562368 212592 562420
rect 58992 562300 59044 562352
rect 102232 562300 102284 562352
rect 189080 562300 189132 562352
rect 288624 562300 288676 562352
rect 4804 561688 4856 561740
rect 321560 561688 321612 561740
rect 178040 561144 178092 561196
rect 233884 561144 233936 561196
rect 73252 561076 73304 561128
rect 107660 561076 107712 561128
rect 187792 561076 187844 561128
rect 253940 561076 253992 561128
rect 256792 561076 256844 561128
rect 323952 561076 324004 561128
rect 80152 561008 80204 561060
rect 121092 561008 121144 561060
rect 138020 561008 138072 561060
rect 211620 561008 211672 561060
rect 249800 561008 249852 561060
rect 323860 561008 323912 561060
rect 59268 560940 59320 560992
rect 117320 560940 117372 560992
rect 147220 560940 147272 560992
rect 173992 560940 174044 560992
rect 200212 560940 200264 560992
rect 302792 560940 302844 560992
rect 207020 559716 207072 559768
rect 220176 559716 220228 559768
rect 197360 559648 197412 559700
rect 214748 559648 214800 559700
rect 259460 559648 259512 559700
rect 305736 559648 305788 559700
rect 88432 559580 88484 559632
rect 103520 559580 103572 559632
rect 127072 559580 127124 559632
rect 204260 559580 204312 559632
rect 216772 559580 216824 559632
rect 273904 559580 273956 559632
rect 59176 559512 59228 559564
rect 107660 559512 107712 559564
rect 182180 559512 182232 559564
rect 300676 559512 300728 559564
rect 40040 558832 40092 558884
rect 321560 558832 321612 558884
rect 281540 558288 281592 558340
rect 304264 558288 304316 558340
rect 190460 558220 190512 558272
rect 222844 558220 222896 558272
rect 242900 558220 242952 558272
rect 320916 558220 320968 558272
rect 67824 558152 67876 558204
rect 107752 558152 107804 558204
rect 133144 558152 133196 558204
rect 198832 558152 198884 558204
rect 205640 558152 205692 558204
rect 285680 558152 285732 558204
rect 199200 556996 199252 557048
rect 216128 556996 216180 557048
rect 76012 556928 76064 556980
rect 86776 556928 86828 556980
rect 206376 556928 206428 556980
rect 262220 556928 262272 556980
rect 266544 556928 266596 556980
rect 322296 556928 322348 556980
rect 62212 556860 62264 556912
rect 109684 556860 109736 556912
rect 124680 556860 124732 556912
rect 210976 556860 211028 556912
rect 250076 556860 250128 556912
rect 314200 556860 314252 556912
rect 71688 556792 71740 556844
rect 121644 556792 121696 556844
rect 179144 556792 179196 556844
rect 291292 556792 291344 556844
rect 215760 556180 215812 556232
rect 217416 556180 217468 556232
rect 125600 556044 125652 556096
rect 126888 556044 126940 556096
rect 193496 555704 193548 555756
rect 232504 555704 232556 555756
rect 154120 555636 154172 555688
rect 212908 555636 212960 555688
rect 121092 555568 121144 555620
rect 198004 555568 198056 555620
rect 251548 555568 251600 555620
rect 323768 555568 323820 555620
rect 71044 555500 71096 555552
rect 105360 555500 105412 555552
rect 191380 555500 191432 555552
rect 277400 555500 277452 555552
rect 279516 555500 279568 555552
rect 313924 555500 313976 555552
rect 57612 555432 57664 555484
rect 77208 555432 77260 555484
rect 82452 555432 82504 555484
rect 116676 555432 116728 555484
rect 148692 555432 148744 555484
rect 160560 555432 160612 555484
rect 198556 555432 198608 555484
rect 287704 555432 287756 555484
rect 259460 554208 259512 554260
rect 320824 554208 320876 554260
rect 184940 554140 184992 554192
rect 235356 554140 235408 554192
rect 253664 554140 253716 554192
rect 323676 554140 323728 554192
rect 76748 554072 76800 554124
rect 116584 554072 116636 554124
rect 148416 554072 148468 554124
rect 172520 554072 172572 554124
rect 192760 554072 192812 554124
rect 280804 554072 280856 554124
rect 63132 554004 63184 554056
rect 110604 554004 110656 554056
rect 140504 554004 140556 554056
rect 193864 554004 193916 554056
rect 197084 554004 197136 554056
rect 302608 554004 302660 554056
rect 290924 552916 290976 552968
rect 295340 552916 295392 552968
rect 145012 552848 145064 552900
rect 146208 552848 146260 552900
rect 107752 552780 107804 552832
rect 108948 552780 109000 552832
rect 64972 552712 65024 552764
rect 65984 552712 66036 552764
rect 67640 552712 67692 552764
rect 68836 552712 68888 552764
rect 69020 552712 69072 552764
rect 70308 552712 70360 552764
rect 78680 552712 78732 552764
rect 79600 552712 79652 552764
rect 89720 552712 89772 552764
rect 91008 552712 91060 552764
rect 94596 552712 94648 552764
rect 123300 552780 123352 552832
rect 171324 552780 171376 552832
rect 210884 552780 210936 552832
rect 211160 552780 211212 552832
rect 212172 552780 212224 552832
rect 213552 552780 213604 552832
rect 235264 552848 235316 552900
rect 283748 552848 283800 552900
rect 309876 552848 309928 552900
rect 222200 552780 222252 552832
rect 222844 552780 222896 552832
rect 227720 552780 227772 552832
rect 228640 552780 228692 552832
rect 124220 552712 124272 552764
rect 125416 552712 125468 552764
rect 126980 552712 127032 552764
rect 128268 552712 128320 552764
rect 129740 552712 129792 552764
rect 130476 552712 130528 552764
rect 136640 552712 136692 552764
rect 137652 552712 137704 552764
rect 140780 552712 140832 552764
rect 141884 552712 141936 552764
rect 142160 552712 142212 552764
rect 143356 552712 143408 552764
rect 143540 552712 143592 552764
rect 144736 552712 144788 552764
rect 147680 552712 147732 552764
rect 191104 552712 191156 552764
rect 198740 552712 198792 552764
rect 199936 552712 199988 552764
rect 200120 552712 200172 552764
rect 201408 552712 201460 552764
rect 208584 552712 208636 552764
rect 238300 552780 238352 552832
rect 255320 552780 255372 552832
rect 256516 552780 256568 552832
rect 256792 552780 256844 552832
rect 257988 552780 258040 552832
rect 267280 552780 267332 552832
rect 311164 552780 311216 552832
rect 231860 552712 231912 552764
rect 232872 552712 232924 552764
rect 233240 552712 233292 552764
rect 234344 552712 234396 552764
rect 246488 552712 246540 552764
rect 311256 552712 311308 552764
rect 57704 552644 57756 552696
rect 103244 552644 103296 552696
rect 104900 552644 104952 552696
rect 106096 552644 106148 552696
rect 106280 552644 106332 552696
rect 107568 552644 107620 552696
rect 121460 552644 121512 552696
rect 122564 552644 122616 552696
rect 122840 552644 122892 552696
rect 124036 552644 124088 552696
rect 151176 552644 151228 552696
rect 163412 552644 163464 552696
rect 168380 552644 168432 552696
rect 169116 552644 169168 552696
rect 179420 552644 179472 552696
rect 180616 552644 180668 552696
rect 180800 552644 180852 552696
rect 181996 552644 182048 552696
rect 181352 552576 181404 552628
rect 301228 552644 301280 552696
rect 219440 552576 219492 552628
rect 220728 552576 220780 552628
rect 273260 552576 273312 552628
rect 274456 552576 274508 552628
rect 291200 552576 291252 552628
rect 292396 552576 292448 552628
rect 293960 552576 294012 552628
rect 295248 552576 295300 552628
rect 295340 552576 295392 552628
rect 322480 552576 322532 552628
rect 286692 552508 286744 552560
rect 319536 552508 319588 552560
rect 285680 552440 285732 552492
rect 321008 552440 321060 552492
rect 285956 552372 286008 552424
rect 322664 552372 322716 552424
rect 285220 552304 285272 552356
rect 322296 552304 322348 552356
rect 258724 552236 258776 552288
rect 321100 552236 321152 552288
rect 252284 552168 252336 552220
rect 321560 552168 321612 552220
rect 241612 552100 241664 552152
rect 320916 552100 320968 552152
rect 237932 552032 237984 552084
rect 320824 552032 320876 552084
rect 113272 551964 113324 552016
rect 121920 551964 121972 552016
rect 148508 551964 148560 552016
rect 149060 551964 149112 552016
rect 211436 551964 211488 552016
rect 214656 551964 214708 552016
rect 207112 551488 207164 551540
rect 229744 551488 229796 551540
rect 244372 551488 244424 551540
rect 304264 551488 304316 551540
rect 189908 551420 189960 551472
rect 238116 551420 238168 551472
rect 249432 551420 249484 551472
rect 321192 551420 321244 551472
rect 147496 551352 147548 551404
rect 167000 551352 167052 551404
rect 202788 551352 202840 551404
rect 256700 551352 256752 551404
rect 86224 551284 86276 551336
rect 114652 551284 114704 551336
rect 120448 551284 120500 551336
rect 130384 551284 130436 551336
rect 142620 551284 142672 551336
rect 211528 551284 211580 551336
rect 271604 551284 271656 551336
rect 312544 551284 312596 551336
rect 262312 551216 262364 551268
rect 300124 551216 300176 551268
rect 264428 551148 264480 551200
rect 302884 551148 302936 551200
rect 254400 551080 254452 551132
rect 302976 551080 303028 551132
rect 273720 551012 273772 551064
rect 322572 551012 322624 551064
rect 272340 550944 272392 550996
rect 323676 550944 323728 550996
rect 273076 550876 273128 550928
rect 324780 550876 324832 550928
rect 265900 550808 265952 550860
rect 324688 550808 324740 550860
rect 135444 550740 135496 550792
rect 144184 550740 144236 550792
rect 287336 550740 287388 550792
rect 322388 550740 322440 550792
rect 164332 550672 164384 550724
rect 165528 550672 165580 550724
rect 255872 550672 255924 550724
rect 324872 550672 324924 550724
rect 291660 550604 291712 550656
rect 319444 550604 319496 550656
rect 61660 550536 61712 550588
rect 62764 550536 62816 550588
rect 79324 550536 79376 550588
rect 81716 550536 81768 550588
rect 108304 550536 108356 550588
rect 111800 550536 111852 550588
rect 115480 550536 115532 550588
rect 116124 550536 116176 550588
rect 136180 550536 136232 550588
rect 140044 550536 140096 550588
rect 144092 550536 144144 550588
rect 146852 550536 146904 550588
rect 146944 550536 146996 550588
rect 148324 550536 148376 550588
rect 149888 550536 149940 550588
rect 151268 550536 151320 550588
rect 219992 550536 220044 550588
rect 228364 550536 228416 550588
rect 230020 550536 230072 550588
rect 231124 550536 231176 550588
rect 235080 550536 235132 550588
rect 236644 550536 236696 550588
rect 55128 550468 55180 550520
rect 67364 550468 67416 550520
rect 209228 550468 209280 550520
rect 216036 550468 216088 550520
rect 118240 550400 118292 550452
rect 126244 550400 126296 550452
rect 209964 550400 210016 550452
rect 220084 550400 220136 550452
rect 54944 550332 54996 550384
rect 88892 550332 88944 550384
rect 118976 550332 119028 550384
rect 129096 550332 129148 550384
rect 203524 550332 203576 550384
rect 214564 550332 214616 550384
rect 225052 550332 225104 550384
rect 235540 550332 235592 550384
rect 57796 550264 57848 550316
rect 93216 550264 93268 550316
rect 114008 550264 114060 550316
rect 124404 550264 124456 550316
rect 151084 550264 151136 550316
rect 153384 550264 153436 550316
rect 157340 550264 157392 550316
rect 167092 550264 167144 550316
rect 204260 550264 204312 550316
rect 217324 550264 217376 550316
rect 230756 550264 230808 550316
rect 246304 550264 246356 550316
rect 56508 550196 56560 550248
rect 83924 550196 83976 550248
rect 85304 550196 85356 550248
rect 120908 550196 120960 550248
rect 195612 550196 195664 550248
rect 215944 550196 215996 550248
rect 225788 550196 225840 550248
rect 241520 550196 241572 550248
rect 295984 550196 296036 550248
rect 300676 550196 300728 550248
rect 58624 550128 58676 550180
rect 95332 550128 95384 550180
rect 96068 550128 96120 550180
rect 119344 550128 119396 550180
rect 147588 550128 147640 550180
rect 157708 550128 157760 550180
rect 160192 550128 160244 550180
rect 172704 550128 172756 550180
rect 215024 550128 215076 550180
rect 236736 550128 236788 550180
rect 242256 550128 242308 550180
rect 303160 550128 303212 550180
rect 55036 550060 55088 550112
rect 98920 550060 98972 550112
rect 106832 550060 106884 550112
rect 124312 550060 124364 550112
rect 146116 550060 146168 550112
rect 156972 550060 157024 550112
rect 170588 550060 170640 550112
rect 195244 550060 195296 550112
rect 212816 550060 212868 550112
rect 249064 550060 249116 550112
rect 270868 550060 270920 550112
rect 322756 550060 322808 550112
rect 56416 549992 56468 550044
rect 73804 549992 73856 550044
rect 78128 549992 78180 550044
rect 121552 549992 121604 550044
rect 152004 549992 152056 550044
rect 56324 549924 56376 549976
rect 99656 549924 99708 549976
rect 103980 549924 104032 549976
rect 125784 549924 125836 549976
rect 148968 549924 149020 549976
rect 167000 549992 167052 550044
rect 175556 549992 175608 550044
rect 183468 549992 183520 550044
rect 231216 549992 231268 550044
rect 252928 549992 252980 550044
rect 321284 549992 321336 550044
rect 60372 549856 60424 549908
rect 116860 549856 116912 549908
rect 121828 549856 121880 549908
rect 167736 549924 167788 549976
rect 176292 549924 176344 549976
rect 238208 549924 238260 549976
rect 299572 549924 299624 549976
rect 316684 549924 316736 549976
rect 171968 549856 172020 549908
rect 169760 549720 169812 549772
rect 173440 549720 173492 549772
rect 192484 549856 192536 549908
rect 194232 549856 194284 549908
rect 226984 549856 227036 549908
rect 237196 549856 237248 549908
rect 285680 549856 285732 549908
rect 298836 549856 298888 549908
rect 323584 549856 323636 549908
rect 283104 549788 283156 549840
rect 301872 549788 301924 549840
rect 280160 549720 280212 549772
rect 300308 549720 300360 549772
rect 275928 549652 275980 549704
rect 300216 549652 300268 549704
rect 277308 549584 277360 549636
rect 305736 549584 305788 549636
rect 257252 549516 257304 549568
rect 301596 549516 301648 549568
rect 240048 549448 240100 549500
rect 273260 549448 273312 549500
rect 278044 549448 278096 549500
rect 324136 549448 324188 549500
rect 138296 549380 138348 549432
rect 142804 549380 142856 549432
rect 284484 549380 284536 549432
rect 300492 549380 300544 549432
rect 296720 549312 296772 549364
rect 323768 549312 323820 549364
rect 131212 549244 131264 549296
rect 133144 549244 133196 549296
rect 281632 549244 281684 549296
rect 300584 549244 300636 549296
rect 293776 548768 293828 548820
rect 322848 548768 322900 548820
rect 268752 548700 268804 548752
rect 303068 548700 303120 548752
rect 265164 548632 265216 548684
rect 307024 548632 307076 548684
rect 278780 548564 278832 548616
rect 321560 548564 321612 548616
rect 273260 548496 273312 548548
rect 322112 548496 322164 548548
rect 276572 548428 276624 548480
rect 324596 548428 324648 548480
rect 247224 548360 247276 548412
rect 301780 548360 301832 548412
rect 243636 548292 243688 548344
rect 301964 548292 302016 548344
rect 263048 548224 263100 548276
rect 324504 548224 324556 548276
rect 260840 548156 260892 548208
rect 323860 548156 323912 548208
rect 235816 548088 235868 548140
rect 236460 548088 236512 548140
rect 301044 548088 301096 548140
rect 323584 548020 323636 548072
rect 301044 543668 301096 543720
rect 321560 543668 321612 543720
rect 302792 539588 302844 539640
rect 311164 539588 311216 539640
rect 301964 539520 302016 539572
rect 321560 539520 321612 539572
rect 324688 533400 324740 533452
rect 324780 533196 324832 533248
rect 300676 529864 300728 529916
rect 457444 529864 457496 529916
rect 300584 529796 300636 529848
rect 436468 529796 436520 529848
rect 300492 529728 300544 529780
rect 436192 529728 436244 529780
rect 301872 529660 301924 529712
rect 436100 529660 436152 529712
rect 303160 529592 303212 529644
rect 436560 529592 436612 529644
rect 305736 529524 305788 529576
rect 436376 529524 436428 529576
rect 322756 529456 322808 529508
rect 436284 529456 436336 529508
rect 319536 528504 319588 528556
rect 512184 528504 512236 528556
rect 322664 528436 322716 528488
rect 495440 528436 495492 528488
rect 322480 528368 322532 528420
rect 488540 528368 488592 528420
rect 322848 528300 322900 528352
rect 465080 528300 465132 528352
rect 323768 528232 323820 528284
rect 459560 528232 459612 528284
rect 300308 528164 300360 528216
rect 436928 528164 436980 528216
rect 301596 528096 301648 528148
rect 436836 528096 436888 528148
rect 321284 528028 321336 528080
rect 436652 528028 436704 528080
rect 324136 527960 324188 528012
rect 436744 527960 436796 528012
rect 305644 527892 305696 527944
rect 374276 527892 374328 527944
rect 300216 527824 300268 527876
rect 356244 527824 356296 527876
rect 307024 527076 307076 527128
rect 324964 527144 325016 527196
rect 324596 527076 324648 527128
rect 420000 527076 420052 527128
rect 323860 527008 323912 527060
rect 347228 527008 347280 527060
rect 323584 526940 323636 526992
rect 338212 526940 338264 526992
rect 324872 526872 324924 526924
rect 411260 526872 411312 526924
rect 324504 526804 324556 526856
rect 406476 526804 406528 526856
rect 322572 526736 322624 526788
rect 401968 526736 402020 526788
rect 302884 526668 302936 526720
rect 379520 526668 379572 526720
rect 324780 526600 324832 526652
rect 388444 526600 388496 526652
rect 301780 526532 301832 526584
rect 365260 526532 365312 526584
rect 302976 526464 303028 526516
rect 351920 526464 351972 526516
rect 324688 526396 324740 526448
rect 369860 526396 369912 526448
rect 323676 526328 323728 526380
rect 415584 526328 415636 526380
rect 303068 526260 303120 526312
rect 393320 526260 393372 526312
rect 300124 526192 300176 526244
rect 333980 526192 334032 526244
rect 301504 525716 301556 525768
rect 512276 525716 512328 525768
rect 322388 525648 322440 525700
rect 476120 525648 476172 525700
rect 322296 525580 322348 525632
rect 470600 525580 470652 525632
rect 321100 525512 321152 525564
rect 433340 525512 433392 525564
rect 302884 524424 302936 524476
rect 519544 524424 519596 524476
rect 319444 524356 319496 524408
rect 457628 524356 457680 524408
rect 321008 524288 321060 524340
rect 434628 524288 434680 524340
rect 320824 524220 320876 524272
rect 433524 524220 433576 524272
rect 320916 524152 320968 524204
rect 433432 524152 433484 524204
rect 329748 524084 329800 524136
rect 434720 524084 434772 524136
rect 53748 517488 53800 517540
rect 57888 517488 57940 517540
rect 311164 515380 311216 515432
rect 580264 515380 580316 515432
rect 560944 511912 560996 511964
rect 580172 511912 580224 511964
rect 302240 495456 302292 495508
rect 520924 495456 520976 495508
rect 274656 487772 274708 487824
rect 274824 487772 274876 487824
rect 64880 487024 64932 487076
rect 65156 487024 65208 487076
rect 128360 487024 128412 487076
rect 128636 487024 128688 487076
rect 207112 487024 207164 487076
rect 207388 487024 207440 487076
rect 140872 486684 140924 486736
rect 199108 486684 199160 486736
rect 121184 486616 121236 486668
rect 197912 486616 197964 486668
rect 109408 486548 109460 486600
rect 198372 486548 198424 486600
rect 109500 486480 109552 486532
rect 204812 486480 204864 486532
rect 15844 486412 15896 486464
rect 383660 486412 383712 486464
rect 73988 485732 74040 485784
rect 105084 485732 105136 485784
rect 107844 485732 107896 485784
rect 108028 485732 108080 485784
rect 151268 485732 151320 485784
rect 204904 485732 204956 485784
rect 60004 485664 60056 485716
rect 91836 485664 91888 485716
rect 149520 485664 149572 485716
rect 201316 485664 201368 485716
rect 201408 485664 201460 485716
rect 212080 485732 212132 485784
rect 262404 485732 262456 485784
rect 262588 485732 262640 485784
rect 285772 485732 285824 485784
rect 285956 485732 286008 485784
rect 234528 485664 234580 485716
rect 56508 485596 56560 485648
rect 89628 485596 89680 485648
rect 154304 485596 154356 485648
rect 212540 485596 212592 485648
rect 59084 485528 59136 485580
rect 92296 485528 92348 485580
rect 162124 485528 162176 485580
rect 244556 485664 244608 485716
rect 356796 485664 356848 485716
rect 239680 485596 239732 485648
rect 358268 485596 358320 485648
rect 64144 485460 64196 485512
rect 72424 485460 72476 485512
rect 79324 485460 79376 485512
rect 106372 485460 106424 485512
rect 152188 485460 152240 485512
rect 204260 485460 204312 485512
rect 55128 485392 55180 485444
rect 88340 485392 88392 485444
rect 149428 485392 149480 485444
rect 200488 485392 200540 485444
rect 201316 485392 201368 485444
rect 208492 485392 208544 485444
rect 364984 485528 365036 485580
rect 211068 485460 211120 485512
rect 217416 485460 217468 485512
rect 226064 485460 226116 485512
rect 356704 485460 356756 485512
rect 211160 485392 211212 485444
rect 230848 485392 230900 485444
rect 362224 485392 362276 485444
rect 56416 485324 56468 485376
rect 90548 485324 90600 485376
rect 148232 485324 148284 485376
rect 197452 485324 197504 485376
rect 209688 485324 209740 485376
rect 221740 485324 221792 485376
rect 225604 485324 225656 485376
rect 358176 485324 358228 485376
rect 50988 485256 51040 485308
rect 93584 485256 93636 485308
rect 156696 485256 156748 485308
rect 162124 485256 162176 485308
rect 162216 485256 162268 485308
rect 205640 485256 205692 485308
rect 240048 485256 240100 485308
rect 373264 485256 373316 485308
rect 51816 485188 51868 485240
rect 99380 485188 99432 485240
rect 150440 485188 150492 485240
rect 42432 485120 42484 485172
rect 102876 485120 102928 485172
rect 161480 485120 161532 485172
rect 43628 485052 43680 485104
rect 104624 485052 104676 485104
rect 110328 485052 110380 485104
rect 170404 485052 170456 485104
rect 197360 485120 197412 485172
rect 201500 485188 201552 485240
rect 199384 485120 199436 485172
rect 209780 485188 209832 485240
rect 209872 485188 209924 485240
rect 219900 485188 219952 485240
rect 224040 485188 224092 485240
rect 360844 485188 360896 485240
rect 206836 485120 206888 485172
rect 219164 485120 219216 485172
rect 231768 485120 231820 485172
rect 369124 485120 369176 485172
rect 200212 485052 200264 485104
rect 217416 485052 217468 485104
rect 223488 485052 223540 485104
rect 371884 485052 371936 485104
rect 52184 484984 52236 485036
rect 81716 484984 81768 485036
rect 157432 484984 157484 485036
rect 162216 484984 162268 485036
rect 50620 484916 50672 484968
rect 73252 484916 73304 484968
rect 73804 484916 73856 484968
rect 79324 484916 79376 484968
rect 139400 484916 139452 484968
rect 73896 484848 73948 484900
rect 95332 484848 95384 484900
rect 50896 484780 50948 484832
rect 73344 484780 73396 484832
rect 68284 484712 68336 484764
rect 84384 484712 84436 484764
rect 158720 484916 158772 484968
rect 204260 484984 204312 485036
rect 209780 484984 209832 485036
rect 214748 484984 214800 485036
rect 155592 484848 155644 484900
rect 161480 484848 161532 484900
rect 185584 484916 185636 484968
rect 195336 484916 195388 484968
rect 211620 484916 211672 484968
rect 166264 484780 166316 484832
rect 203524 484848 203576 484900
rect 204904 484780 204956 484832
rect 211160 484780 211212 484832
rect 212540 484440 212592 484492
rect 212724 484440 212776 484492
rect 195152 484372 195204 484424
rect 197084 484372 197136 484424
rect 201960 484372 202012 484424
rect 203984 484372 204036 484424
rect 211896 484372 211948 484424
rect 212908 484372 212960 484424
rect 213368 484372 213420 484424
rect 216220 484372 216272 484424
rect 216588 484372 216640 484424
rect 219164 484372 219216 484424
rect 219992 484372 220044 484424
rect 222660 484372 222712 484424
rect 129832 484304 129884 484356
rect 130016 484304 130068 484356
rect 129740 484236 129792 484288
rect 129924 484236 129976 484288
rect 281632 484236 281684 484288
rect 70492 484168 70544 484220
rect 71228 484168 71280 484220
rect 78680 484168 78732 484220
rect 79140 484168 79192 484220
rect 172520 484168 172572 484220
rect 173532 484168 173584 484220
rect 191840 484168 191892 484220
rect 192392 484168 192444 484220
rect 193220 484168 193272 484220
rect 194140 484168 194192 484220
rect 198740 484168 198792 484220
rect 199476 484168 199528 484220
rect 205732 484168 205784 484220
rect 206468 484168 206520 484220
rect 219532 484168 219584 484220
rect 220084 484168 220136 484220
rect 70400 484100 70452 484152
rect 70860 484100 70912 484152
rect 71872 484100 71924 484152
rect 72608 484100 72660 484152
rect 74632 484100 74684 484152
rect 75276 484100 75328 484152
rect 75920 484100 75972 484152
rect 76564 484100 76616 484152
rect 78772 484100 78824 484152
rect 79692 484100 79744 484152
rect 93860 484100 93912 484152
rect 94596 484100 94648 484152
rect 131120 484100 131172 484152
rect 132132 484100 132184 484152
rect 132592 484100 132644 484152
rect 133420 484100 133472 484152
rect 133880 484100 133932 484152
rect 134708 484100 134760 484152
rect 139400 484100 139452 484152
rect 140044 484100 140096 484152
rect 140872 484100 140924 484152
rect 141332 484100 141384 484152
rect 142160 484100 142212 484152
rect 142620 484100 142672 484152
rect 143540 484100 143592 484152
rect 144460 484100 144512 484152
rect 147680 484100 147732 484152
rect 148324 484100 148376 484152
rect 167092 484100 167144 484152
rect 167736 484100 167788 484152
rect 171140 484100 171192 484152
rect 171692 484100 171744 484152
rect 172612 484100 172664 484152
rect 172980 484100 173032 484152
rect 175280 484100 175332 484152
rect 175740 484100 175792 484152
rect 186320 484100 186372 484152
rect 187148 484100 187200 484152
rect 187792 484100 187844 484152
rect 188436 484100 188488 484152
rect 190460 484100 190512 484152
rect 191012 484100 191064 484152
rect 191932 484100 191984 484152
rect 192116 484100 192168 484152
rect 193312 484100 193364 484152
rect 193772 484100 193824 484152
rect 197452 484100 197504 484152
rect 198188 484100 198240 484152
rect 201592 484100 201644 484152
rect 202052 484100 202104 484152
rect 204444 484100 204496 484152
rect 205180 484100 205232 484152
rect 205640 484100 205692 484152
rect 206100 484100 206152 484152
rect 207020 484100 207072 484152
rect 207756 484100 207808 484152
rect 208492 484100 208544 484152
rect 209136 484100 209188 484152
rect 209780 484100 209832 484152
rect 210516 484100 210568 484152
rect 212632 484100 212684 484152
rect 213460 484100 213512 484152
rect 213920 484100 213972 484152
rect 214932 484100 214984 484152
rect 216772 484100 216824 484152
rect 217508 484100 217560 484152
rect 219440 484100 219492 484152
rect 219716 484100 219768 484152
rect 223580 484100 223632 484152
rect 224132 484100 224184 484152
rect 226340 484100 226392 484152
rect 226708 484100 226760 484152
rect 229100 484100 229152 484152
rect 229468 484100 229520 484152
rect 240232 484100 240284 484152
rect 240876 484100 240928 484152
rect 241520 484100 241572 484152
rect 242164 484100 242216 484152
rect 263692 484100 263744 484152
rect 264244 484100 264296 484152
rect 264980 484100 265032 484152
rect 265532 484100 265584 484152
rect 269120 484100 269172 484152
rect 269948 484100 270000 484152
rect 270500 484100 270552 484152
rect 270868 484100 270920 484152
rect 271972 484100 272024 484152
rect 272524 484100 272576 484152
rect 273352 484100 273404 484152
rect 273812 484100 273864 484152
rect 293960 484100 294012 484152
rect 371700 484100 371752 484152
rect 359464 484032 359516 484084
rect 129832 483964 129884 484016
rect 130292 483964 130344 484016
rect 202972 483964 203024 484016
rect 203892 483964 203944 484016
rect 226432 483964 226484 484016
rect 227260 483964 227312 484016
rect 280068 483964 280120 484016
rect 362776 483964 362828 484016
rect 279792 483896 279844 483948
rect 372344 483896 372396 483948
rect 275560 483828 275612 483880
rect 370412 483828 370464 483880
rect 176568 483760 176620 483812
rect 206376 483760 206428 483812
rect 260104 483760 260156 483812
rect 370688 483760 370740 483812
rect 165528 483692 165580 483744
rect 214564 483692 214616 483744
rect 236736 483692 236788 483744
rect 362316 483692 362368 483744
rect 60648 483624 60700 483676
rect 80704 483624 80756 483676
rect 161572 483624 161624 483676
rect 215944 483624 215996 483676
rect 246948 483624 247000 483676
rect 378784 483624 378836 483676
rect 189080 483352 189132 483404
rect 189356 483352 189408 483404
rect 50436 482944 50488 482996
rect 97172 482944 97224 482996
rect 48044 482876 48096 482928
rect 97540 482876 97592 482928
rect 290096 482876 290148 482928
rect 367008 482876 367060 482928
rect 49240 482808 49292 482860
rect 98000 482808 98052 482860
rect 203708 482808 203760 482860
rect 209412 482808 209464 482860
rect 274824 482808 274876 482860
rect 365536 482808 365588 482860
rect 47860 482740 47912 482792
rect 111708 482740 111760 482792
rect 271788 482740 271840 482792
rect 366916 482740 366968 482792
rect 46572 482672 46624 482724
rect 111248 482672 111300 482724
rect 159272 482672 159324 482724
rect 207756 482672 207808 482724
rect 276664 482672 276716 482724
rect 374460 482672 374512 482724
rect 50528 482604 50580 482656
rect 115664 482604 115716 482656
rect 135628 482604 135680 482656
rect 141792 482604 141844 482656
rect 160560 482604 160612 482656
rect 211804 482604 211856 482656
rect 276848 482604 276900 482656
rect 375840 482604 375892 482656
rect 46388 482536 46440 482588
rect 112536 482536 112588 482588
rect 138480 482536 138532 482588
rect 200304 482536 200356 482588
rect 261392 482536 261444 482588
rect 368020 482536 368072 482588
rect 46480 482468 46532 482520
rect 112076 482468 112128 482520
rect 136824 482468 136876 482520
rect 199108 482468 199160 482520
rect 257528 482468 257580 482520
rect 366640 482468 366692 482520
rect 49148 482400 49200 482452
rect 115204 482400 115256 482452
rect 140780 482400 140832 482452
rect 141700 482400 141752 482452
rect 141792 482400 141844 482452
rect 198004 482400 198056 482452
rect 244648 482400 244700 482452
rect 373356 482400 373408 482452
rect 48136 482332 48188 482384
rect 119620 482332 119672 482384
rect 137928 482332 137980 482384
rect 201868 482332 201920 482384
rect 248328 482332 248380 482384
rect 378968 482332 379020 482384
rect 46664 482264 46716 482316
rect 120080 482264 120132 482316
rect 138572 482264 138624 482316
rect 207296 482264 207348 482316
rect 222568 482264 222620 482316
rect 376024 482264 376076 482316
rect 51908 482196 51960 482248
rect 98460 482196 98512 482248
rect 54852 482128 54904 482180
rect 96712 482128 96764 482180
rect 58716 482060 58768 482112
rect 96252 482060 96304 482112
rect 189172 481720 189224 481772
rect 189724 481720 189776 481772
rect 291292 481448 291344 481500
rect 291476 481448 291528 481500
rect 295524 481448 295576 481500
rect 295708 481448 295760 481500
rect 285496 481380 285548 481432
rect 359740 481380 359792 481432
rect 281448 481312 281500 481364
rect 357072 481312 357124 481364
rect 269028 481244 269080 481296
rect 361396 481244 361448 481296
rect 261208 481176 261260 481228
rect 358360 481176 358412 481228
rect 251364 481108 251416 481160
rect 251548 481108 251600 481160
rect 269304 481108 269356 481160
rect 377496 481108 377548 481160
rect 67732 481040 67784 481092
rect 67916 481040 67968 481092
rect 179604 481040 179656 481092
rect 179788 481040 179840 481092
rect 182364 481040 182416 481092
rect 182548 481040 182600 481092
rect 243084 481040 243136 481092
rect 370504 481040 370556 481092
rect 57888 480972 57940 481024
rect 114284 480972 114336 481024
rect 159088 480972 159140 481024
rect 209044 480972 209096 481024
rect 248052 480972 248104 481024
rect 376116 480972 376168 481024
rect 3792 480904 3844 480956
rect 434812 480904 434864 480956
rect 62120 480836 62172 480888
rect 62948 480836 63000 480888
rect 69112 480836 69164 480888
rect 69940 480836 69992 480888
rect 81532 480836 81584 480888
rect 82268 480836 82320 480888
rect 82820 480836 82872 480888
rect 83556 480836 83608 480888
rect 84292 480836 84344 480888
rect 84936 480836 84988 480888
rect 85580 480836 85632 480888
rect 86316 480836 86368 480888
rect 99472 480836 99524 480888
rect 100300 480836 100352 480888
rect 100760 480836 100812 480888
rect 101588 480836 101640 480888
rect 106372 480836 106424 480888
rect 106924 480836 106976 480888
rect 113272 480836 113324 480888
rect 113548 480836 113600 480888
rect 125600 480836 125652 480888
rect 126336 480836 126388 480888
rect 161480 480836 161532 480888
rect 161940 480836 161992 480888
rect 176660 480836 176712 480888
rect 177396 480836 177448 480888
rect 180800 480836 180852 480888
rect 181444 480836 181496 480888
rect 182180 480836 182232 480888
rect 182732 480836 182784 480888
rect 183560 480836 183612 480888
rect 184388 480836 184440 480888
rect 248420 480836 248472 480888
rect 248788 480836 248840 480888
rect 249800 480836 249852 480888
rect 250536 480836 250588 480888
rect 251180 480836 251232 480888
rect 251916 480836 251968 480888
rect 252560 480836 252612 480888
rect 253204 480836 253256 480888
rect 258080 480836 258132 480888
rect 258540 480836 258592 480888
rect 262312 480836 262364 480888
rect 262864 480836 262916 480888
rect 282920 480836 282972 480888
rect 283564 480836 283616 480888
rect 284300 480836 284352 480888
rect 284484 480836 284536 480888
rect 287060 480836 287112 480888
rect 287980 480836 288032 480888
rect 289820 480836 289872 480888
rect 290556 480836 290608 480888
rect 293960 480836 294012 480888
rect 294604 480836 294656 480888
rect 295340 480836 295392 480888
rect 295892 480836 295944 480888
rect 296720 480836 296772 480888
rect 297180 480836 297232 480888
rect 179512 480700 179564 480752
rect 180064 480700 180116 480752
rect 220820 480224 220872 480276
rect 221004 480224 221056 480276
rect 57244 480156 57296 480208
rect 123024 480156 123076 480208
rect 46756 480088 46808 480140
rect 116216 480088 116268 480140
rect 293316 480088 293368 480140
rect 370320 480088 370372 480140
rect 48228 480020 48280 480072
rect 117504 480020 117556 480072
rect 299480 480020 299532 480072
rect 379244 480020 379296 480072
rect 59728 479952 59780 480004
rect 129832 479952 129884 480004
rect 278780 479952 278832 480004
rect 365628 479952 365680 480004
rect 45468 479884 45520 479936
rect 117596 479884 117648 479936
rect 256332 479884 256384 479936
rect 356888 479884 356940 479936
rect 43720 479816 43772 479868
rect 117964 479816 118016 479868
rect 265900 479816 265952 479868
rect 366732 479816 366784 479868
rect 47676 479748 47728 479800
rect 129740 479748 129792 479800
rect 259552 479748 259604 479800
rect 365352 479748 365404 479800
rect 47768 479680 47820 479732
rect 129924 479680 129976 479732
rect 254492 479680 254544 479732
rect 369492 479680 369544 479732
rect 46112 479612 46164 479664
rect 128912 479612 128964 479664
rect 189264 479612 189316 479664
rect 200764 479612 200816 479664
rect 243452 479612 243504 479664
rect 360936 479612 360988 479664
rect 47584 479544 47636 479596
rect 134340 479544 134392 479596
rect 160192 479544 160244 479596
rect 210516 479544 210568 479596
rect 246120 479544 246172 479596
rect 369216 479544 369268 479596
rect 62396 479476 62448 479528
rect 199292 479476 199344 479528
rect 238208 479476 238260 479528
rect 374736 479476 374788 479528
rect 51724 479408 51776 479460
rect 116124 479408 116176 479460
rect 58532 479340 58584 479392
rect 123668 479340 123720 479392
rect 54760 479272 54812 479324
rect 116676 479272 116728 479324
rect 107752 478524 107804 478576
rect 108212 478524 108264 478576
rect 270592 478524 270644 478576
rect 358544 478524 358596 478576
rect 254860 478456 254912 478508
rect 358452 478456 358504 478508
rect 269396 478388 269448 478440
rect 373908 478388 373960 478440
rect 252744 478320 252796 478372
rect 374920 478320 374972 478372
rect 241704 478252 241756 478304
rect 367836 478252 367888 478304
rect 177028 478184 177080 478236
rect 204996 478184 205048 478236
rect 237472 478184 237524 478236
rect 363880 478184 363932 478236
rect 61660 478116 61712 478168
rect 199384 478116 199436 478168
rect 205824 478116 205876 478168
rect 217324 478116 217376 478168
rect 233332 478116 233384 478168
rect 366364 478116 366416 478168
rect 298008 478048 298060 478100
rect 298284 478048 298336 478100
rect 60740 477912 60792 477964
rect 61108 477912 61160 477964
rect 183652 477640 183704 477692
rect 184020 477640 184072 477692
rect 185032 477640 185084 477692
rect 185860 477640 185912 477692
rect 298192 477572 298244 477624
rect 299020 477572 299072 477624
rect 59636 477436 59688 477488
rect 135996 477436 136048 477488
rect 289268 477436 289320 477488
rect 373816 477436 373868 477488
rect 45376 477368 45428 477420
rect 123300 477368 123352 477420
rect 287336 477368 287388 477420
rect 379336 477368 379388 477420
rect 57428 477300 57480 477352
rect 135260 477300 135312 477352
rect 265164 477300 265216 477352
rect 362592 477300 362644 477352
rect 55956 477232 56008 477284
rect 133880 477232 133932 477284
rect 268108 477232 268160 477284
rect 366272 477232 366324 477284
rect 54484 477164 54536 477216
rect 133972 477164 134024 477216
rect 275652 477164 275704 477216
rect 373724 477164 373776 477216
rect 50068 477096 50120 477148
rect 131212 477096 131264 477148
rect 265072 477096 265124 477148
rect 365444 477096 365496 477148
rect 49056 477028 49108 477080
rect 130660 477028 130712 477080
rect 263692 477028 263744 477080
rect 368112 477028 368164 477080
rect 48964 476960 49016 477012
rect 132592 476960 132644 477012
rect 263784 476960 263836 477012
rect 375012 476960 375064 477012
rect 46296 476892 46348 476944
rect 132868 476892 132920 476944
rect 237380 476892 237432 476944
rect 366456 476892 366508 476944
rect 42156 476824 42208 476876
rect 131580 476824 131632 476876
rect 162952 476824 163004 476876
rect 207664 476824 207716 476876
rect 236828 476824 236880 476876
rect 365076 476824 365128 476876
rect 44732 476756 44784 476808
rect 143632 476756 143684 476808
rect 165712 476756 165764 476808
rect 218796 476756 218848 476808
rect 247040 476756 247092 476808
rect 376300 476756 376352 476808
rect 58440 476688 58492 476740
rect 128452 476688 128504 476740
rect 292764 476688 292816 476740
rect 375748 476688 375800 476740
rect 59820 476620 59872 476672
rect 127624 476620 127676 476672
rect 43996 476552 44048 476604
rect 80980 476552 81032 476604
rect 100852 476484 100904 476536
rect 101220 476484 101272 476536
rect 88432 476416 88484 476468
rect 88892 476416 88944 476468
rect 292580 475736 292632 475788
rect 376760 475736 376812 475788
rect 269120 475668 269172 475720
rect 374368 475668 374420 475720
rect 258908 475600 258960 475652
rect 372160 475600 372212 475652
rect 185032 475532 185084 475584
rect 213184 475532 213236 475584
rect 254032 475532 254084 475584
rect 379060 475532 379112 475584
rect 176752 475464 176804 475516
rect 207848 475464 207900 475516
rect 245292 475464 245344 475516
rect 370596 475464 370648 475516
rect 57612 475396 57664 475448
rect 114744 475396 114796 475448
rect 164608 475396 164660 475448
rect 211896 475396 211948 475448
rect 226616 475396 226668 475448
rect 363604 475396 363656 475448
rect 60832 475328 60884 475380
rect 199476 475328 199528 475380
rect 238760 475328 238812 475380
rect 378876 475328 378928 475380
rect 291936 474648 291988 474700
rect 368388 474648 368440 474700
rect 85672 474580 85724 474632
rect 85856 474580 85908 474632
rect 273444 474580 273496 474632
rect 361488 474580 361540 474632
rect 280436 474512 280488 474564
rect 369676 474512 369728 474564
rect 278228 474444 278280 474496
rect 368296 474444 368348 474496
rect 257620 474376 257672 474428
rect 362684 474376 362736 474428
rect 176660 474308 176712 474360
rect 209228 474308 209280 474360
rect 262588 474308 262640 474360
rect 373540 474308 373592 474360
rect 179788 474240 179840 474292
rect 216128 474240 216180 474292
rect 259460 474240 259512 474292
rect 373632 474240 373684 474292
rect 159364 474172 159416 474224
rect 218888 474172 218940 474224
rect 241612 474172 241664 474224
rect 361028 474172 361080 474224
rect 51632 474104 51684 474156
rect 99564 474104 99616 474156
rect 139492 474104 139544 474156
rect 205824 474104 205876 474156
rect 244280 474104 244332 474156
rect 371976 474104 372028 474156
rect 57796 474036 57848 474088
rect 113272 474036 113324 474088
rect 126980 474036 127032 474088
rect 201500 474036 201552 474088
rect 207204 474036 207256 474088
rect 217232 474036 217284 474088
rect 229836 474036 229888 474088
rect 363788 474036 363840 474088
rect 59360 473968 59412 474020
rect 180156 473968 180208 474020
rect 186412 473968 186464 474020
rect 212080 473968 212132 474020
rect 229192 473968 229244 474020
rect 363696 473968 363748 474020
rect 290188 473900 290240 473952
rect 357164 473900 357216 473952
rect 289820 473016 289872 473068
rect 360752 473016 360804 473068
rect 294052 472948 294104 473000
rect 369768 472948 369820 473000
rect 273352 472880 273404 472932
rect 362868 472880 362920 472932
rect 262312 472812 262364 472864
rect 370780 472812 370832 472864
rect 188068 472744 188120 472796
rect 210700 472744 210752 472796
rect 263600 472744 263652 472796
rect 372252 472744 372304 472796
rect 175372 472676 175424 472728
rect 202144 472676 202196 472728
rect 226432 472676 226484 472728
rect 367744 472676 367796 472728
rect 58624 472608 58676 472660
rect 110604 472608 110656 472660
rect 184940 472608 184992 472660
rect 212172 472608 212224 472660
rect 227720 472608 227772 472660
rect 374644 472608 374696 472660
rect 46204 471928 46256 471980
rect 64880 471928 64932 471980
rect 192760 471928 192812 471980
rect 213460 471928 213512 471980
rect 296260 471928 296312 471980
rect 362040 471928 362092 471980
rect 50988 471860 51040 471912
rect 82820 471860 82872 471912
rect 183100 471860 183152 471912
rect 205088 471860 205140 471912
rect 287152 471860 287204 471912
rect 358728 471860 358780 471912
rect 51540 471792 51592 471844
rect 84476 471792 84528 471844
rect 192024 471792 192076 471844
rect 217692 471792 217744 471844
rect 298192 471792 298244 471844
rect 372436 471792 372488 471844
rect 50620 471724 50672 471776
rect 82912 471724 82964 471776
rect 190644 471724 190696 471776
rect 216404 471724 216456 471776
rect 298100 471724 298152 471776
rect 372620 471724 372672 471776
rect 49424 471656 49476 471708
rect 83188 471656 83240 471708
rect 190552 471656 190604 471708
rect 217508 471656 217560 471708
rect 298284 471656 298336 471708
rect 375196 471656 375248 471708
rect 54668 471588 54720 471640
rect 100760 471588 100812 471640
rect 183652 471588 183704 471640
rect 210792 471588 210844 471640
rect 297732 471588 297784 471640
rect 375104 471588 375156 471640
rect 57336 471520 57388 471572
rect 103612 471520 103664 471572
rect 161572 471520 161624 471572
rect 214656 471520 214708 471572
rect 288532 471520 288584 471572
rect 371148 471520 371200 471572
rect 53288 471452 53340 471504
rect 100852 471452 100904 471504
rect 140964 471452 141016 471504
rect 200396 471452 200448 471504
rect 276940 471452 276992 471504
rect 358636 471452 358688 471504
rect 53196 471384 53248 471436
rect 100944 471384 100996 471436
rect 140872 471384 140924 471436
rect 203156 471384 203208 471436
rect 285864 471384 285916 471436
rect 376484 471384 376536 471436
rect 50252 471316 50304 471368
rect 98644 471316 98696 471368
rect 140780 471316 140832 471368
rect 205916 471316 205968 471368
rect 240140 471316 240192 471368
rect 362408 471316 362460 471368
rect 57704 471248 57756 471300
rect 113364 471248 113416 471300
rect 125692 471248 125744 471300
rect 196900 471248 196952 471300
rect 240232 471248 240284 471300
rect 363972 471248 364024 471300
rect 47400 471180 47452 471232
rect 65524 471180 65576 471232
rect 183560 471180 183612 471232
rect 203800 471180 203852 471232
rect 47492 471112 47544 471164
rect 64972 471112 65024 471164
rect 182364 471112 182416 471164
rect 202420 471112 202472 471164
rect 52092 471044 52144 471096
rect 68284 471044 68336 471096
rect 183744 471044 183796 471096
rect 200856 471044 200908 471096
rect 282920 470432 282972 470484
rect 358084 470432 358136 470484
rect 283104 470364 283156 470416
rect 359924 470364 359976 470416
rect 283012 470296 283064 470348
rect 359832 470296 359884 470348
rect 285680 470228 285732 470280
rect 364248 470228 364300 470280
rect 287060 470160 287112 470212
rect 367652 470160 367704 470212
rect 285772 470092 285824 470144
rect 377680 470092 377732 470144
rect 178132 470024 178184 470076
rect 202328 470024 202380 470076
rect 284300 470024 284352 470076
rect 377404 470024 377456 470076
rect 179512 469956 179564 470008
rect 206468 469956 206520 470008
rect 284392 469956 284444 470008
rect 377588 469956 377640 470008
rect 50804 469888 50856 469940
rect 81624 469888 81676 469940
rect 164240 469888 164292 469940
rect 218980 469888 219032 469940
rect 281540 469888 281592 469940
rect 376576 469888 376628 469940
rect 57520 469820 57572 469872
rect 111984 469820 112036 469872
rect 143540 469820 143592 469872
rect 210424 469820 210476 469872
rect 281632 469820 281684 469872
rect 379980 469820 380032 469872
rect 49516 469140 49568 469192
rect 80060 469140 80112 469192
rect 193404 469140 193456 469192
rect 216496 469140 216548 469192
rect 273260 469140 273312 469192
rect 363420 469140 363472 469192
rect 50712 469072 50764 469124
rect 78772 469072 78824 469124
rect 178040 469072 178092 469124
rect 210884 469072 210936 469124
rect 266544 469072 266596 469124
rect 359556 469072 359608 469124
rect 46020 469004 46072 469056
rect 63592 469004 63644 469056
rect 168564 469004 168616 469056
rect 202236 469004 202288 469056
rect 266452 469004 266504 469056
rect 359648 469004 359700 469056
rect 48780 468936 48832 468988
rect 70584 468936 70636 468988
rect 167092 468936 167144 468988
rect 209136 468936 209188 468988
rect 266360 468936 266412 468988
rect 361304 468936 361356 468988
rect 56140 468868 56192 468920
rect 85580 468868 85632 468920
rect 167184 468868 167236 468920
rect 210608 468868 210660 468920
rect 272064 468868 272116 468920
rect 369032 468868 369084 468920
rect 56232 468800 56284 468852
rect 87144 468800 87196 468852
rect 168472 468800 168524 468852
rect 214748 468800 214800 468852
rect 264980 468800 265032 468852
rect 364064 468800 364116 468852
rect 54944 468732 54996 468784
rect 86960 468732 87012 468784
rect 139400 468732 139452 468784
rect 196992 468732 197044 468784
rect 255320 468732 255372 468784
rect 361212 468732 361264 468784
rect 53380 468664 53432 468716
rect 85672 468664 85724 468716
rect 142344 468664 142396 468716
rect 200488 468664 200540 468716
rect 267740 468664 267792 468716
rect 377312 468664 377364 468716
rect 59912 468596 59964 468648
rect 92572 468596 92624 468648
rect 109040 468596 109092 468648
rect 197728 468596 197780 468648
rect 249984 468596 250036 468648
rect 365168 468596 365220 468648
rect 53472 468528 53524 468580
rect 87052 468528 87104 468580
rect 107844 468528 107896 468580
rect 198924 468528 198976 468580
rect 251364 468528 251416 468580
rect 369308 468528 369360 468580
rect 49332 468460 49384 468512
rect 93952 468460 94004 468512
rect 107752 468460 107804 468512
rect 203064 468460 203116 468512
rect 252560 468460 252612 468512
rect 376208 468460 376260 468512
rect 191932 468392 191984 468444
rect 214380 468392 214432 468444
rect 280160 468392 280212 468444
rect 363512 468392 363564 468444
rect 191840 468324 191892 468376
rect 211528 468324 211580 468376
rect 189172 468256 189224 468308
rect 208032 468256 208084 468308
rect 45100 467780 45152 467832
rect 73804 467780 73856 467832
rect 80704 467780 80756 467832
rect 178040 467780 178092 467832
rect 293960 467780 294012 467832
rect 357992 467780 358044 467832
rect 44824 467712 44876 467764
rect 73988 467712 74040 467764
rect 291292 467712 291344 467764
rect 362132 467712 362184 467764
rect 42524 467644 42576 467696
rect 73896 467644 73948 467696
rect 288440 467644 288492 467696
rect 364800 467644 364852 467696
rect 53104 467576 53156 467628
rect 99656 467576 99708 467628
rect 277492 467576 277544 467628
rect 370228 467576 370280 467628
rect 52368 467508 52420 467560
rect 99472 467508 99524 467560
rect 274640 467508 274692 467560
rect 367560 467508 367612 467560
rect 43904 467440 43956 467492
rect 93860 467440 93912 467492
rect 256700 467440 256752 467492
rect 361120 467440 361172 467492
rect 45008 467372 45060 467424
rect 105084 467372 105136 467424
rect 182180 467372 182232 467424
rect 212264 467372 212316 467424
rect 258172 467372 258224 467424
rect 368204 467372 368256 467424
rect 43444 467304 43496 467356
rect 103704 467304 103756 467356
rect 175280 467304 175332 467356
rect 206560 467304 206612 467356
rect 251272 467304 251324 467356
rect 365260 467304 365312 467356
rect 44916 467236 44968 467288
rect 104992 467236 105044 467288
rect 180156 467236 180208 467288
rect 218060 467236 218112 467288
rect 251180 467236 251232 467288
rect 366824 467236 366876 467288
rect 45284 467168 45336 467220
rect 106372 467168 106424 467220
rect 149060 467168 149112 467220
rect 212908 467168 212960 467220
rect 253940 467168 253992 467220
rect 369584 467168 369636 467220
rect 45192 467100 45244 467152
rect 106464 467100 106516 467152
rect 146300 467100 146352 467152
rect 218704 467100 218756 467152
rect 262220 467100 262272 467152
rect 379152 467100 379204 467152
rect 59268 467032 59320 467084
rect 67732 467032 67784 467084
rect 59176 466964 59228 467016
rect 66352 466964 66404 467016
rect 178040 466556 178092 466608
rect 204628 466556 204680 466608
rect 338488 466556 338540 466608
rect 356980 466556 357032 466608
rect 498476 466556 498528 466608
rect 517796 466556 517848 466608
rect 48872 466488 48924 466540
rect 218060 466488 218112 466540
rect 218244 466488 218296 466540
rect 339776 466488 339828 466540
rect 357532 466488 357584 466540
rect 499764 466488 499816 466540
rect 190920 466420 190972 466472
rect 206284 466420 206336 466472
rect 207112 466420 207164 466472
rect 208124 466420 208176 466472
rect 351000 466420 351052 466472
rect 358820 466420 358872 466472
rect 510896 466488 510948 466540
rect 517520 466488 517572 466540
rect 517888 466420 517940 466472
rect 52276 466352 52328 466404
rect 77300 466352 77352 466404
rect 193312 466352 193364 466404
rect 213092 466352 213144 466404
rect 295432 466352 295484 466404
rect 357256 466352 357308 466404
rect 52000 466284 52052 466336
rect 75920 466284 75972 466336
rect 180984 466284 181036 466336
rect 207940 466284 207992 466336
rect 271972 466284 272024 466336
rect 366180 466284 366232 466336
rect 189080 466216 189132 466268
rect 217600 466216 217652 466268
rect 258080 466216 258132 466268
rect 364156 466216 364208 466268
rect 54392 466148 54444 466200
rect 62120 466148 62172 466200
rect 173900 466148 173952 466200
rect 203892 466148 203944 466200
rect 260840 466148 260892 466200
rect 376392 466148 376444 466200
rect 54300 466080 54352 466132
rect 63500 466080 63552 466132
rect 180892 466080 180944 466132
rect 210976 466080 211028 466132
rect 249800 466080 249852 466132
rect 366548 466080 366600 466132
rect 51448 466012 51500 466064
rect 66260 466012 66312 466064
rect 172520 466012 172572 466064
rect 204904 466012 204956 466064
rect 245660 466012 245712 466064
rect 362500 466012 362552 466064
rect 42064 465944 42116 465996
rect 60740 465944 60792 465996
rect 179420 465944 179472 465996
rect 219072 465944 219124 465996
rect 249892 465944 249944 465996
rect 367928 465944 367980 465996
rect 43352 465876 43404 465928
rect 62212 465876 62264 465928
rect 173992 465876 174044 465928
rect 214840 465876 214892 465928
rect 248512 465876 248564 465928
rect 372068 465876 372120 465928
rect 56048 465808 56100 465860
rect 89812 465808 89864 465860
rect 142252 465808 142304 465860
rect 207112 465808 207164 465860
rect 248604 465808 248656 465860
rect 373448 465808 373500 465860
rect 50804 465740 50856 465792
rect 50988 465740 51040 465792
rect 51540 465740 51592 465792
rect 52000 465740 52052 465792
rect 58808 465740 58860 465792
rect 95424 465740 95476 465792
rect 107660 465740 107712 465792
rect 201776 465740 201828 465792
rect 208308 465740 208360 465792
rect 221004 465740 221056 465792
rect 241520 465740 241572 465792
rect 369400 465740 369452 465792
rect 49516 465672 49568 465724
rect 70400 465672 70452 465724
rect 72424 465672 72476 465724
rect 198832 465672 198884 465724
rect 205364 465672 205416 465724
rect 220912 465672 220964 465724
rect 242900 465672 242952 465724
rect 374828 465672 374880 465724
rect 186320 465604 186372 465656
rect 202512 465604 202564 465656
rect 187792 465536 187844 465588
rect 200948 465536 201000 465588
rect 194600 465468 194652 465520
rect 206652 465468 206704 465520
rect 198832 465060 198884 465112
rect 199016 465060 199068 465112
rect 358912 465060 358964 465112
rect 518900 465060 518952 465112
rect 190460 464788 190512 464840
rect 208952 464788 209004 464840
rect 58992 464720 59044 464772
rect 89904 464720 89956 464772
rect 185584 464720 185636 464772
rect 204720 464720 204772 464772
rect 58900 464652 58952 464704
rect 92664 464652 92716 464704
rect 193220 464652 193272 464704
rect 214288 464652 214340 464704
rect 55864 464584 55916 464636
rect 102324 464584 102376 464636
rect 180800 464584 180852 464636
rect 209320 464584 209372 464636
rect 54576 464516 54628 464568
rect 102232 464516 102284 464568
rect 142160 464516 142212 464568
rect 198096 464516 198148 464568
rect 52920 464448 52972 464500
rect 121460 464448 121512 464500
rect 125600 464448 125652 464500
rect 197820 464448 197872 464500
rect 295340 464448 295392 464500
rect 360660 464448 360712 464500
rect 57060 464380 57112 464432
rect 131120 464380 131172 464432
rect 138020 464380 138072 464432
rect 200580 464380 200632 464432
rect 291200 464380 291252 464432
rect 364892 464380 364944 464432
rect 57152 464312 57204 464364
rect 132500 464312 132552 464364
rect 136640 464312 136692 464364
rect 199568 464312 199620 464364
rect 271880 464312 271932 464364
rect 371608 464312 371660 464364
rect 519544 460164 519596 460216
rect 580356 460164 580408 460216
rect 48872 418072 48924 418124
rect 57060 418072 57112 418124
rect 204536 417732 204588 417784
rect 208216 417732 208268 417784
rect 208124 417392 208176 417444
rect 216680 417392 216732 417444
rect 359740 417392 359792 417444
rect 377220 417392 377272 417444
rect 55772 417120 55824 417172
rect 57244 417120 57296 417172
rect 44640 416780 44692 416832
rect 57244 416780 57296 416832
rect 56876 416168 56928 416220
rect 59636 416168 59688 416220
rect 205732 414808 205784 414860
rect 217140 414808 217192 414860
rect 205456 414672 205508 414724
rect 216772 414672 216824 414724
rect 51540 413992 51592 414044
rect 57060 413992 57112 414044
rect 55680 413924 55732 413976
rect 56968 413924 57020 413976
rect 205640 413244 205692 413296
rect 216864 413244 216916 413296
rect 50160 412700 50212 412752
rect 57244 412700 57296 412752
rect 358084 411884 358136 411936
rect 377220 411884 377272 411936
rect 204444 411544 204496 411596
rect 205640 411544 205692 411596
rect 49608 411272 49660 411324
rect 57244 411272 57296 411324
rect 2964 411204 3016 411256
rect 15844 411204 15896 411256
rect 52276 411068 52328 411120
rect 53012 411068 53064 411120
rect 206744 410660 206796 410712
rect 216956 410660 217008 410712
rect 205640 410524 205692 410576
rect 216680 410524 216732 410576
rect 359924 410524 359976 410576
rect 377220 410524 377272 410576
rect 377680 410524 377732 410576
rect 217692 410048 217744 410100
rect 219256 410048 219308 410100
rect 48872 409844 48924 409896
rect 56692 409844 56744 409896
rect 208216 409096 208268 409148
rect 216680 409096 216732 409148
rect 359832 409096 359884 409148
rect 377404 409096 377456 409148
rect 52368 408484 52420 408536
rect 57244 408484 57296 408536
rect 198832 400868 198884 400920
rect 199476 400868 199528 400920
rect 207204 400868 207256 400920
rect 520924 396720 520976 396772
rect 580356 396720 580408 396772
rect 198188 396312 198240 396364
rect 199200 396312 199252 396364
rect 198004 395972 198056 396024
rect 198832 395972 198884 396024
rect 198280 395496 198332 395548
rect 199568 395496 199620 395548
rect 44732 391892 44784 391944
rect 57244 391892 57296 391944
rect 209412 391892 209464 391944
rect 216680 391892 216732 391944
rect 359464 391892 359516 391944
rect 376944 391892 376996 391944
rect 358820 390464 358872 390516
rect 376944 390464 376996 390516
rect 206284 389784 206336 389836
rect 216680 389784 216732 389836
rect 57060 389512 57112 389564
rect 57428 389512 57480 389564
rect 358084 389172 358136 389224
rect 358820 389172 358872 389224
rect 53748 389104 53800 389156
rect 57244 389104 57296 389156
rect 57520 389104 57572 389156
rect 200764 389104 200816 389156
rect 217692 389104 217744 389156
rect 359648 389104 359700 389156
rect 376944 389104 376996 389156
rect 46112 389036 46164 389088
rect 57152 389036 57204 389088
rect 57060 388356 57112 388408
rect 57428 388356 57480 388408
rect 199292 384276 199344 384328
rect 199660 384276 199712 384328
rect 197176 382168 197228 382220
rect 197912 382168 197964 382220
rect 58532 381828 58584 381880
rect 59636 381828 59688 381880
rect 55864 381692 55916 381744
rect 59360 381692 59412 381744
rect 205548 381488 205600 381540
rect 212908 381488 212960 381540
rect 362040 381488 362092 381540
rect 369860 381488 369912 381540
rect 218244 381012 218296 381064
rect 57336 380944 57388 380996
rect 59452 380944 59504 380996
rect 195888 380944 195940 380996
rect 219532 380944 219584 380996
rect 220084 380944 220136 380996
rect 58440 380876 58492 380928
rect 60740 380876 60792 380928
rect 208400 380876 208452 380928
rect 208676 380876 208728 380928
rect 217600 380876 217652 380928
rect 248236 380876 248288 380928
rect 369860 380876 369912 380928
rect 371056 380876 371108 380928
rect 431132 380876 431184 380928
rect 44640 380808 44692 380860
rect 217232 380808 217284 380860
rect 219164 380808 219216 380860
rect 219348 380808 219400 380860
rect 219900 380808 219952 380860
rect 220728 380808 220780 380860
rect 52920 380740 52972 380792
rect 55864 380740 55916 380792
rect 50160 380672 50212 380724
rect 216864 380740 216916 380792
rect 217692 380740 217744 380792
rect 367008 380740 367060 380792
rect 380992 380740 381044 380792
rect 155960 380672 156012 380724
rect 203156 380672 203208 380724
rect 357992 380672 358044 380724
rect 380900 380672 380952 380724
rect 158536 380604 158588 380656
rect 205916 380604 205968 380656
rect 377312 380604 377364 380656
rect 410708 380604 410760 380656
rect 140964 380536 141016 380588
rect 200580 380536 200632 380588
rect 373908 380536 373960 380588
rect 421104 380536 421156 380588
rect 54484 380468 54536 380520
rect 113548 380468 113600 380520
rect 146024 380468 146076 380520
rect 205824 380468 205876 380520
rect 371608 380468 371660 380520
rect 433616 380468 433668 380520
rect 55956 380400 56008 380452
rect 118424 380400 118476 380452
rect 143540 380400 143592 380452
rect 204720 380400 204772 380452
rect 369032 380400 369084 380452
rect 436008 380400 436060 380452
rect 48964 380332 49016 380384
rect 110972 380332 111024 380384
rect 133512 380332 133564 380384
rect 201868 380332 201920 380384
rect 213644 380332 213696 380384
rect 222016 380332 222068 380384
rect 366180 380332 366232 380384
rect 438492 380332 438544 380384
rect 57428 380264 57480 380316
rect 123484 380264 123536 380316
rect 131028 380264 131080 380316
rect 198280 380264 198332 380316
rect 200120 380264 200172 380316
rect 295340 380264 295392 380316
rect 363420 380264 363472 380316
rect 440884 380264 440936 380316
rect 56876 380196 56928 380248
rect 125968 380196 126020 380248
rect 128360 380196 128412 380248
rect 199108 380196 199160 380248
rect 200212 380196 200264 380248
rect 301504 380196 301556 380248
rect 361488 380196 361540 380248
rect 443460 380196 443512 380248
rect 47584 380128 47636 380180
rect 116032 380128 116084 380180
rect 121000 380128 121052 380180
rect 198832 380128 198884 380180
rect 201684 380128 201736 380180
rect 310428 380128 310480 380180
rect 357072 380128 357124 380180
rect 485964 380128 486016 380180
rect 160928 380060 160980 380112
rect 207112 380060 207164 380112
rect 213552 380060 213604 380112
rect 213828 380060 213880 380112
rect 236000 380060 236052 380112
rect 163412 379992 163464 380044
rect 198096 379992 198148 380044
rect 215852 379992 215904 380044
rect 237104 379992 237156 380044
rect 239128 379992 239180 380044
rect 259460 379992 259512 380044
rect 165988 379924 166040 379976
rect 200488 379924 200540 379976
rect 213828 379924 213880 379976
rect 243084 379924 243136 379976
rect 219808 379856 219860 379908
rect 254492 379856 254544 379908
rect 215300 379788 215352 379840
rect 216220 379788 216272 379840
rect 256976 379788 257028 379840
rect 376484 379788 376536 379840
rect 405464 379788 405516 379840
rect 212540 379720 212592 379772
rect 255872 379720 255924 379772
rect 380992 379720 381044 379772
rect 381360 379720 381412 379772
rect 413468 379720 413520 379772
rect 212632 379652 212684 379704
rect 258080 379652 258132 379704
rect 380900 379652 380952 379704
rect 426440 379652 426492 379704
rect 212724 379584 212776 379636
rect 219808 379584 219860 379636
rect 219900 379584 219952 379636
rect 263876 379584 263928 379636
rect 368388 379584 368440 379636
rect 372528 379584 372580 379636
rect 419448 379584 419500 379636
rect 207112 379516 207164 379568
rect 213828 379516 213880 379568
rect 86592 379448 86644 379500
rect 208492 379448 208544 379500
rect 212448 379448 212500 379500
rect 219348 379448 219400 379500
rect 265256 379516 265308 379568
rect 374552 379516 374604 379568
rect 375104 379516 375156 379568
rect 434352 379516 434404 379568
rect 220084 379448 220136 379500
rect 275652 379448 275704 379500
rect 301504 379448 301556 379500
rect 313372 379448 313424 379500
rect 359556 379448 359608 379500
rect 408316 379448 408368 379500
rect 47768 379380 47820 379432
rect 88340 379380 88392 379432
rect 92388 379380 92440 379432
rect 212816 379380 212868 379432
rect 213828 379380 213880 379432
rect 219440 379380 219492 379432
rect 274364 379380 274416 379432
rect 310428 379380 310480 379432
rect 315764 379380 315816 379432
rect 372436 379380 372488 379432
rect 377404 379380 377456 379432
rect 88800 379312 88852 379364
rect 47676 379244 47728 379296
rect 90640 379244 90692 379296
rect 208492 379312 208544 379364
rect 209596 379312 209648 379364
rect 209872 379244 209924 379296
rect 219624 379312 219676 379364
rect 273260 379312 273312 379364
rect 295340 379312 295392 379364
rect 310980 379312 311032 379364
rect 91376 379176 91428 379228
rect 211344 379176 211396 379228
rect 218336 379244 218388 379296
rect 271052 379244 271104 379296
rect 59728 379108 59780 379160
rect 93492 379108 93544 379160
rect 93584 379108 93636 379160
rect 201408 379108 201460 379160
rect 46296 379040 46348 379092
rect 108212 379040 108264 379092
rect 108856 379040 108908 379092
rect 205456 379040 205508 379092
rect 210332 379040 210384 379092
rect 219532 379176 219584 379228
rect 220176 379176 220228 379228
rect 221004 379040 221056 379092
rect 373816 379040 373868 379092
rect 380900 379040 380952 379092
rect 42156 378972 42208 379024
rect 101036 378972 101088 379024
rect 112352 378972 112404 379024
rect 206836 378972 206888 379024
rect 212356 378972 212408 379024
rect 272156 378972 272208 379024
rect 379796 378972 379848 379024
rect 379980 378972 380032 379024
rect 397092 378972 397144 379024
rect 55680 378904 55732 378956
rect 103520 378904 103572 378956
rect 201408 378904 201460 378956
rect 220912 378904 220964 378956
rect 371148 378904 371200 378956
rect 379520 378904 379572 378956
rect 57060 378836 57112 378888
rect 104900 378836 104952 378888
rect 205640 378836 205692 378888
rect 206836 378836 206888 378888
rect 219440 378836 219492 378888
rect 220728 378836 220780 378888
rect 247592 378836 247644 378888
rect 376576 378836 376628 378888
rect 396080 378836 396132 378888
rect 55772 378768 55824 378820
rect 56968 378768 57020 378820
rect 222016 378768 222068 378820
rect 245384 378768 245436 378820
rect 358728 378768 358780 378820
rect 372620 378768 372672 378820
rect 377404 378768 377456 378820
rect 437848 378768 437900 378820
rect 50068 378700 50120 378752
rect 98460 378700 98512 378752
rect 211068 378700 211120 378752
rect 219716 378700 219768 378752
rect 49056 378632 49108 378684
rect 96068 378632 96120 378684
rect 46204 378564 46256 378616
rect 47676 378564 47728 378616
rect 113456 378564 113508 378616
rect 214196 378564 214248 378616
rect 219624 378564 219676 378616
rect 375288 378700 375340 378752
rect 400404 378700 400456 378752
rect 220176 378632 220228 378684
rect 248604 378632 248656 378684
rect 372712 378632 372764 378684
rect 373172 378632 373224 378684
rect 399484 378632 399536 378684
rect 250076 378564 250128 378616
rect 379336 378564 379388 378616
rect 379888 378564 379940 378616
rect 405832 378564 405884 378616
rect 114468 378496 114520 378548
rect 205640 378496 205692 378548
rect 213828 378496 213880 378548
rect 115848 378428 115900 378480
rect 213368 378428 213420 378480
rect 220084 378428 220136 378480
rect 221004 378496 221056 378548
rect 251180 378496 251232 378548
rect 380900 378496 380952 378548
rect 381176 378496 381228 378548
rect 412364 378496 412416 378548
rect 220820 378428 220872 378480
rect 252284 378428 252336 378480
rect 379520 378428 379572 378480
rect 411260 378428 411312 378480
rect 111340 378360 111392 378412
rect 208492 378360 208544 378412
rect 210332 378360 210384 378412
rect 268660 378360 268712 378412
rect 372620 378360 372672 378412
rect 373908 378360 373960 378412
rect 407580 378360 407632 378412
rect 90088 378292 90140 378344
rect 209780 378292 209832 378344
rect 211068 378292 211120 378344
rect 211712 378292 211764 378344
rect 212448 378292 212500 378344
rect 246212 378292 246264 378344
rect 273260 378292 273312 378344
rect 300860 378292 300912 378344
rect 342260 378292 342312 378344
rect 343180 378292 343232 378344
rect 360200 378292 360252 378344
rect 85488 378224 85540 378276
rect 208584 378224 208636 378276
rect 213000 378224 213052 378276
rect 213644 378224 213696 378276
rect 276020 378224 276072 378276
rect 277032 378224 277084 378276
rect 356612 378224 356664 378276
rect 375380 378292 375432 378344
rect 435180 378292 435232 378344
rect 503076 378224 503128 378276
rect 517612 378224 517664 378276
rect 580264 378224 580316 378276
rect 47676 378156 47728 378208
rect 80428 378156 80480 378208
rect 87880 378156 87932 378208
rect 219624 378156 219676 378208
rect 220728 378156 220780 378208
rect 220912 378156 220964 378208
rect 221188 378156 221240 378208
rect 253388 378156 253440 378208
rect 271788 378156 271840 378208
rect 305828 378156 305880 378208
rect 343548 378156 343600 378208
rect 503536 378156 503588 378208
rect 517704 378156 517756 378208
rect 580172 378156 580224 378208
rect 196716 378088 196768 378140
rect 287612 378088 287664 378140
rect 372344 378088 372396 378140
rect 474832 378088 474884 378140
rect 42064 378020 42116 378072
rect 199476 378020 199528 378072
rect 203984 378020 204036 378072
rect 317420 378020 317472 378072
rect 364248 378020 364300 378072
rect 375288 378020 375340 378072
rect 375840 378020 375892 378072
rect 460940 378020 460992 378072
rect 197452 377952 197504 378004
rect 298468 377952 298520 378004
rect 374460 377952 374512 378004
rect 458364 377952 458416 378004
rect 54392 377884 54444 377936
rect 183468 377884 183520 377936
rect 197636 377884 197688 377936
rect 295432 377884 295484 377936
rect 362868 377884 362920 377936
rect 445852 377884 445904 377936
rect 54300 377816 54352 377868
rect 182272 377816 182324 377868
rect 182824 377816 182876 377868
rect 197544 377816 197596 377868
rect 292672 377816 292724 377868
rect 367560 377816 367612 377868
rect 451004 377816 451056 377868
rect 95976 377748 96028 377800
rect 212540 377748 212592 377800
rect 213276 377748 213328 377800
rect 98276 377680 98328 377732
rect 212632 377680 212684 377732
rect 215760 377748 215812 377800
rect 217416 377748 217468 377800
rect 307852 377748 307904 377800
rect 370412 377748 370464 377800
rect 453028 377748 453080 377800
rect 214932 377680 214984 377732
rect 303252 377680 303304 377732
rect 373724 377680 373776 377732
rect 455512 377680 455564 377732
rect 196808 377612 196860 377664
rect 290924 377612 290976 377664
rect 365536 377612 365588 377664
rect 447508 377612 447560 377664
rect 196624 377544 196676 377596
rect 285956 377544 286008 377596
rect 358544 377544 358596 377596
rect 425980 377544 426032 377596
rect 197084 377476 197136 377528
rect 278228 377476 278280 377528
rect 361396 377476 361448 377528
rect 415676 377476 415728 377528
rect 43352 377408 43404 377460
rect 199568 377408 199620 377460
rect 199752 377408 199804 377460
rect 273260 377408 273312 377460
rect 360752 377408 360804 377460
rect 150992 377340 151044 377392
rect 198188 377340 198240 377392
rect 198740 377340 198792 377392
rect 271788 377340 271840 377392
rect 376668 377408 376720 377460
rect 416872 377408 416924 377460
rect 375196 377340 375248 377392
rect 415860 377340 415912 377392
rect 138480 377272 138532 377324
rect 207296 377272 207348 377324
rect 211620 377272 211672 377324
rect 280252 377272 280304 377324
rect 364800 377272 364852 377324
rect 379336 377272 379388 377324
rect 409972 377272 410024 377324
rect 48872 377204 48924 377256
rect 216772 377204 216824 377256
rect 216956 377204 217008 377256
rect 374552 377204 374604 377256
rect 375288 377204 375340 377256
rect 402980 377204 403032 377256
rect 154028 377136 154080 377188
rect 200396 377136 200448 377188
rect 213000 377136 213052 377188
rect 213552 377136 213604 377188
rect 362132 377136 362184 377188
rect 375932 377136 375984 377188
rect 376668 377136 376720 377188
rect 380992 377136 381044 377188
rect 381360 377136 381412 377188
rect 374460 377068 374512 377120
rect 375288 377068 375340 377120
rect 376484 377000 376536 377052
rect 376668 377000 376720 377052
rect 375380 376864 375432 376916
rect 376484 376864 376536 376916
rect 368388 376728 368440 376780
rect 372620 376728 372672 376780
rect 77208 376660 77260 376712
rect 204352 376660 204404 376712
rect 215852 376660 215904 376712
rect 362776 376660 362828 376712
rect 477592 376660 477644 376712
rect 206652 376592 206704 376644
rect 283380 376592 283432 376644
rect 369676 376592 369728 376644
rect 483388 376592 483440 376644
rect 135904 376524 135956 376576
rect 200304 376524 200356 376576
rect 201592 376524 201644 376576
rect 320916 376524 320968 376576
rect 365628 376524 365680 376576
rect 473452 376524 473504 376576
rect 94688 376456 94740 376508
rect 212724 376456 212776 376508
rect 214288 376456 214340 376508
rect 276112 376456 276164 376508
rect 358636 376456 358688 376508
rect 463516 376456 463568 376508
rect 83280 376388 83332 376440
rect 207112 376388 207164 376440
rect 213092 376388 213144 376440
rect 273444 376388 273496 376440
rect 368296 376388 368348 376440
rect 470784 376388 470836 376440
rect 99472 376320 99524 376372
rect 214012 376320 214064 376372
rect 216496 376320 216548 376372
rect 270960 376320 271012 376372
rect 370228 376320 370280 376372
rect 467932 376320 467984 376372
rect 148692 376252 148744 376304
rect 196992 376252 197044 376304
rect 213460 376252 213512 376304
rect 268108 376252 268160 376304
rect 366916 376252 366968 376304
rect 430672 376252 430724 376304
rect 211528 376184 211580 376236
rect 265900 376184 265952 376236
rect 372620 376184 372672 376236
rect 436192 376184 436244 376236
rect 214380 376116 214432 376168
rect 263600 376116 263652 376168
rect 374368 376116 374420 376168
rect 422852 376116 422904 376168
rect 208032 376048 208084 376100
rect 250628 376048 250680 376100
rect 366272 376048 366324 376100
rect 413284 376048 413336 376100
rect 97816 375980 97868 376032
rect 215024 375980 215076 376032
rect 215300 375980 215352 376032
rect 219256 375980 219308 376032
rect 260932 375980 260984 376032
rect 377496 375980 377548 376032
rect 418436 375980 418488 376032
rect 208952 375912 209004 375964
rect 258356 375912 258408 375964
rect 357164 375912 357216 375964
rect 379980 375912 380032 375964
rect 414572 375912 414624 375964
rect 100852 375844 100904 375896
rect 214472 375844 214524 375896
rect 216404 375844 216456 375896
rect 255964 375844 256016 375896
rect 217508 375776 217560 375828
rect 253572 375776 253624 375828
rect 202880 375708 202932 375760
rect 325884 375708 325936 375760
rect 105728 375640 105780 375692
rect 218520 375640 218572 375692
rect 219348 375640 219400 375692
rect 372988 375368 373040 375420
rect 376760 375368 376812 375420
rect 377404 375368 377456 375420
rect 84384 375300 84436 375352
rect 208400 375300 208452 375352
rect 208676 375300 208728 375352
rect 102968 375232 103020 375284
rect 215392 375300 215444 375352
rect 217232 375300 217284 375352
rect 372436 375300 372488 375352
rect 379704 375300 379756 375352
rect 432236 375300 432288 375352
rect 213920 375232 213972 375284
rect 216496 375232 216548 375284
rect 369768 375232 369820 375284
rect 376760 375232 376812 375284
rect 425152 375232 425204 375284
rect 101864 375164 101916 375216
rect 375748 375164 375800 375216
rect 421196 375164 421248 375216
rect 107568 375096 107620 375148
rect 106464 375028 106516 375080
rect 377404 375096 377456 375148
rect 420644 375096 420696 375148
rect 367652 375028 367704 375080
rect 377496 375028 377548 375080
rect 408684 375028 408736 375080
rect 208400 374824 208452 374876
rect 216404 374960 216456 375012
rect 244280 374960 244332 375012
rect 216496 374892 216548 374944
rect 261668 374892 261720 374944
rect 364892 374892 364944 374944
rect 377128 374960 377180 375012
rect 418160 374960 418212 375012
rect 378140 374892 378192 374944
rect 423956 374892 424008 374944
rect 217232 374824 217284 374876
rect 262772 374824 262824 374876
rect 370320 374824 370372 374876
rect 374000 374824 374052 374876
rect 422668 374824 422720 374876
rect 211068 374756 211120 374808
rect 219440 374756 219492 374808
rect 267556 374756 267608 374808
rect 360660 374756 360712 374808
rect 372344 374756 372396 374808
rect 429660 374756 429712 374808
rect 206744 374688 206796 374740
rect 219348 374688 219400 374740
rect 266360 374688 266412 374740
rect 428556 374688 428608 374740
rect 183468 374620 183520 374672
rect 197636 374620 197688 374672
rect 342260 374620 342312 374672
rect 357256 374620 357308 374672
rect 369676 374620 369728 374672
rect 371700 374620 371752 374672
rect 378140 374620 378192 374672
rect 379428 374620 379480 374672
rect 439044 374620 439096 374672
rect 199384 371832 199436 371884
rect 199568 371832 199620 371884
rect 359188 371832 359240 371884
rect 359464 371832 359516 371884
rect 359740 371832 359792 371884
rect 519360 371900 519412 371952
rect 519544 371900 519596 371952
rect 199476 370472 199528 370524
rect 359096 370472 359148 370524
rect 359096 369860 359148 369912
rect 359648 369860 359700 369912
rect 207020 369792 207072 369844
rect 207204 369792 207256 369844
rect 359004 369792 359056 369844
rect 199568 369112 199620 369164
rect 207020 369112 207072 369164
rect 359464 369112 359516 369164
rect 519176 369112 519228 369164
rect 359004 366324 359056 366376
rect 359556 366324 359608 366376
rect 519084 366324 519136 366376
rect 519360 366324 519412 366376
rect 359648 363672 359700 363724
rect 518900 363672 518952 363724
rect 199752 363604 199804 363656
rect 359004 363604 359056 363656
rect 359004 362924 359056 362976
rect 359740 362924 359792 362976
rect 199660 362176 199712 362228
rect 359188 362176 359240 362228
rect 519084 362176 519136 362228
rect 519268 362176 519320 362228
rect 201408 360204 201460 360256
rect 206284 360204 206336 360256
rect 180156 360136 180208 360188
rect 195888 360136 195940 360188
rect 195888 359660 195940 359712
rect 197544 359660 197596 359712
rect 340052 359592 340104 359644
rect 357532 359592 357584 359644
rect 500408 359592 500460 359644
rect 517980 359592 518032 359644
rect 197360 359524 197412 359576
rect 204628 359524 204680 359576
rect 338488 359524 338540 359576
rect 356980 359524 357032 359576
rect 498936 359524 498988 359576
rect 517796 359524 517848 359576
rect 190920 359456 190972 359508
rect 200764 359456 200816 359508
rect 201408 359456 201460 359508
rect 351736 359456 351788 359508
rect 358084 359456 358136 359508
rect 178592 358776 178644 358828
rect 197360 358776 197412 358828
rect 342260 358776 342312 358828
rect 343548 358776 343600 358828
rect 358820 358776 358872 358828
rect 510896 358776 510948 358828
rect 517520 358776 517572 358828
rect 219256 358708 219308 358760
rect 220820 358708 220872 358760
rect 57152 358640 57204 358692
rect 59452 358640 59504 358692
rect 218612 358640 218664 358692
rect 221004 358640 221056 358692
rect 377036 358572 377088 358624
rect 381176 358572 381228 358624
rect 217140 358232 217192 358284
rect 219440 358232 219492 358284
rect 379244 358096 379296 358148
rect 380992 358096 381044 358148
rect 54484 358028 54536 358080
rect 59360 358028 59412 358080
rect 182824 358028 182876 358080
rect 201592 358028 201644 358080
rect 342260 358028 342312 358080
rect 373816 358028 373868 358080
rect 381084 358028 381136 358080
rect 379428 357960 379480 358012
rect 381268 357960 381320 358012
rect 219164 357824 219216 357876
rect 220912 357824 220964 357876
rect 378692 357824 378744 357876
rect 380900 357824 380952 357876
rect 58532 357348 58584 357400
rect 60740 357348 60792 357400
rect 46388 303560 46440 303612
rect 57336 303560 57388 303612
rect 57520 303560 57572 303612
rect 46480 300772 46532 300824
rect 56784 300772 56836 300824
rect 56968 300772 57020 300824
rect 58440 300772 58492 300824
rect 57060 300704 57112 300756
rect 520188 288396 520240 288448
rect 580264 288396 580316 288448
rect 518992 287036 519044 287088
rect 580356 287036 580408 287088
rect 200948 284248 201000 284300
rect 216680 284248 216732 284300
rect 361304 284248 361356 284300
rect 376852 284248 376904 284300
rect 203892 282820 203944 282872
rect 216772 282820 216824 282872
rect 366824 282820 366876 282872
rect 377588 282820 377640 282872
rect 55864 282616 55916 282668
rect 58624 282616 58676 282668
rect 51540 282140 51592 282192
rect 58348 282140 58400 282192
rect 200764 282140 200816 282192
rect 201408 282140 201460 282192
rect 216680 282140 216732 282192
rect 358084 282140 358136 282192
rect 376944 282140 376996 282192
rect 370412 273912 370464 273964
rect 370872 273912 370924 273964
rect 43628 273572 43680 273624
rect 133420 273572 133472 273624
rect 371056 273572 371108 273624
rect 378140 273572 378192 273624
rect 378692 273572 378744 273624
rect 379704 273572 379756 273624
rect 426440 273572 426492 273624
rect 44824 273504 44876 273556
rect 135904 273504 135956 273556
rect 369492 273504 369544 273556
rect 421104 273504 421156 273556
rect 44916 273436 44968 273488
rect 138480 273436 138532 273488
rect 370964 273436 371016 273488
rect 373080 273436 373132 273488
rect 431132 273436 431184 273488
rect 45008 273368 45060 273420
rect 140872 273368 140924 273420
rect 219348 273368 219400 273420
rect 219900 273368 219952 273420
rect 266360 273368 266412 273420
rect 373816 273368 373868 273420
rect 433340 273368 433392 273420
rect 45100 273300 45152 273352
rect 143540 273300 143592 273352
rect 214196 273300 214248 273352
rect 214932 273300 214984 273352
rect 273260 273300 273312 273352
rect 356888 273300 356940 273352
rect 430948 273300 431000 273352
rect 45192 273232 45244 273284
rect 145932 273232 145984 273284
rect 210976 273232 211028 273284
rect 283472 273232 283524 273284
rect 369768 273232 369820 273284
rect 373632 273232 373684 273284
rect 453396 273232 453448 273284
rect 374000 273164 374052 273216
rect 422852 273164 422904 273216
rect 361212 273096 361264 273148
rect 425980 273096 426032 273148
rect 46664 273028 46716 273080
rect 51540 273028 51592 273080
rect 95884 273028 95936 273080
rect 209320 273028 209372 273080
rect 288164 273028 288216 273080
rect 358452 273028 358504 273080
rect 423404 273028 423456 273080
rect 49148 272960 49200 273012
rect 54300 272960 54352 273012
rect 83004 272960 83056 273012
rect 207940 272960 207992 273012
rect 285956 272960 286008 273012
rect 370780 272960 370832 273012
rect 468484 272960 468536 273012
rect 58440 272892 58492 272944
rect 61016 272892 61068 272944
rect 61476 272892 61528 272944
rect 212264 272892 212316 272944
rect 295892 272892 295944 272944
rect 372252 272892 372304 272944
rect 470876 272892 470928 272944
rect 202420 272824 202472 272876
rect 290924 272824 290976 272876
rect 375012 272824 375064 272876
rect 473452 272824 473504 272876
rect 50344 272756 50396 272808
rect 53840 272756 53892 272808
rect 210792 272756 210844 272808
rect 303436 272756 303488 272808
rect 368112 272756 368164 272808
rect 475844 272756 475896 272808
rect 50436 272688 50488 272740
rect 90732 272688 90784 272740
rect 205088 272688 205140 272740
rect 298468 272688 298520 272740
rect 365444 272688 365496 272740
rect 478420 272688 478472 272740
rect 48044 272620 48096 272672
rect 93676 272620 93728 272672
rect 200856 272620 200908 272672
rect 300860 272620 300912 272672
rect 362592 272620 362644 272672
rect 480812 272620 480864 272672
rect 49240 272552 49292 272604
rect 96068 272552 96120 272604
rect 203800 272552 203852 272604
rect 305828 272552 305880 272604
rect 364064 272552 364116 272604
rect 483204 272552 483256 272604
rect 51908 272484 51960 272536
rect 98460 272484 98512 272536
rect 47860 272416 47912 272468
rect 77116 272416 77168 272468
rect 98092 272416 98144 272468
rect 197176 272484 197228 272536
rect 202512 272484 202564 272536
rect 320916 272484 320968 272536
rect 366732 272484 366784 272536
rect 485964 272484 486016 272536
rect 378140 272416 378192 272468
rect 423772 272416 423824 272468
rect 46572 272348 46624 272400
rect 76012 272348 76064 272400
rect 59636 272280 59688 272332
rect 60832 272280 60884 272332
rect 62212 272280 62264 272332
rect 94412 272280 94464 272332
rect 54116 272212 54168 272264
rect 54760 272212 54812 272264
rect 87604 272212 87656 272264
rect 58348 272144 58400 272196
rect 59728 272144 59780 272196
rect 99380 272144 99432 272196
rect 58624 272076 58676 272128
rect 100760 272076 100812 272128
rect 356888 272076 356940 272128
rect 358820 272076 358872 272128
rect 47952 272008 48004 272060
rect 52828 272008 52880 272060
rect 96620 272008 96672 272060
rect 85764 271940 85816 271992
rect 106556 271940 106608 271992
rect 427084 271940 427136 271992
rect 436100 271940 436152 271992
rect 60832 271872 60884 271924
rect 106280 271872 106332 271924
rect 112352 271872 112404 271924
rect 196624 271872 196676 271924
rect 396724 271872 396776 271924
rect 415860 271872 415912 271924
rect 425704 271872 425756 271924
rect 427820 271872 427872 271924
rect 42432 271804 42484 271856
rect 123116 271804 123168 271856
rect 154488 271804 154540 271856
rect 201776 271804 201828 271856
rect 213184 271804 213236 271856
rect 313280 271804 313332 271856
rect 358360 271804 358412 271856
rect 455788 271804 455840 271856
rect 517704 271804 517756 271856
rect 517888 271804 517940 271856
rect 57152 271736 57204 271788
rect 128360 271736 128412 271788
rect 151360 271736 151412 271788
rect 198924 271736 198976 271788
rect 212172 271736 212224 271788
rect 307760 271736 307812 271788
rect 368020 271736 368072 271788
rect 458180 271736 458232 271788
rect 54484 271668 54536 271720
rect 125600 271668 125652 271720
rect 157248 271668 157300 271720
rect 203064 271668 203116 271720
rect 206468 271668 206520 271720
rect 280252 271668 280304 271720
rect 365352 271668 365404 271720
rect 447140 271668 447192 271720
rect 54576 271600 54628 271652
rect 120080 271600 120132 271652
rect 158628 271600 158680 271652
rect 198372 271600 198424 271652
rect 202328 271600 202380 271652
rect 270500 271600 270552 271652
rect 370688 271600 370740 271652
rect 449900 271600 449952 271652
rect 54668 271532 54720 271584
rect 117320 271532 117372 271584
rect 161296 271532 161348 271584
rect 204812 271532 204864 271584
rect 216128 271532 216180 271584
rect 276020 271532 276072 271584
rect 364156 271532 364208 271584
rect 443000 271532 443052 271584
rect 53196 271464 53248 271516
rect 115940 271464 115992 271516
rect 164148 271464 164200 271516
rect 197728 271464 197780 271516
rect 204996 271464 205048 271516
rect 263600 271464 263652 271516
rect 362684 271464 362736 271516
rect 437480 271464 437532 271516
rect 53104 271396 53156 271448
rect 52920 271328 52972 271380
rect 53012 271260 53064 271312
rect 51632 271192 51684 271244
rect 104900 271192 104952 271244
rect 51816 271124 51868 271176
rect 103520 271124 103572 271176
rect 50252 271056 50304 271108
rect 100760 271056 100812 271108
rect 197360 271396 197412 271448
rect 197636 271396 197688 271448
rect 219072 271396 219124 271448
rect 277952 271396 278004 271448
rect 343548 271396 343600 271448
rect 356888 271396 356940 271448
rect 372160 271396 372212 271448
rect 445760 271396 445812 271448
rect 210884 271328 210936 271380
rect 268016 271328 268068 271380
rect 361120 271328 361172 271380
rect 433340 271328 433392 271380
rect 183468 271260 183520 271312
rect 197360 271260 197412 271312
rect 209228 271260 209280 271312
rect 264980 271260 265032 271312
rect 343456 271260 343508 271312
rect 360200 271260 360252 271312
rect 368204 271260 368256 271312
rect 440240 271260 440292 271312
rect 503628 271260 503680 271312
rect 517612 271260 517664 271312
rect 113180 271192 113232 271244
rect 207848 271192 207900 271244
rect 260840 271192 260892 271244
rect 280068 271192 280120 271244
rect 357440 271192 357492 271244
rect 366640 271192 366692 271244
rect 434720 271192 434772 271244
rect 110420 271124 110472 271176
rect 183468 271124 183520 271176
rect 201592 271124 201644 271176
rect 206376 271124 206428 271176
rect 258264 271124 258316 271176
rect 277216 271124 277268 271176
rect 356612 271124 356664 271176
rect 369584 271124 369636 271176
rect 416044 271124 416096 271176
rect 503536 271124 503588 271176
rect 517888 271124 517940 271176
rect 107660 271056 107712 271108
rect 202144 271056 202196 271108
rect 252560 271056 252612 271108
rect 379060 271056 379112 271108
rect 418160 271056 418212 271108
rect 54852 270988 54904 271040
rect 88340 270988 88392 271040
rect 106924 270988 106976 271040
rect 113272 270988 113324 271040
rect 206560 270988 206612 271040
rect 255320 270988 255372 271040
rect 376208 270988 376260 271040
rect 412732 270988 412784 271040
rect 46112 270920 46164 270972
rect 77300 270920 77352 270972
rect 214840 270920 214892 270972
rect 247040 270920 247092 270972
rect 374920 270920 374972 270972
rect 409880 270920 409932 270972
rect 43444 270444 43496 270496
rect 129740 270444 129792 270496
rect 196716 270444 196768 270496
rect 197820 270444 197872 270496
rect 211712 270444 211764 270496
rect 212356 270444 212408 270496
rect 213092 270444 213144 270496
rect 213552 270444 213604 270496
rect 220544 270444 220596 270496
rect 248512 270444 248564 270496
rect 50528 270376 50580 270428
rect 84200 270376 84252 270428
rect 220728 270376 220780 270428
rect 247040 270376 247092 270428
rect 377036 270376 377088 270428
rect 378048 270376 378100 270428
rect 411260 270444 411312 270496
rect 380532 270376 380584 270428
rect 411352 270376 411404 270428
rect 81440 270308 81492 270360
rect 107660 270308 107712 270360
rect 218612 270308 218664 270360
rect 219348 270308 219400 270360
rect 252560 270308 252612 270360
rect 370964 270308 371016 270360
rect 401692 270308 401744 270360
rect 80060 270240 80112 270292
rect 109224 270240 109276 270292
rect 212356 270240 212408 270292
rect 245660 270240 245712 270292
rect 379244 270240 379296 270292
rect 379428 270240 379480 270292
rect 63500 270172 63552 270224
rect 92480 270172 92532 270224
rect 219164 270172 219216 270224
rect 251180 270172 251232 270224
rect 376668 270172 376720 270224
rect 404360 270240 404412 270292
rect 379888 270172 379940 270224
rect 405740 270172 405792 270224
rect 51724 270104 51776 270156
rect 54576 270104 54628 270156
rect 84660 270104 84712 270156
rect 216772 270104 216824 270156
rect 219256 270104 219308 270156
rect 251272 270104 251324 270156
rect 373172 270104 373224 270156
rect 398840 270104 398892 270156
rect 57980 270036 58032 270088
rect 91100 270036 91152 270088
rect 213552 270036 213604 270088
rect 244280 270036 244332 270088
rect 373908 270036 373960 270088
rect 374460 270036 374512 270088
rect 375104 270036 375156 270088
rect 400220 270036 400272 270088
rect 53196 269968 53248 270020
rect 58624 269968 58676 270020
rect 77392 269968 77444 270020
rect 110420 269968 110472 270020
rect 220360 269968 220412 270020
rect 249800 269968 249852 270020
rect 370412 269968 370464 270020
rect 373724 269968 373776 270020
rect 397460 269968 397512 270020
rect 55956 269900 56008 269952
rect 88340 269900 88392 269952
rect 220636 269900 220688 269952
rect 262220 269900 262272 269952
rect 371792 269900 371844 269952
rect 373632 269900 373684 269952
rect 403348 269900 403400 269952
rect 57152 269832 57204 269884
rect 89720 269832 89772 269884
rect 115848 269832 115900 269884
rect 197728 269832 197780 269884
rect 201500 269832 201552 269884
rect 220728 269832 220780 269884
rect 265164 269832 265216 269884
rect 374460 269832 374512 269884
rect 407120 269832 407172 269884
rect 51724 269764 51776 269816
rect 85580 269764 85632 269816
rect 113364 269764 113416 269816
rect 196716 269764 196768 269816
rect 217140 269764 217192 269816
rect 218612 269764 218664 269816
rect 266360 269764 266412 269816
rect 372252 269764 372304 269816
rect 375104 269764 375156 269816
rect 379520 269764 379572 269816
rect 413008 269764 413060 269816
rect 205272 269696 205324 269748
rect 209504 269696 209556 269748
rect 237380 269696 237432 269748
rect 376484 269696 376536 269748
rect 377128 269696 377180 269748
rect 391940 269696 391992 269748
rect 212264 269628 212316 269680
rect 271880 269628 271932 269680
rect 375104 269628 375156 269680
rect 380164 269628 380216 269680
rect 216680 269560 216732 269612
rect 217968 269560 218020 269612
rect 263600 269560 263652 269612
rect 378416 269560 378468 269612
rect 379612 269560 379664 269612
rect 380532 269560 380584 269612
rect 214380 269492 214432 269544
rect 219532 269492 219584 269544
rect 220544 269492 220596 269544
rect 378600 269492 378652 269544
rect 379888 269492 379940 269544
rect 215852 269424 215904 269476
rect 219716 269424 219768 269476
rect 220360 269424 220412 269476
rect 218520 269356 218572 269408
rect 219624 269356 219676 269408
rect 220728 269356 220780 269408
rect 217232 269220 217284 269272
rect 219440 269220 219492 269272
rect 220636 269220 220688 269272
rect 370780 269084 370832 269136
rect 373172 269084 373224 269136
rect 46756 269016 46808 269068
rect 51724 269016 51776 269068
rect 210332 269016 210384 269068
rect 210884 269016 210936 269068
rect 213276 269016 213328 269068
rect 216128 269016 216180 269068
rect 216404 269016 216456 269068
rect 219072 269016 219124 269068
rect 43720 268948 43772 269000
rect 57980 268948 58032 269000
rect 215760 268948 215812 269000
rect 218520 268948 218572 269000
rect 45468 268880 45520 268932
rect 57152 268880 57204 268932
rect 215024 268880 215076 268932
rect 217140 268880 217192 268932
rect 48228 268812 48280 268864
rect 55956 268812 56008 268864
rect 210884 268812 210936 268864
rect 267924 269016 267976 269068
rect 374368 269016 374420 269068
rect 375932 269016 375984 269068
rect 416780 269016 416832 269068
rect 219808 268948 219860 269000
rect 253940 268948 253992 269000
rect 379980 268948 380032 269000
rect 414020 268948 414072 269000
rect 232504 268880 232556 268932
rect 259460 268880 259512 268932
rect 387892 268880 387944 268932
rect 420920 268880 420972 268932
rect 231124 268812 231176 268864
rect 259552 268812 259604 268864
rect 377496 268812 377548 268864
rect 377956 268812 378008 268864
rect 408500 268812 408552 268864
rect 45284 268744 45336 268796
rect 147680 268744 147732 268796
rect 216496 268744 216548 268796
rect 229100 268744 229152 268796
rect 260840 268744 260892 268796
rect 379152 268744 379204 268796
rect 379336 268744 379388 268796
rect 409880 268744 409932 268796
rect 216128 268676 216180 268728
rect 255320 268676 255372 268728
rect 390560 268676 390612 268728
rect 419540 268676 419592 268728
rect 49240 268608 49292 268660
rect 63500 268608 63552 268660
rect 213736 268608 213788 268660
rect 216496 268608 216548 268660
rect 217140 268608 217192 268660
rect 256700 268608 256752 268660
rect 391940 268608 391992 268660
rect 418160 268608 418212 268660
rect 49056 268540 49108 268592
rect 80060 268540 80112 268592
rect 218520 268540 218572 268592
rect 258080 268540 258132 268592
rect 42340 268472 42392 268524
rect 46664 268472 46716 268524
rect 81440 268472 81492 268524
rect 208216 268472 208268 268524
rect 213644 268472 213696 268524
rect 269120 268472 269172 268524
rect 43812 268404 43864 268456
rect 49240 268404 49292 268456
rect 58716 268404 58768 268456
rect 104900 268404 104952 268456
rect 209596 268404 209648 268456
rect 212172 268404 212224 268456
rect 270500 268404 270552 268456
rect 43536 268336 43588 268388
rect 49056 268336 49108 268388
rect 50436 268336 50488 268388
rect 98092 268336 98144 268388
rect 206836 268336 206888 268388
rect 213460 268336 213512 268388
rect 273168 268336 273220 268388
rect 374552 268336 374604 268388
rect 376576 268336 376628 268388
rect 402980 268336 403032 268388
rect 216496 268268 216548 268320
rect 242900 268268 242952 268320
rect 219072 268200 219124 268252
rect 244372 268200 244424 268252
rect 45376 267656 45428 267708
rect 58072 267656 58124 267708
rect 213368 267656 213420 267708
rect 274640 267656 274692 267708
rect 377680 267656 377732 267708
rect 437480 267656 437532 267708
rect 216312 267588 216364 267640
rect 277400 267588 277452 267640
rect 380072 267588 380124 267640
rect 438860 267588 438912 267640
rect 375288 267520 375340 267572
rect 433340 267520 433392 267572
rect 58072 267180 58124 267232
rect 58716 267180 58768 267232
rect 379060 266364 379112 266416
rect 380072 266364 380124 266416
rect 191748 253852 191800 253904
rect 201408 253852 201460 253904
rect 202880 253852 202932 253904
rect 339408 253852 339460 253904
rect 356980 253920 357032 253972
rect 357808 253920 357860 253972
rect 500868 253308 500920 253360
rect 517704 253308 517756 253360
rect 180524 253240 180576 253292
rect 197544 253240 197596 253292
rect 340788 253240 340840 253292
rect 357532 253240 357584 253292
rect 357716 253240 357768 253292
rect 499212 253240 499264 253292
rect 517796 253240 517848 253292
rect 179328 253172 179380 253224
rect 197452 253172 197504 253224
rect 197636 253172 197688 253224
rect 351828 253172 351880 253224
rect 358084 253172 358136 253224
rect 517704 253172 517756 253224
rect 517980 253172 518032 253224
rect 510896 252560 510948 252612
rect 517520 252560 517572 252612
rect 214472 252492 214524 252544
rect 231124 252492 231176 252544
rect 375196 252492 375248 252544
rect 377680 252492 377732 252544
rect 396724 252492 396776 252544
rect 217968 252424 218020 252476
rect 232504 252424 232556 252476
rect 368388 252424 368440 252476
rect 376208 252424 376260 252476
rect 58624 252084 58676 252136
rect 60832 252084 60884 252136
rect 375932 252016 375984 252068
rect 376208 252016 376260 252068
rect 427084 252016 427136 252068
rect 54392 251948 54444 252000
rect 60924 251948 60976 252000
rect 369676 251948 369728 252000
rect 372528 251948 372580 252000
rect 425704 251948 425756 252000
rect 54484 251880 54536 251932
rect 61108 251880 61160 251932
rect 372344 251880 372396 251932
rect 373540 251880 373592 251932
rect 429200 251880 429252 251932
rect 52460 251812 52512 251864
rect 106924 251812 106976 251864
rect 214840 251812 214892 251864
rect 229100 251812 229152 251864
rect 375196 251812 375248 251864
rect 431960 251812 432012 251864
rect 58716 251744 58768 251796
rect 61016 251744 61068 251796
rect 56968 251336 57020 251388
rect 62120 251336 62172 251388
rect 46848 251132 46900 251184
rect 52460 251132 52512 251184
rect 53012 251132 53064 251184
rect 372436 251132 372488 251184
rect 374552 251132 374604 251184
rect 375196 251132 375248 251184
rect 519084 183540 519136 183592
rect 520188 183540 520240 183592
rect 580264 183540 580316 183592
rect 520096 183472 520148 183524
rect 580356 183472 580408 183524
rect 216864 178168 216916 178220
rect 204904 177964 204956 178016
rect 216772 177964 216824 178016
rect 216864 177964 216916 178016
rect 365260 177964 365312 178016
rect 376944 177964 376996 178016
rect 202880 176604 202932 176656
rect 216680 176604 216732 176656
rect 202144 176128 202196 176180
rect 202880 176128 202932 176180
rect 358084 175924 358136 175976
rect 376944 175924 376996 175976
rect 43996 175176 44048 175228
rect 57060 175176 57112 175228
rect 207756 175176 207808 175228
rect 217048 175176 217100 175228
rect 365076 175176 365128 175228
rect 376944 175176 376996 175228
rect 216772 175108 216824 175160
rect 216956 175108 217008 175160
rect 49424 166948 49476 167000
rect 98460 166948 98512 167000
rect 197452 166948 197504 167000
rect 201592 166948 201644 167000
rect 373264 166948 373316 167000
rect 421012 166948 421064 167000
rect 50804 166880 50856 166932
rect 101036 166880 101088 166932
rect 362408 166880 362460 166932
rect 423404 166880 423456 166932
rect 52000 166812 52052 166864
rect 105820 166812 105872 166864
rect 358268 166812 358320 166864
rect 418436 166812 418488 166864
rect 53564 166744 53616 166796
rect 108212 166744 108264 166796
rect 210884 166744 210936 166796
rect 220820 166744 220872 166796
rect 363972 166744 364024 166796
rect 428188 166744 428240 166796
rect 56416 166676 56468 166728
rect 138480 166676 138532 166728
rect 214656 166676 214708 166728
rect 260932 166676 260984 166728
rect 356796 166676 356848 166728
rect 445852 166676 445904 166728
rect 58992 166608 59044 166660
rect 140872 166608 140924 166660
rect 203616 166608 203668 166660
rect 265900 166608 265952 166660
rect 372068 166608 372120 166660
rect 470968 166608 471020 166660
rect 60004 166540 60056 166592
rect 145932 166540 145984 166592
rect 210608 166540 210660 166592
rect 293408 166540 293460 166592
rect 373448 166540 373500 166592
rect 475844 166540 475896 166592
rect 59084 166472 59136 166524
rect 148508 166472 148560 166524
rect 203524 166472 203576 166524
rect 285956 166472 286008 166524
rect 367928 166472 367980 166524
rect 478420 166472 478472 166524
rect 58900 166404 58952 166456
rect 153292 166404 153344 166456
rect 203708 166404 203760 166456
rect 288256 166404 288308 166456
rect 365168 166404 365220 166456
rect 480904 166404 480956 166456
rect 43904 166336 43956 166388
rect 163320 166336 163372 166388
rect 209136 166336 209188 166388
rect 295892 166336 295944 166388
rect 369308 166336 369360 166388
rect 485964 166336 486016 166388
rect 42524 166268 42576 166320
rect 165896 166268 165948 166320
rect 202236 166268 202288 166320
rect 303528 166268 303580 166320
rect 366548 166268 366600 166320
rect 483388 166268 483440 166320
rect 50620 166200 50672 166252
rect 96068 166200 96120 166252
rect 517612 165860 517664 165912
rect 517980 165860 518032 165912
rect 53012 165656 53064 165708
rect 114376 165656 114428 165708
rect 54024 165588 54076 165640
rect 54392 165588 54444 165640
rect 116952 165588 117004 165640
rect 357440 165588 357492 165640
rect 360200 165588 360252 165640
rect 375840 165588 375892 165640
rect 436100 165588 436152 165640
rect 56508 165520 56560 165572
rect 132500 165520 132552 165572
rect 214748 165520 214800 165572
rect 300860 165520 300912 165572
rect 362500 165520 362552 165572
rect 455420 165520 455472 165572
rect 517612 165520 517664 165572
rect 517888 165520 517940 165572
rect 55036 165452 55088 165504
rect 129740 165452 129792 165504
rect 214564 165452 214616 165504
rect 280252 165452 280304 165504
rect 369216 165452 369268 165504
rect 458364 165452 458416 165504
rect 56324 165384 56376 165436
rect 128360 165384 128412 165436
rect 211896 165384 211948 165436
rect 277400 165384 277452 165436
rect 360936 165384 360988 165436
rect 443000 165384 443052 165436
rect 55128 165316 55180 165368
rect 125876 165316 125928 165368
rect 218796 165316 218848 165368
rect 283380 165316 283432 165368
rect 370596 165316 370648 165368
rect 452660 165316 452712 165368
rect 53472 165248 53524 165300
rect 120908 165248 120960 165300
rect 207664 165248 207716 165300
rect 267740 165248 267792 165300
rect 371976 165248 372028 165300
rect 449900 165248 449952 165300
rect 56232 165180 56284 165232
rect 123484 165180 123536 165232
rect 183284 165180 183336 165232
rect 197360 165180 197412 165232
rect 216036 165180 216088 165232
rect 273444 165180 273496 165232
rect 373356 165180 373408 165232
rect 447324 165180 447376 165232
rect 54944 165112 54996 165164
rect 118332 165112 118384 165164
rect 218980 165112 219032 165164
rect 276204 165112 276256 165164
rect 370504 165112 370556 165164
rect 438032 165112 438084 165164
rect 53380 165044 53432 165096
rect 113548 165044 113600 165096
rect 183376 165044 183428 165096
rect 197452 165044 197504 165096
rect 215944 165044 215996 165096
rect 258080 165044 258132 165096
rect 367836 165044 367888 165096
rect 419264 165044 419316 165096
rect 503260 165044 503312 165096
rect 517980 165044 518032 165096
rect 56140 164976 56192 165028
rect 115940 164976 115992 165028
rect 211804 164976 211856 165028
rect 252560 164976 252612 165028
rect 343456 164976 343508 165028
rect 356888 164976 356940 165028
rect 374828 164976 374880 165028
rect 440332 164976 440384 165028
rect 52092 164908 52144 164960
rect 103520 164908 103572 164960
rect 114560 164908 114612 164960
rect 196716 164908 196768 164960
rect 210516 164908 210568 164960
rect 249800 164908 249852 164960
rect 369400 164908 369452 164960
rect 434720 164908 434772 164960
rect 503352 164908 503404 164960
rect 50712 164840 50764 164892
rect 89996 164840 90048 164892
rect 113180 164840 113232 164892
rect 196624 164840 196676 164892
rect 218888 164840 218940 164892
rect 247684 164840 247736 164892
rect 343548 164840 343600 164892
rect 357440 164840 357492 164892
rect 357624 164840 357676 164892
rect 363880 164840 363932 164892
rect 409880 164840 409932 164892
rect 419264 164840 419316 164892
rect 433340 164840 433392 164892
rect 510528 164908 510580 164960
rect 517520 164908 517572 164960
rect 517612 164840 517664 164892
rect 52184 164772 52236 164824
rect 88340 164772 88392 164824
rect 115940 164772 115992 164824
rect 197728 164772 197780 164824
rect 366456 164772 366508 164824
rect 407120 164772 407172 164824
rect 428924 164772 428976 164824
rect 433432 164772 433484 164824
rect 374736 164704 374788 164756
rect 412640 164704 412692 164756
rect 378876 164636 378928 164688
rect 416044 164636 416096 164688
rect 98644 164432 98696 164484
rect 100760 164432 100812 164484
rect 83464 164364 83516 164416
rect 107660 164364 107712 164416
rect 87604 164296 87656 164348
rect 106280 164296 106332 164348
rect 49056 164160 49108 164212
rect 50896 164160 50948 164212
rect 58624 164160 58676 164212
rect 60004 164160 60056 164212
rect 46388 164092 46440 164144
rect 50804 164092 50856 164144
rect 58164 164024 58216 164076
rect 117964 164160 118016 164212
rect 211988 164160 212040 164212
rect 323308 164160 323360 164212
rect 361028 164160 361080 164212
rect 430580 164160 430632 164212
rect 56968 163956 57020 164008
rect 59360 163956 59412 164008
rect 53656 163888 53708 163940
rect 110880 164092 110932 164144
rect 219624 164092 219676 164144
rect 264980 164092 265032 164144
rect 374276 164092 374328 164144
rect 374920 164092 374972 164144
rect 434812 164092 434864 164144
rect 213184 164024 213236 164076
rect 236000 164024 236052 164076
rect 374552 164024 374604 164076
rect 431960 164024 432012 164076
rect 216220 163956 216272 164008
rect 236092 163956 236144 164008
rect 379704 163956 379756 164008
rect 426532 163956 426584 164008
rect 375012 163888 375064 163940
rect 396172 163888 396224 163940
rect 51540 163820 51592 163872
rect 56876 163820 56928 163872
rect 95240 163820 95292 163872
rect 375748 163820 375800 163872
rect 396080 163820 396132 163872
rect 52920 163752 52972 163804
rect 56508 163752 56560 163804
rect 96620 163752 96672 163804
rect 60004 163684 60056 163736
rect 106372 163684 106424 163736
rect 50896 163616 50948 163668
rect 109500 163616 109552 163668
rect 59360 163548 59412 163600
rect 118976 163548 119028 163600
rect 373540 163548 373592 163600
rect 375196 163548 375248 163600
rect 429292 163548 429344 163600
rect 50804 163480 50856 163532
rect 111156 163480 111208 163532
rect 216680 163480 216732 163532
rect 218980 163480 219032 163532
rect 263784 163480 263836 163532
rect 373080 163480 373132 163532
rect 375104 163480 375156 163532
rect 430672 163480 430724 163532
rect 57152 162800 57204 162852
rect 59084 162800 59136 162852
rect 214288 162800 214340 162852
rect 214472 162800 214524 162852
rect 214840 162800 214892 162852
rect 260840 162800 260892 162852
rect 376484 162800 376536 162852
rect 379612 162800 379664 162852
rect 379980 162800 380032 162852
rect 428924 162800 428976 162852
rect 259552 162732 259604 162784
rect 376760 162732 376812 162784
rect 420920 162732 420972 162784
rect 217968 162664 218020 162716
rect 259460 162664 259512 162716
rect 376208 162664 376260 162716
rect 418528 162664 418580 162716
rect 218520 162596 218572 162648
rect 218888 162596 218940 162648
rect 258080 162596 258132 162648
rect 375748 162596 375800 162648
rect 378692 162596 378744 162648
rect 419540 162596 419592 162648
rect 375288 162528 375340 162580
rect 379980 162528 380032 162580
rect 374368 162460 374420 162512
rect 378968 162460 379020 162512
rect 59084 162120 59136 162172
rect 89904 162120 89956 162172
rect 218612 162120 218664 162172
rect 219532 162120 219584 162172
rect 266360 162120 266412 162172
rect 379612 162120 379664 162172
rect 418160 162120 418212 162172
rect 376300 161848 376352 161900
rect 376760 161848 376812 161900
rect 216128 161576 216180 161628
rect 235264 161508 235316 161560
rect 217140 161440 217192 161492
rect 236644 161440 236696 161492
rect 378968 161440 379020 161492
rect 396724 161440 396776 161492
rect 58072 148996 58124 149048
rect 106280 148996 106332 149048
rect 213276 148996 213328 149048
rect 276112 148996 276164 149048
rect 379060 148996 379112 149048
rect 440240 148996 440292 149048
rect 58716 148928 58768 148980
rect 103520 148928 103572 148980
rect 213460 148928 213512 148980
rect 274732 148928 274784 148980
rect 373816 148928 373868 148980
rect 434720 148928 434772 148980
rect 216312 148860 216364 148912
rect 277400 148860 277452 148912
rect 379796 148860 379848 148912
rect 427820 148860 427872 148912
rect 46664 148792 46716 148844
rect 59912 148792 59964 148844
rect 83464 148792 83516 148844
rect 214932 148792 214984 148844
rect 274640 148792 274692 148844
rect 373724 148792 373776 148844
rect 397460 148792 397512 148844
rect 48044 148724 48096 148776
rect 55036 148724 55088 148776
rect 80060 148724 80112 148776
rect 213552 148724 213604 148776
rect 241520 148724 241572 148776
rect 46480 148656 46532 148708
rect 58992 148656 59044 148708
rect 87604 148656 87656 148708
rect 49148 148588 49200 148640
rect 52184 148588 52236 148640
rect 81440 148588 81492 148640
rect 54484 148520 54536 148572
rect 56232 148520 56284 148572
rect 102140 148520 102192 148572
rect 213736 148520 213788 148572
rect 238760 148520 238812 148572
rect 372252 148520 372304 148572
rect 374736 148520 374788 148572
rect 400220 148520 400272 148572
rect 53472 148452 53524 148504
rect 113180 148452 113232 148504
rect 215024 148452 215076 148504
rect 240140 148452 240192 148504
rect 370780 148452 370832 148504
rect 373264 148452 373316 148504
rect 398840 148452 398892 148504
rect 53564 148384 53616 148436
rect 114560 148384 114612 148436
rect 212172 148384 212224 148436
rect 214656 148384 214708 148436
rect 270500 148384 270552 148436
rect 370964 148384 371016 148436
rect 373356 148384 373408 148436
rect 401600 148384 401652 148436
rect 53380 148316 53432 148368
rect 115940 148316 115992 148368
rect 215760 148316 215812 148368
rect 271880 148316 271932 148368
rect 372528 148316 372580 148368
rect 379980 148316 380032 148368
rect 429200 148316 429252 148368
rect 56324 147636 56376 147688
rect 58716 147636 58768 147688
rect 213368 147636 213420 147688
rect 214932 147636 214984 147688
rect 379336 147636 379388 147688
rect 379796 147636 379848 147688
rect 206744 147568 206796 147620
rect 213184 147568 213236 147620
rect 213736 147568 213788 147620
rect 212264 147500 212316 147552
rect 215760 147500 215812 147552
rect 215944 147500 215996 147552
rect 213276 147432 213328 147484
rect 213736 147432 213788 147484
rect 210976 147364 211028 147416
rect 214564 147364 214616 147416
rect 215024 147364 215076 147416
rect 215024 146276 215076 146328
rect 276020 146276 276072 146328
rect 46296 146208 46348 146260
rect 52092 146208 52144 146260
rect 57060 146208 57112 146260
rect 57980 146208 58032 146260
rect 59820 146208 59872 146260
rect 93860 146208 93912 146260
rect 179052 146208 179104 146260
rect 197636 146208 197688 146260
rect 236644 146208 236696 146260
rect 256700 146208 256752 146260
rect 356612 146208 356664 146260
rect 375932 146208 375984 146260
rect 377956 146208 378008 146260
rect 378600 146208 378652 146260
rect 379244 146208 379296 146260
rect 379888 146208 379940 146260
rect 414020 146208 414072 146260
rect 91192 146140 91244 146192
rect 179696 146140 179748 146192
rect 197544 146140 197596 146192
rect 235264 146140 235316 146192
rect 255320 146140 255372 146192
rect 338488 146140 338540 146192
rect 357808 146140 357860 146192
rect 378416 146140 378468 146192
rect 379428 146140 379480 146192
rect 396724 146140 396776 146192
rect 416780 146140 416832 146192
rect 500224 146140 500276 146192
rect 517704 146140 517756 146192
rect 55956 146072 56008 146124
rect 88432 146072 88484 146124
rect 215852 146072 215904 146124
rect 219348 146072 219400 146124
rect 252560 146072 252612 146124
rect 340236 146072 340288 146124
rect 357716 146072 357768 146124
rect 379060 146072 379112 146124
rect 379520 146072 379572 146124
rect 412732 146072 412784 146124
rect 498660 146072 498712 146124
rect 517520 146072 517572 146124
rect 517796 146072 517848 146124
rect 53656 146004 53708 146056
rect 54116 146004 54168 146056
rect 86960 146004 87012 146056
rect 216496 146004 216548 146056
rect 249800 146004 249852 146056
rect 379428 146004 379480 146056
rect 411352 146004 411404 146056
rect 54300 145936 54352 145988
rect 54852 145936 54904 145988
rect 82820 145936 82872 145988
rect 219164 145936 219216 145988
rect 251180 145936 251232 145988
rect 377312 145936 377364 145988
rect 379152 145936 379204 145988
rect 409880 145936 409932 145988
rect 58808 145868 58860 145920
rect 84200 145868 84252 145920
rect 216128 145868 216180 145920
rect 217324 145868 217376 145920
rect 247040 145868 247092 145920
rect 377956 145868 378008 145920
rect 408500 145868 408552 145920
rect 47860 145800 47912 145852
rect 53104 145800 53156 145852
rect 78680 145800 78732 145852
rect 216404 145800 216456 145852
rect 242900 145800 242952 145852
rect 375840 145800 375892 145852
rect 376576 145800 376628 145852
rect 376668 145800 376720 145852
rect 404360 145800 404412 145852
rect 56416 145732 56468 145784
rect 84292 145732 84344 145784
rect 214932 145732 214984 145784
rect 219072 145732 219124 145784
rect 244372 145732 244424 145784
rect 403072 145732 403124 145784
rect 53840 145664 53892 145716
rect 85580 145664 85632 145716
rect 218060 145664 218112 145716
rect 245660 145664 245712 145716
rect 375012 145664 375064 145716
rect 402980 145664 403032 145716
rect 58624 145596 58676 145648
rect 91100 145596 91152 145648
rect 216036 145596 216088 145648
rect 244280 145596 244332 145648
rect 280068 145596 280120 145648
rect 356612 145596 356664 145648
rect 357532 145596 357584 145648
rect 376116 145596 376168 145648
rect 407212 145596 407264 145648
rect 517520 145596 517572 145648
rect 580356 145596 580408 145648
rect 53932 145528 53984 145580
rect 98000 145528 98052 145580
rect 191288 145528 191340 145580
rect 202144 145528 202196 145580
rect 204904 145528 204956 145580
rect 217048 145528 217100 145580
rect 248420 145528 248472 145580
rect 351644 145528 351696 145580
rect 358084 145528 358136 145580
rect 358728 145528 358780 145580
rect 510528 145528 510580 145580
rect 517704 145528 517756 145580
rect 580264 145528 580316 145580
rect 52092 145460 52144 145512
rect 77300 145460 77352 145512
rect 218520 145460 218572 145512
rect 236092 145460 236144 145512
rect 379244 145460 379296 145512
rect 405740 145460 405792 145512
rect 47952 145392 48004 145444
rect 54392 145392 54444 145444
rect 76012 145392 76064 145444
rect 218612 145392 218664 145444
rect 236000 145392 236052 145444
rect 378692 145392 378744 145444
rect 396172 145392 396224 145444
rect 46572 145324 46624 145376
rect 54944 145324 54996 145376
rect 75920 145324 75972 145376
rect 219808 145324 219860 145376
rect 253940 145324 253992 145376
rect 378784 145324 378836 145376
rect 396080 145324 396132 145376
rect 216772 145256 216824 145308
rect 217232 145256 217284 145308
rect 251272 145256 251324 145308
rect 378048 145256 378100 145308
rect 411260 145256 411312 145308
rect 51724 144848 51776 144900
rect 53840 144848 53892 144900
rect 54484 144848 54536 144900
rect 54576 144848 54628 144900
rect 58808 144848 58860 144900
rect 209504 144848 209556 144900
rect 213276 144848 213328 144900
rect 214380 144848 214432 144900
rect 217048 144848 217100 144900
rect 373632 144848 373684 144900
rect 374828 144848 374880 144900
rect 375012 144848 375064 144900
rect 51816 144780 51868 144832
rect 58624 144780 58676 144832
rect 213644 144780 213696 144832
rect 214472 144780 214524 144832
rect 374460 144780 374512 144832
rect 376116 144780 376168 144832
rect 50436 144712 50488 144764
rect 53932 144712 53984 144764
rect 54668 144712 54720 144764
rect 213092 144712 213144 144764
rect 216036 144712 216088 144764
rect 50528 144644 50580 144696
rect 55864 144644 55916 144696
rect 56416 144644 56468 144696
rect 212356 144644 212408 144696
rect 218060 144644 218112 144696
rect 218796 144644 218848 144696
rect 49240 144576 49292 144628
rect 58716 144576 58768 144628
rect 53196 144508 53248 144560
rect 58900 144508 58952 144560
rect 55956 144372 56008 144424
rect 56324 144372 56376 144424
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 42616 70320 42668 70372
rect 57612 70320 57664 70372
rect 209044 70320 209096 70372
rect 216680 70320 216732 70372
rect 362316 70320 362368 70372
rect 376944 70320 376996 70372
rect 358728 68280 358780 68332
rect 376944 68280 376996 68332
rect 358084 68144 358136 68196
rect 358728 68144 358780 68196
rect 204904 67600 204956 67652
rect 216680 67600 216732 67652
rect 218612 61208 218664 61260
rect 219072 61208 219124 61260
rect 54392 59644 54444 59696
rect 77116 59644 77168 59696
rect 218520 59644 218572 59696
rect 237104 59644 237156 59696
rect 378784 59644 378836 59696
rect 396080 59644 396132 59696
rect 54852 59576 54904 59628
rect 83096 59576 83148 59628
rect 216956 59576 217008 59628
rect 256976 59576 257028 59628
rect 378692 59576 378744 59628
rect 397092 59576 397144 59628
rect 58900 59508 58952 59560
rect 100760 59508 100812 59560
rect 216220 59508 216272 59560
rect 255872 59508 255924 59560
rect 378968 59508 379020 59560
rect 416964 59508 417016 59560
rect 54760 59440 54812 59492
rect 101772 59440 101824 59492
rect 218980 59440 219032 59492
rect 263876 59440 263928 59492
rect 377496 59440 377548 59492
rect 423956 59440 424008 59492
rect 49516 59372 49568 59424
rect 113548 59372 113600 59424
rect 215852 59372 215904 59424
rect 262864 59372 262916 59424
rect 358176 59372 358228 59424
rect 423496 59372 423548 59424
rect 55864 59304 55916 59356
rect 84200 59304 84252 59356
rect 217968 59304 218020 59356
rect 358084 59304 358136 59356
rect 379612 59304 379664 59356
rect 418160 59304 418212 59356
rect 59084 59236 59136 59288
rect 89996 59236 90048 59288
rect 218888 59236 218940 59288
rect 258080 59236 258132 59288
rect 371884 59236 371936 59288
rect 410708 59236 410760 59288
rect 59820 59168 59872 59220
rect 94504 59168 94556 59220
rect 214288 59168 214340 59220
rect 260656 59168 260708 59220
rect 376208 59168 376260 59220
rect 419448 59168 419500 59220
rect 56876 59100 56928 59152
rect 95884 59100 95936 59152
rect 214748 59100 214800 59152
rect 261760 59100 261812 59152
rect 279240 59100 279292 59152
rect 356612 59100 356664 59152
rect 375748 59100 375800 59152
rect 420644 59100 420696 59152
rect 56508 59032 56560 59084
rect 96988 59032 97040 59084
rect 205180 59032 205232 59084
rect 290924 59032 290976 59084
rect 376300 59032 376352 59084
rect 421748 59032 421800 59084
rect 54668 58964 54720 59016
rect 98092 58964 98144 59016
rect 213828 58964 213880 59016
rect 300860 58964 300912 59016
rect 360844 58964 360896 59016
rect 416044 58964 416096 59016
rect 56232 58896 56284 58948
rect 102784 58896 102836 58948
rect 212448 58896 212500 58948
rect 315856 58896 315908 58948
rect 356704 58896 356756 58948
rect 425980 58896 426032 58948
rect 58992 58828 59044 58880
rect 107568 58828 107620 58880
rect 202788 58828 202840 58880
rect 308496 58828 308548 58880
rect 369124 58828 369176 58880
rect 458456 58828 458508 58880
rect 48780 58760 48832 58812
rect 110972 58760 111024 58812
rect 206928 58760 206980 58812
rect 320916 58760 320968 58812
rect 362224 58760 362276 58812
rect 453396 58760 453448 58812
rect 53288 58692 53340 58744
rect 148508 58692 148560 58744
rect 205364 58692 205416 58744
rect 325884 58692 325936 58744
rect 364984 58692 365036 58744
rect 475844 58692 475896 58744
rect 50988 58624 51040 58676
rect 150900 58624 150952 58676
rect 219256 58624 219308 58676
rect 428188 58624 428240 58676
rect 374828 58556 374880 58608
rect 404176 58556 404228 58608
rect 375840 58420 375892 58472
rect 403072 58420 403124 58472
rect 57888 57876 57940 57928
rect 204904 57876 204956 57928
rect 210240 57876 210292 57928
rect 323308 57876 323360 57928
rect 343180 57876 343232 57928
rect 357624 57876 357676 57928
rect 376668 57876 376720 57928
rect 485964 57876 486016 57928
rect 503352 57876 503404 57928
rect 517612 57876 517664 57928
rect 52368 57808 52420 57860
rect 145564 57808 145616 57860
rect 183468 57808 183520 57860
rect 197452 57808 197504 57860
rect 208308 57808 208360 57860
rect 313372 57808 313424 57860
rect 343456 57808 343508 57860
rect 356796 57808 356848 57860
rect 366364 57808 366416 57860
rect 470876 57808 470928 57860
rect 503260 57808 503312 57860
rect 517980 57808 518032 57860
rect 53748 57740 53800 57792
rect 133420 57740 133472 57792
rect 183192 57740 183244 57792
rect 197360 57740 197412 57792
rect 218704 57740 218756 57792
rect 318248 57740 318300 57792
rect 361488 57740 361540 57792
rect 465908 57740 465960 57792
rect 52276 57672 52328 57724
rect 130844 57672 130896 57724
rect 215116 57672 215168 57724
rect 310980 57672 311032 57724
rect 378508 57672 378560 57724
rect 478420 57672 478472 57724
rect 42708 57604 42760 57656
rect 115940 57604 115992 57656
rect 216588 57604 216640 57656
rect 305828 57604 305880 57656
rect 371148 57604 371200 57656
rect 460940 57604 460992 57656
rect 56416 57536 56468 57588
rect 103796 57536 103848 57588
rect 215208 57536 215260 57588
rect 303436 57536 303488 57588
rect 363788 57536 363840 57588
rect 451004 57536 451056 57588
rect 56140 57468 56192 57520
rect 99380 57468 99432 57520
rect 208860 57468 208912 57520
rect 295892 57468 295944 57520
rect 363696 57468 363748 57520
rect 445852 57468 445904 57520
rect 51448 57400 51500 57452
rect 88340 57400 88392 57452
rect 218428 57400 218480 57452
rect 298100 57400 298152 57452
rect 363604 57400 363656 57452
rect 430948 57400 431000 57452
rect 59268 57332 59320 57384
rect 93676 57332 93728 57384
rect 205548 57332 205600 57384
rect 278320 57332 278372 57384
rect 367744 57332 367796 57384
rect 435916 57332 435968 57384
rect 59176 57264 59228 57316
rect 90732 57264 90784 57316
rect 218612 57264 218664 57316
rect 258356 57264 258408 57316
rect 374644 57264 374696 57316
rect 438492 57264 438544 57316
rect 52092 57196 52144 57248
rect 78220 57196 78272 57248
rect 210424 57196 210476 57248
rect 248236 57196 248288 57248
rect 378876 57196 378928 57248
rect 415492 57196 415544 57248
rect 57244 57128 57296 57180
rect 57888 57128 57940 57180
rect 54944 57060 54996 57112
rect 76012 57128 76064 57180
rect 53380 56516 53432 56568
rect 115756 56516 115808 56568
rect 219992 56516 220044 56568
rect 408316 56516 408368 56568
rect 50804 56448 50856 56500
rect 111156 56448 111208 56500
rect 215024 56448 215076 56500
rect 276940 56448 276992 56500
rect 375656 56448 375708 56500
rect 436284 56448 436336 56500
rect 53472 56380 53524 56432
rect 112076 56380 112128 56432
rect 219072 56380 219124 56432
rect 236000 56380 236052 56432
rect 375288 56380 375340 56432
rect 434444 56380 434496 56432
rect 59912 56312 59964 56364
rect 108212 56312 108264 56364
rect 213368 56312 213420 56364
rect 273260 56312 273312 56364
rect 374552 56312 374604 56364
rect 432236 56312 432288 56364
rect 58716 56244 58768 56296
rect 93308 56244 93360 56296
rect 214656 56244 214708 56296
rect 271052 56244 271104 56296
rect 379336 56244 379388 56296
rect 427636 56244 427688 56296
rect 56324 56176 56376 56228
rect 88708 56176 88760 56228
rect 219900 56176 219952 56228
rect 268108 56176 268160 56228
rect 379888 56176 379940 56228
rect 414572 56176 414624 56228
rect 54484 56108 54536 56160
rect 86500 56108 86552 56160
rect 218244 56108 218296 56160
rect 266360 56108 266412 56160
rect 379060 56108 379112 56160
rect 412640 56108 412692 56160
rect 58808 56040 58860 56092
rect 85396 56040 85448 56092
rect 219348 56040 219400 56092
rect 253388 56040 253440 56092
rect 375932 56040 375984 56092
rect 408684 56040 408736 56092
rect 55036 55972 55088 56024
rect 80428 55972 80480 56024
rect 219164 55972 219216 56024
rect 251180 55972 251232 56024
rect 379428 55972 379480 56024
rect 411260 55972 411312 56024
rect 217140 55904 217192 55956
rect 248604 55904 248656 55956
rect 373356 55904 373408 55956
rect 401692 55904 401744 55956
rect 213552 55836 213604 55888
rect 241612 55836 241664 55888
rect 373264 55836 373316 55888
rect 399484 55836 399536 55888
rect 216036 55768 216088 55820
rect 245292 55768 245344 55820
rect 213184 55700 213236 55752
rect 239220 55700 239272 55752
rect 213736 55632 213788 55684
rect 275100 55632 275152 55684
rect 53104 55156 53156 55208
rect 78680 55156 78732 55208
rect 216404 55156 216456 55208
rect 242900 55156 242952 55208
rect 379244 55156 379296 55208
rect 405832 55156 405884 55208
rect 54024 55088 54076 55140
rect 116124 55088 116176 55140
rect 214564 55088 214616 55140
rect 240140 55088 240192 55140
rect 374736 55088 374788 55140
rect 400220 55088 400272 55140
rect 53564 55020 53616 55072
rect 113180 55020 113232 55072
rect 215944 55020 215996 55072
rect 271880 55020 271932 55072
rect 373816 55020 373868 55072
rect 433432 55020 433484 55072
rect 53012 54952 53064 55004
rect 113272 54952 113324 55004
rect 219532 54952 219584 55004
rect 266452 54952 266504 55004
rect 375104 54952 375156 55004
rect 430580 54952 430632 55004
rect 50896 54884 50948 54936
rect 109040 54884 109092 54936
rect 219624 54884 219676 54936
rect 264980 54884 265032 54936
rect 375196 54884 375248 54936
rect 429200 54884 429252 54936
rect 60004 54816 60056 54868
rect 106280 54816 106332 54868
rect 219808 54816 219860 54868
rect 253940 54816 253992 54868
rect 379980 54816 380032 54868
rect 427820 54816 427872 54868
rect 57060 54748 57112 54800
rect 91100 54748 91152 54800
rect 217232 54748 217284 54800
rect 251364 54748 251416 54800
rect 379704 54748 379756 54800
rect 426532 54748 426584 54800
rect 53656 54680 53708 54732
rect 86960 54680 87012 54732
rect 216496 54680 216548 54732
rect 249800 54680 249852 54732
rect 378048 54680 378100 54732
rect 411352 54680 411404 54732
rect 58624 54612 58676 54664
rect 91468 54612 91520 54664
rect 216128 54612 216180 54664
rect 247040 54612 247092 54664
rect 377312 54612 377364 54664
rect 409880 54612 409932 54664
rect 52184 54544 52236 54596
rect 81440 54544 81492 54596
rect 214932 54544 214984 54596
rect 244372 54544 244424 54596
rect 376116 54544 376168 54596
rect 407212 54544 407264 54596
rect 44088 54476 44140 54528
rect 122840 54476 122892 54528
rect 218796 54476 218848 54528
rect 245660 54476 245712 54528
rect 376484 54476 376536 54528
rect 404360 54476 404412 54528
rect 216312 54408 216364 54460
rect 277400 54408 277452 54460
rect 375564 54408 375616 54460
rect 437480 54408 437532 54460
rect 213460 54340 213512 54392
rect 273352 54340 273404 54392
rect 374276 54340 374328 54392
rect 434720 54340 434772 54392
rect 213276 54272 213328 54324
rect 237380 54272 237432 54324
rect 373724 54272 373776 54324
rect 397460 54272 397512 54324
rect 3424 20612 3476 20664
rect 10324 20612 10376 20664
rect 572 3408 624 3460
rect 57244 3408 57296 3460
rect 125876 2796 125928 2848
rect 365720 2796 365772 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 639736 3476 639742
rect 3424 639678 3476 639684
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3436 201929 3464 639678
rect 3528 638246 3556 684247
rect 3608 639668 3660 639674
rect 3608 639610 3660 639616
rect 3516 638240 3568 638246
rect 3516 638182 3568 638188
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3528 573374 3556 632023
rect 3516 573368 3568 573374
rect 3516 573310 3568 573316
rect 3514 548040 3570 548049
rect 3514 547975 3570 547984
rect 3528 514865 3556 547975
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3514 482216 3570 482225
rect 3514 482151 3570 482160
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3528 58585 3556 482151
rect 3620 306241 3648 639610
rect 3700 639600 3752 639606
rect 3700 639542 3752 639548
rect 3712 358465 3740 639542
rect 3790 580000 3846 580009
rect 3790 579935 3846 579944
rect 3804 575482 3832 579935
rect 3792 575476 3844 575482
rect 3792 575418 3844 575424
rect 10324 570648 10376 570654
rect 10324 570590 10376 570596
rect 4804 561740 4856 561746
rect 4804 561682 4856 561688
rect 3792 480956 3844 480962
rect 3792 480898 3844 480904
rect 3804 462641 3832 480898
rect 3790 462632 3846 462641
rect 3790 462567 3846 462576
rect 3698 358456 3754 358465
rect 3698 358391 3754 358400
rect 3606 306232 3662 306241
rect 3606 306167 3662 306176
rect 4816 97782 4844 561682
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 10336 20670 10364 570590
rect 40052 558890 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 57704 700324 57756 700330
rect 57704 700266 57756 700272
rect 54852 640552 54904 640558
rect 54852 640494 54904 640500
rect 54864 574938 54892 640494
rect 55128 640484 55180 640490
rect 55128 640426 55180 640432
rect 55036 640416 55088 640422
rect 55036 640358 55088 640364
rect 54944 637900 54996 637906
rect 54944 637842 54996 637848
rect 54852 574932 54904 574938
rect 54852 574874 54904 574880
rect 40040 558884 40092 558890
rect 40040 558826 40092 558832
rect 54956 550390 54984 637842
rect 54944 550384 54996 550390
rect 54944 550326 54996 550332
rect 55048 550118 55076 640358
rect 55140 550526 55168 640426
rect 56508 640348 56560 640354
rect 56508 640290 56560 640296
rect 56416 637832 56468 637838
rect 56416 637774 56468 637780
rect 56324 637764 56376 637770
rect 56324 637706 56376 637712
rect 55128 550520 55180 550526
rect 55128 550462 55180 550468
rect 55036 550112 55088 550118
rect 55036 550054 55088 550060
rect 56336 549982 56364 637706
rect 56428 550050 56456 637774
rect 56520 550254 56548 640290
rect 57610 635624 57666 635633
rect 57610 635559 57666 635568
rect 57518 626784 57574 626793
rect 57518 626719 57574 626728
rect 57426 605024 57482 605033
rect 57426 604959 57482 604968
rect 57242 598904 57298 598913
rect 57242 598839 57298 598848
rect 57150 596184 57206 596193
rect 57150 596119 57206 596128
rect 57058 590064 57114 590073
rect 57058 589999 57114 590008
rect 57072 575346 57100 589999
rect 57164 575754 57192 596119
rect 57152 575748 57204 575754
rect 57152 575690 57204 575696
rect 57060 575340 57112 575346
rect 57060 575282 57112 575288
rect 57256 566642 57284 598839
rect 57334 586664 57390 586673
rect 57334 586599 57390 586608
rect 57348 572082 57376 586599
rect 57440 574326 57468 604959
rect 57428 574320 57480 574326
rect 57428 574262 57480 574268
rect 57532 573510 57560 626719
rect 57520 573504 57572 573510
rect 57520 573446 57572 573452
rect 57336 572076 57388 572082
rect 57336 572018 57388 572024
rect 57244 566636 57296 566642
rect 57244 566578 57296 566584
rect 57624 555490 57652 635559
rect 57716 614553 57744 700266
rect 104912 647902 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 700398 170352 703520
rect 235184 700466 235212 703520
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 147220 683188 147272 683194
rect 147220 683130 147272 683136
rect 104900 647896 104952 647902
rect 104900 647838 104952 647844
rect 131120 641028 131172 641034
rect 131120 640970 131172 640976
rect 115388 640892 115440 640898
rect 115388 640834 115440 640840
rect 124680 640892 124732 640898
rect 124680 640834 124732 640840
rect 69020 640756 69072 640762
rect 69020 640698 69072 640704
rect 60740 640620 60792 640626
rect 60740 640562 60792 640568
rect 60752 637974 60780 640562
rect 65800 640416 65852 640422
rect 65800 640358 65852 640364
rect 65812 638044 65840 640358
rect 69032 638044 69060 640698
rect 112168 640688 112220 640694
rect 112168 640630 112220 640636
rect 98000 640620 98052 640626
rect 98000 640562 98052 640568
rect 106372 640620 106424 640626
rect 106372 640562 106424 640568
rect 88984 640552 89036 640558
rect 88984 640494 89036 640500
rect 77392 640348 77444 640354
rect 77392 640290 77444 640296
rect 77404 638044 77432 640290
rect 88996 638044 89024 640494
rect 92204 640484 92256 640490
rect 92204 640426 92256 640432
rect 94780 640484 94832 640490
rect 94780 640426 94832 640432
rect 92216 638044 92244 640426
rect 94792 638044 94820 640426
rect 98012 638044 98040 640562
rect 103796 640552 103848 640558
rect 103796 640494 103848 640500
rect 100576 640416 100628 640422
rect 100576 640358 100628 640364
rect 100588 638044 100616 640358
rect 103808 638044 103836 640494
rect 106384 638044 106412 640562
rect 109592 640348 109644 640354
rect 109592 640290 109644 640296
rect 109604 638044 109632 640290
rect 112180 638044 112208 640630
rect 115400 638044 115428 640834
rect 124404 640824 124456 640830
rect 124404 640766 124456 640772
rect 117964 640756 118016 640762
rect 117964 640698 118016 640704
rect 117976 640422 118004 640698
rect 122840 640688 122892 640694
rect 122840 640630 122892 640636
rect 121460 640620 121512 640626
rect 121460 640562 121512 640568
rect 120908 640484 120960 640490
rect 120908 640426 120960 640432
rect 117964 640416 118016 640422
rect 117964 640358 118016 640364
rect 118240 640348 118292 640354
rect 118240 640290 118292 640296
rect 118252 638058 118280 640290
rect 117990 638030 118280 638058
rect 59360 637968 59412 637974
rect 59360 637910 59412 637916
rect 60740 637968 60792 637974
rect 60740 637910 60792 637916
rect 57796 637696 57848 637702
rect 57796 637638 57848 637644
rect 57702 614544 57758 614553
rect 57702 614479 57758 614488
rect 57702 602304 57758 602313
rect 57702 602239 57758 602248
rect 57716 589286 57744 602239
rect 57704 589280 57756 589286
rect 57704 589222 57756 589228
rect 57702 580544 57758 580553
rect 57702 580479 57758 580488
rect 57612 555484 57664 555490
rect 57612 555426 57664 555432
rect 57716 552702 57744 580479
rect 57704 552696 57756 552702
rect 57704 552638 57756 552644
rect 57808 550322 57836 637638
rect 57888 637628 57940 637634
rect 57888 637570 57940 637576
rect 57900 611153 57928 637570
rect 59082 632904 59138 632913
rect 59082 632839 59138 632848
rect 58898 623384 58954 623393
rect 58898 623319 58954 623328
rect 57886 611144 57942 611153
rect 57886 611079 57942 611088
rect 57796 550316 57848 550322
rect 57796 550258 57848 550264
rect 56508 550248 56560 550254
rect 56508 550190 56560 550196
rect 56416 550044 56468 550050
rect 56416 549986 56468 549992
rect 56324 549976 56376 549982
rect 56324 549918 56376 549924
rect 57900 517993 57928 611079
rect 58806 608424 58862 608433
rect 58806 608359 58862 608368
rect 58714 592784 58770 592793
rect 58714 592719 58770 592728
rect 58624 589280 58676 589286
rect 58624 589222 58676 589228
rect 58530 583944 58586 583953
rect 58530 583879 58586 583888
rect 58544 569294 58572 583879
rect 58532 569288 58584 569294
rect 58532 569230 58584 569236
rect 58636 550186 58664 589222
rect 58728 574870 58756 592719
rect 58716 574864 58768 574870
rect 58716 574806 58768 574812
rect 58820 570790 58848 608359
rect 58912 575006 58940 623319
rect 58990 617264 59046 617273
rect 58990 617199 59046 617208
rect 58900 575000 58952 575006
rect 58900 574942 58952 574948
rect 58808 570784 58860 570790
rect 58808 570726 58860 570732
rect 59004 562358 59032 617199
rect 59096 573578 59124 632839
rect 59266 629504 59322 629513
rect 59266 629439 59322 629448
rect 59174 620664 59230 620673
rect 59174 620599 59230 620608
rect 59084 573572 59136 573578
rect 59084 573514 59136 573520
rect 58992 562352 59044 562358
rect 58992 562294 59044 562300
rect 59188 559570 59216 620599
rect 59280 560998 59308 629439
rect 59268 560992 59320 560998
rect 59268 560934 59320 560940
rect 59176 559564 59228 559570
rect 59176 559506 59228 559512
rect 59372 552786 59400 637910
rect 62960 637906 63250 637922
rect 62948 637900 63250 637906
rect 63000 637894 63250 637900
rect 62948 637842 63000 637848
rect 71228 637832 71280 637838
rect 86776 637832 86828 637838
rect 71280 637780 71622 637786
rect 71228 637774 71622 637780
rect 71240 637758 71622 637774
rect 74644 637770 74842 637786
rect 74632 637764 74842 637770
rect 74684 637758 74842 637764
rect 86434 637780 86776 637786
rect 86434 637774 86828 637780
rect 86434 637758 86816 637774
rect 74632 637706 74684 637712
rect 80244 637696 80296 637702
rect 83464 637696 83516 637702
rect 80296 637644 80638 637650
rect 80244 637638 80638 637644
rect 80256 637622 80638 637638
rect 83214 637644 83464 637650
rect 83214 637638 83516 637644
rect 83214 637622 83504 637638
rect 59464 637350 60030 637378
rect 120566 637350 120764 637378
rect 59464 568002 59492 637350
rect 120736 581670 120764 637350
rect 120814 613320 120870 613329
rect 120814 613255 120870 613264
rect 120724 581664 120776 581670
rect 120724 581606 120776 581612
rect 59542 577788 59598 577797
rect 59542 577723 59598 577732
rect 59452 567996 59504 568002
rect 59452 567938 59504 567944
rect 59556 563786 59584 577723
rect 120722 576872 120778 576881
rect 120722 576807 120778 576816
rect 59912 575748 59964 575754
rect 59912 575690 59964 575696
rect 59544 563780 59596 563786
rect 59544 563722 59596 563728
rect 59924 557534 59952 575690
rect 62120 575340 62172 575346
rect 62120 575282 62172 575288
rect 106280 575340 106332 575346
rect 106280 575282 106332 575288
rect 60016 572014 60044 575076
rect 60740 574320 60792 574326
rect 60740 574262 60792 574268
rect 60004 572008 60056 572014
rect 60004 571950 60056 571956
rect 60752 557534 60780 574262
rect 59924 557506 60412 557534
rect 60752 557506 60964 557534
rect 59372 552758 60320 552786
rect 58624 550180 58676 550186
rect 58624 550122 58676 550128
rect 60292 547963 60320 552758
rect 60384 549914 60412 557506
rect 60372 549908 60424 549914
rect 60372 549850 60424 549856
rect 60936 547963 60964 557506
rect 62132 552786 62160 575282
rect 99564 575272 99616 575278
rect 99564 575214 99616 575220
rect 98092 575204 98144 575210
rect 98092 575146 98144 575152
rect 96804 575136 96856 575142
rect 62224 575062 62606 575090
rect 62224 556918 62252 575062
rect 63500 574796 63552 574802
rect 63500 574738 63552 574744
rect 62764 572552 62816 572558
rect 62764 572494 62816 572500
rect 62212 556912 62264 556918
rect 62212 556854 62264 556860
rect 62132 552758 62436 552786
rect 61660 550588 61712 550594
rect 61660 550530 61712 550536
rect 61672 547963 61700 550530
rect 62408 547963 62436 552758
rect 62776 550594 62804 572494
rect 63132 554056 63184 554062
rect 63132 553998 63184 554004
rect 62764 550588 62816 550594
rect 62764 550530 62816 550536
rect 63144 547963 63172 553998
rect 63512 552786 63540 574738
rect 65064 573436 65116 573442
rect 65064 573378 65116 573384
rect 63592 566500 63644 566506
rect 63592 566442 63644 566448
rect 63604 557534 63632 566442
rect 64972 565140 65024 565146
rect 64972 565082 65024 565088
rect 63604 557506 64552 557534
rect 63512 552758 63816 552786
rect 63788 547963 63816 552758
rect 64524 547963 64552 557506
rect 64984 552770 65012 565082
rect 65076 557534 65104 573378
rect 65168 572558 65196 575076
rect 67836 575062 68402 575090
rect 67640 574864 67692 574870
rect 67640 574806 67692 574812
rect 65156 572552 65208 572558
rect 65156 572494 65208 572500
rect 66352 570716 66404 570722
rect 66352 570658 66404 570664
rect 66364 557534 66392 570658
rect 65076 557506 65288 557534
rect 66364 557506 66760 557534
rect 64972 552764 65024 552770
rect 64972 552706 65024 552712
rect 65260 547963 65288 557506
rect 65984 552764 66036 552770
rect 65984 552706 66036 552712
rect 65996 547963 66024 552706
rect 66732 547963 66760 557506
rect 67652 552770 67680 574806
rect 67732 569220 67784 569226
rect 67732 569162 67784 569168
rect 67744 557534 67772 569162
rect 67836 558210 67864 575062
rect 69020 574864 69072 574870
rect 69020 574806 69072 574812
rect 67824 558204 67876 558210
rect 67824 558146 67876 558152
rect 67744 557506 68140 557534
rect 67640 552764 67692 552770
rect 67640 552706 67692 552712
rect 67364 550520 67416 550526
rect 67364 550462 67416 550468
rect 67376 547963 67404 550462
rect 68112 547963 68140 557506
rect 69032 552770 69060 574806
rect 70964 572218 70992 575076
rect 70952 572212 71004 572218
rect 70952 572154 71004 572160
rect 71044 572008 71096 572014
rect 71044 571950 71096 571956
rect 69112 567928 69164 567934
rect 69112 567870 69164 567876
rect 69124 557534 69152 567870
rect 70400 567860 70452 567866
rect 70400 567802 70452 567808
rect 70412 557534 70440 567802
rect 69124 557506 69612 557534
rect 70412 557506 70992 557534
rect 68836 552764 68888 552770
rect 68836 552706 68888 552712
rect 69020 552764 69072 552770
rect 69020 552706 69072 552712
rect 68848 547963 68876 552706
rect 69584 547963 69612 557506
rect 70308 552764 70360 552770
rect 70308 552706 70360 552712
rect 70320 547963 70348 552706
rect 70964 547963 70992 557506
rect 71056 555558 71084 571950
rect 74184 571402 74212 575076
rect 76024 575062 76774 575090
rect 74540 575000 74592 575006
rect 74540 574942 74592 574948
rect 71780 571396 71832 571402
rect 71780 571338 71832 571344
rect 74172 571396 74224 571402
rect 74172 571338 74224 571344
rect 71792 557534 71820 571338
rect 73252 561128 73304 561134
rect 73252 561070 73304 561076
rect 71792 557506 72464 557534
rect 71688 556844 71740 556850
rect 71688 556786 71740 556792
rect 71044 555552 71096 555558
rect 71044 555494 71096 555500
rect 71700 547963 71728 556786
rect 72436 547963 72464 557506
rect 73264 548162 73292 561070
rect 73804 550044 73856 550050
rect 73804 549986 73856 549992
rect 73188 548134 73292 548162
rect 73188 547944 73216 548134
rect 73816 547963 73844 549986
rect 74552 547963 74580 574942
rect 74632 572144 74684 572150
rect 74632 572086 74684 572092
rect 74644 557534 74672 572086
rect 75920 567996 75972 568002
rect 75920 567938 75972 567944
rect 74644 557506 75316 557534
rect 75288 547963 75316 557506
rect 75932 552786 75960 567938
rect 76024 556986 76052 575062
rect 78680 574932 78732 574938
rect 78680 574874 78732 574880
rect 76012 556980 76064 556986
rect 76012 556922 76064 556928
rect 77208 555484 77260 555490
rect 77208 555426 77260 555432
rect 76748 554124 76800 554130
rect 76748 554066 76800 554072
rect 75932 552758 76052 552786
rect 76024 547963 76052 552758
rect 76760 547963 76788 554066
rect 77220 550610 77248 555426
rect 78692 552770 78720 574874
rect 79324 572076 79376 572082
rect 79324 572018 79376 572024
rect 78772 563712 78824 563718
rect 78772 563654 78824 563660
rect 78784 557534 78812 563654
rect 78784 557506 78904 557534
rect 78680 552764 78732 552770
rect 78680 552706 78732 552712
rect 77220 550582 77432 550610
rect 77404 547963 77432 550582
rect 78128 550044 78180 550050
rect 78128 549986 78180 549992
rect 78140 547963 78168 549986
rect 78876 547963 78904 557506
rect 79336 550594 79364 572018
rect 79980 572014 80008 575076
rect 81452 575062 82570 575090
rect 79968 572008 80020 572014
rect 79968 571950 80020 571956
rect 80060 569356 80112 569362
rect 80060 569298 80112 569304
rect 80072 552786 80100 569298
rect 81452 563854 81480 575062
rect 82912 573504 82964 573510
rect 82912 573446 82964 573452
rect 84200 573504 84252 573510
rect 84200 573446 84252 573452
rect 81440 563848 81492 563854
rect 81440 563790 81492 563796
rect 80152 561060 80204 561066
rect 80152 561002 80204 561008
rect 80164 557534 80192 561002
rect 82924 557534 82952 573446
rect 84212 557534 84240 573446
rect 85776 572082 85804 575076
rect 88366 575062 88472 575090
rect 96804 575078 96856 575084
rect 86960 575000 87012 575006
rect 86960 574942 87012 574948
rect 86224 572212 86276 572218
rect 86224 572154 86276 572160
rect 85764 572076 85816 572082
rect 85764 572018 85816 572024
rect 85580 566568 85632 566574
rect 85580 566510 85632 566516
rect 85592 557534 85620 566510
rect 80164 557506 81020 557534
rect 82924 557506 83228 557534
rect 84212 557506 84608 557534
rect 85592 557506 86080 557534
rect 79600 552764 79652 552770
rect 80072 552758 80376 552786
rect 79600 552706 79652 552712
rect 79324 550588 79376 550594
rect 79324 550530 79376 550536
rect 79612 547963 79640 552706
rect 80348 547963 80376 552758
rect 80992 547963 81020 557506
rect 82452 555484 82504 555490
rect 82452 555426 82504 555432
rect 81716 550588 81768 550594
rect 81716 550530 81768 550536
rect 81728 547963 81756 550530
rect 82464 547963 82492 555426
rect 83200 547963 83228 557506
rect 83924 550248 83976 550254
rect 83924 550190 83976 550196
rect 83936 547963 83964 550190
rect 84580 547963 84608 557506
rect 85304 550248 85356 550254
rect 85304 550190 85356 550196
rect 85316 547963 85344 550190
rect 86052 547963 86080 557506
rect 86236 551342 86264 572154
rect 86776 556980 86828 556986
rect 86776 556922 86828 556928
rect 86224 551336 86276 551342
rect 86224 551278 86276 551284
rect 86788 547963 86816 556922
rect 86972 552786 87000 574942
rect 87052 574932 87104 574938
rect 87052 574874 87104 574880
rect 87064 557534 87092 574874
rect 88444 559638 88472 575062
rect 91572 570790 91600 575076
rect 93860 575068 93912 575074
rect 93860 575010 93912 575016
rect 92572 573572 92624 573578
rect 92572 573514 92624 573520
rect 91100 570784 91152 570790
rect 91100 570726 91152 570732
rect 91560 570784 91612 570790
rect 91560 570726 91612 570732
rect 89720 566636 89772 566642
rect 89720 566578 89772 566584
rect 88524 565208 88576 565214
rect 88524 565150 88576 565156
rect 88432 559632 88484 559638
rect 88432 559574 88484 559580
rect 88536 557534 88564 565150
rect 87064 557506 88196 557534
rect 88536 557506 89668 557534
rect 86972 552758 87460 552786
rect 87432 547963 87460 552758
rect 88168 547963 88196 557506
rect 88892 550384 88944 550390
rect 88892 550326 88944 550332
rect 88904 547963 88932 550326
rect 89640 547963 89668 557506
rect 89732 552770 89760 566578
rect 89812 563848 89864 563854
rect 89812 563790 89864 563796
rect 89824 557534 89852 563790
rect 91112 557534 91140 570726
rect 89824 557506 90404 557534
rect 91112 557506 91784 557534
rect 89720 552764 89772 552770
rect 89720 552706 89772 552712
rect 90376 547963 90404 557506
rect 91008 552764 91060 552770
rect 91008 552706 91060 552712
rect 91020 547963 91048 552706
rect 91756 547963 91784 557506
rect 92584 548162 92612 573514
rect 93872 557534 93900 575010
rect 94148 572218 94176 575076
rect 94136 572212 94188 572218
rect 94136 572154 94188 572160
rect 96712 570784 96764 570790
rect 96712 570726 96764 570732
rect 93872 557506 93992 557534
rect 93216 550316 93268 550322
rect 93216 550258 93268 550264
rect 92508 548134 92612 548162
rect 92508 547944 92536 548134
rect 93228 547963 93256 550258
rect 93964 547963 93992 557506
rect 96724 552786 96752 570726
rect 96816 557534 96844 575078
rect 97368 572150 97396 575076
rect 97356 572144 97408 572150
rect 97356 572086 97408 572092
rect 98104 557534 98132 575146
rect 99576 557534 99604 575214
rect 99944 572150 99972 575076
rect 102152 575062 103178 575090
rect 105004 575062 105754 575090
rect 99932 572144 99984 572150
rect 99932 572086 99984 572092
rect 100760 563780 100812 563786
rect 100760 563722 100812 563728
rect 100772 557534 100800 563722
rect 96816 557506 97488 557534
rect 98104 557506 98224 557534
rect 99576 557506 100432 557534
rect 100772 557506 101076 557534
rect 94596 552764 94648 552770
rect 96724 552758 96844 552786
rect 94596 552706 94648 552712
rect 94608 547963 94636 552706
rect 95332 550180 95384 550186
rect 95332 550122 95384 550128
rect 96068 550180 96120 550186
rect 96068 550122 96120 550128
rect 95344 547963 95372 550122
rect 96080 547963 96108 550122
rect 96816 547963 96844 552758
rect 97460 547963 97488 557506
rect 98196 547963 98224 557506
rect 98920 550112 98972 550118
rect 98920 550054 98972 550060
rect 98932 547963 98960 550054
rect 99656 549976 99708 549982
rect 99656 549918 99708 549924
rect 99668 547963 99696 549918
rect 100404 547963 100432 557506
rect 101048 547963 101076 557506
rect 102152 549386 102180 575062
rect 104900 572212 104952 572218
rect 104900 572154 104952 572160
rect 102232 562352 102284 562358
rect 102232 562294 102284 562300
rect 102244 557534 102272 562294
rect 103520 559632 103572 559638
rect 103520 559574 103572 559580
rect 103532 557534 103560 559574
rect 102244 557506 102548 557534
rect 103532 557506 104664 557534
rect 101876 549358 102180 549386
rect 101876 548162 101904 549358
rect 101800 548134 101904 548162
rect 101800 547944 101828 548134
rect 102520 547963 102548 557506
rect 103244 552696 103296 552702
rect 103244 552638 103296 552644
rect 103256 547963 103284 552638
rect 103980 549976 104032 549982
rect 103980 549918 104032 549924
rect 103992 547963 104020 549918
rect 104636 547963 104664 557506
rect 104912 552702 104940 572154
rect 105004 565214 105032 575062
rect 104992 565208 105044 565214
rect 104992 565150 105044 565156
rect 105360 555552 105412 555558
rect 105360 555494 105412 555500
rect 104900 552696 104952 552702
rect 104900 552638 104952 552644
rect 105372 547963 105400 555494
rect 106292 552702 106320 575282
rect 107672 575062 108974 575090
rect 110616 575062 111550 575090
rect 114572 575062 114770 575090
rect 107672 561134 107700 575062
rect 108304 572076 108356 572082
rect 108304 572018 108356 572024
rect 110420 572076 110472 572082
rect 110420 572018 110472 572024
rect 107660 561128 107712 561134
rect 107660 561070 107712 561076
rect 107660 559564 107712 559570
rect 107660 559506 107712 559512
rect 106096 552696 106148 552702
rect 106096 552638 106148 552644
rect 106280 552696 106332 552702
rect 106280 552638 106332 552644
rect 107568 552696 107620 552702
rect 107672 552684 107700 559506
rect 107752 558204 107804 558210
rect 107752 558146 107804 558152
rect 107764 552838 107792 558146
rect 107752 552832 107804 552838
rect 107752 552774 107804 552780
rect 107672 552656 108252 552684
rect 107568 552638 107620 552644
rect 106108 547963 106136 552638
rect 106832 550112 106884 550118
rect 106832 550054 106884 550060
rect 106844 547963 106872 550054
rect 107580 547963 107608 552638
rect 108224 547963 108252 552656
rect 108316 550594 108344 572018
rect 109684 556912 109736 556918
rect 109684 556854 109736 556860
rect 108948 552832 109000 552838
rect 108948 552774 109000 552780
rect 108304 550588 108356 550594
rect 108304 550530 108356 550536
rect 108960 547963 108988 552774
rect 109696 547963 109724 556854
rect 110432 547963 110460 572018
rect 110512 569288 110564 569294
rect 110512 569230 110564 569236
rect 110524 552684 110552 569230
rect 110616 554062 110644 575062
rect 111892 573640 111944 573646
rect 111892 573582 111944 573588
rect 111904 557534 111932 573582
rect 114572 567934 114600 575062
rect 115204 572144 115256 572150
rect 115204 572086 115256 572092
rect 114744 572008 114796 572014
rect 114744 571950 114796 571956
rect 114560 567928 114612 567934
rect 114560 567870 114612 567876
rect 111904 557506 112576 557534
rect 110604 554056 110656 554062
rect 110604 553998 110656 554004
rect 110524 552656 111104 552684
rect 111076 547963 111104 552656
rect 111800 550588 111852 550594
rect 111800 550530 111852 550536
rect 111812 547963 111840 550530
rect 112548 547963 112576 557506
rect 114756 552786 114784 571950
rect 115216 557534 115244 572086
rect 116676 571464 116728 571470
rect 116676 571406 116728 571412
rect 116584 571396 116636 571402
rect 116584 571338 116636 571344
rect 115216 557506 115520 557534
rect 114756 552758 115428 552786
rect 113272 552016 113324 552022
rect 113272 551958 113324 551964
rect 113284 547963 113312 551958
rect 114652 551336 114704 551342
rect 114652 551278 114704 551284
rect 114008 550316 114060 550322
rect 114008 550258 114060 550264
rect 114020 547963 114048 550258
rect 114664 547963 114692 551278
rect 115400 547963 115428 552758
rect 115492 550594 115520 557506
rect 116596 554130 116624 571338
rect 116688 555490 116716 571406
rect 117332 571402 117360 575076
rect 119344 574660 119396 574666
rect 119344 574602 119396 574608
rect 117320 571396 117372 571402
rect 117320 571338 117372 571344
rect 118700 569424 118752 569430
rect 118700 569366 118752 569372
rect 117320 560992 117372 560998
rect 117320 560934 117372 560940
rect 117332 557534 117360 560934
rect 118712 557534 118740 569366
rect 117332 557506 117636 557534
rect 118712 557506 119108 557534
rect 116676 555484 116728 555490
rect 116676 555426 116728 555432
rect 116584 554124 116636 554130
rect 116584 554066 116636 554072
rect 115480 550588 115532 550594
rect 115480 550530 115532 550536
rect 116124 550588 116176 550594
rect 116124 550530 116176 550536
rect 116136 547963 116164 550530
rect 116860 549908 116912 549914
rect 116860 549850 116912 549856
rect 116872 547963 116900 549850
rect 117608 547963 117636 557506
rect 118240 550452 118292 550458
rect 118240 550394 118292 550400
rect 118252 547963 118280 550394
rect 118976 550384 119028 550390
rect 118976 550326 119028 550332
rect 118988 547963 119016 550326
rect 119080 550066 119108 557506
rect 119356 550186 119384 574602
rect 120552 571470 120580 575076
rect 120540 571464 120592 571470
rect 120540 571406 120592 571412
rect 120736 570722 120764 576807
rect 120724 570716 120776 570722
rect 120724 570658 120776 570664
rect 120828 569362 120856 613255
rect 120816 569356 120868 569362
rect 120816 569298 120868 569304
rect 120448 551336 120500 551342
rect 120448 551278 120500 551284
rect 119344 550180 119396 550186
rect 119344 550122 119396 550128
rect 119080 550038 119752 550066
rect 119724 547963 119752 550038
rect 120460 547963 120488 551278
rect 120920 550254 120948 640426
rect 121000 640416 121052 640422
rect 121000 640358 121052 640364
rect 121012 575210 121040 640358
rect 121090 598224 121146 598233
rect 121090 598159 121146 598168
rect 121000 575204 121052 575210
rect 121000 575146 121052 575152
rect 121104 561066 121132 598159
rect 121184 581664 121236 581670
rect 121184 581606 121236 581612
rect 121196 572082 121224 581606
rect 121472 575006 121500 640562
rect 121552 640552 121604 640558
rect 121552 640494 121604 640500
rect 121460 575000 121512 575006
rect 121460 574942 121512 574948
rect 121184 572076 121236 572082
rect 121184 572018 121236 572024
rect 121460 570784 121512 570790
rect 121460 570726 121512 570732
rect 121092 561060 121144 561066
rect 121092 561002 121144 561008
rect 121092 555620 121144 555626
rect 121092 555562 121144 555568
rect 120908 550248 120960 550254
rect 120908 550190 120960 550196
rect 121104 547963 121132 555562
rect 121472 552702 121500 570726
rect 121460 552696 121512 552702
rect 121460 552638 121512 552644
rect 121564 550050 121592 640494
rect 121734 628824 121790 628833
rect 121734 628759 121790 628768
rect 121642 622704 121698 622713
rect 121642 622639 121698 622648
rect 121656 556850 121684 622639
rect 121748 566574 121776 628759
rect 121826 616584 121882 616593
rect 121826 616519 121882 616528
rect 121840 567866 121868 616519
rect 122010 601624 122066 601633
rect 122010 601559 122066 601568
rect 121918 579864 121974 579873
rect 121918 579799 121974 579808
rect 121828 567860 121880 567866
rect 121828 567802 121880 567808
rect 121736 566568 121788 566574
rect 121736 566510 121788 566516
rect 121644 556844 121696 556850
rect 121644 556786 121696 556792
rect 121932 552022 121960 579799
rect 122024 573442 122052 601559
rect 122102 595504 122158 595513
rect 122102 595439 122158 595448
rect 122116 573510 122144 595439
rect 122194 592104 122250 592113
rect 122194 592039 122250 592048
rect 122208 574870 122236 592039
rect 122286 589384 122342 589393
rect 122286 589319 122342 589328
rect 122300 575278 122328 589319
rect 122288 575272 122340 575278
rect 122288 575214 122340 575220
rect 122852 575142 122880 640630
rect 124220 637764 124272 637770
rect 124220 637706 124272 637712
rect 122930 634944 122986 634953
rect 122930 634879 122986 634888
rect 122840 575136 122892 575142
rect 122840 575078 122892 575084
rect 122196 574864 122248 574870
rect 122196 574806 122248 574812
rect 122840 573572 122892 573578
rect 122840 573514 122892 573520
rect 122104 573504 122156 573510
rect 122104 573446 122156 573452
rect 122012 573436 122064 573442
rect 122012 573378 122064 573384
rect 122852 552702 122880 573514
rect 122944 566506 122972 634879
rect 123022 632224 123078 632233
rect 123022 632159 123078 632168
rect 123036 573646 123064 632159
rect 123114 626104 123170 626113
rect 123114 626039 123170 626048
rect 123024 573640 123076 573646
rect 123024 573582 123076 573588
rect 123128 569226 123156 626039
rect 123206 619984 123262 619993
rect 123206 619919 123262 619928
rect 123116 569220 123168 569226
rect 123116 569162 123168 569168
rect 123024 566636 123076 566642
rect 123024 566578 123076 566584
rect 122932 566500 122984 566506
rect 122932 566442 122984 566448
rect 122564 552696 122616 552702
rect 122564 552638 122616 552644
rect 122840 552696 122892 552702
rect 123036 552684 123064 566578
rect 123220 565146 123248 619919
rect 123390 610464 123446 610473
rect 123390 610399 123446 610408
rect 123300 601044 123352 601050
rect 123300 600986 123352 600992
rect 123208 565140 123260 565146
rect 123208 565082 123260 565088
rect 123312 552838 123340 600986
rect 123404 574666 123432 610399
rect 123482 607744 123538 607753
rect 123482 607679 123538 607688
rect 123496 601050 123524 607679
rect 124126 604344 124182 604353
rect 124126 604279 124182 604288
rect 124140 603158 124168 604279
rect 124128 603152 124180 603158
rect 124128 603094 124180 603100
rect 123484 601044 123536 601050
rect 123484 600986 123536 600992
rect 123482 585984 123538 585993
rect 123482 585919 123538 585928
rect 123392 574660 123444 574666
rect 123392 574602 123444 574608
rect 123496 563718 123524 585919
rect 123574 583264 123630 583273
rect 123574 583199 123630 583208
rect 123588 574802 123616 583199
rect 123576 574796 123628 574802
rect 123576 574738 123628 574744
rect 123484 563712 123536 563718
rect 123484 563654 123536 563660
rect 123300 552832 123352 552838
rect 123300 552774 123352 552780
rect 124232 552770 124260 637706
rect 124312 637696 124364 637702
rect 124312 637638 124364 637644
rect 124220 552764 124272 552770
rect 124220 552706 124272 552712
rect 124036 552696 124088 552702
rect 123036 552656 123340 552684
rect 122840 552638 122892 552644
rect 121920 552016 121972 552022
rect 121920 551958 121972 551964
rect 121552 550044 121604 550050
rect 121552 549986 121604 549992
rect 121828 549908 121880 549914
rect 121828 549850 121880 549856
rect 121840 547963 121868 549850
rect 122576 547963 122604 552638
rect 123312 547963 123340 552656
rect 124036 552638 124088 552644
rect 124048 547963 124076 552638
rect 124324 550118 124352 637638
rect 124416 550322 124444 640766
rect 124496 640756 124548 640762
rect 124496 640698 124548 640704
rect 124508 575074 124536 640698
rect 124588 640348 124640 640354
rect 124588 640290 124640 640296
rect 124496 575068 124548 575074
rect 124496 575010 124548 575016
rect 124600 574938 124628 640290
rect 124692 575346 124720 640834
rect 126244 638036 126296 638042
rect 126244 637978 126296 637984
rect 125784 637832 125836 637838
rect 125784 637774 125836 637780
rect 125600 592068 125652 592074
rect 125600 592010 125652 592016
rect 124680 575340 124732 575346
rect 124680 575282 124732 575288
rect 124588 574932 124640 574938
rect 124588 574874 124640 574880
rect 124680 556912 124732 556918
rect 124680 556854 124732 556860
rect 124404 550316 124456 550322
rect 124404 550258 124456 550264
rect 124312 550112 124364 550118
rect 124312 550054 124364 550060
rect 124692 547963 124720 556854
rect 125612 556102 125640 592010
rect 125692 567928 125744 567934
rect 125692 567870 125744 567876
rect 125600 556096 125652 556102
rect 125600 556038 125652 556044
rect 125416 552764 125468 552770
rect 125416 552706 125468 552712
rect 125428 547963 125456 552706
rect 125704 549794 125732 567870
rect 125796 549982 125824 637774
rect 126256 550458 126284 637978
rect 129004 604512 129056 604518
rect 129004 604454 129056 604460
rect 126980 574932 127032 574938
rect 126980 574874 127032 574880
rect 126888 556096 126940 556102
rect 126888 556038 126940 556044
rect 126244 550452 126296 550458
rect 126244 550394 126296 550400
rect 125784 549976 125836 549982
rect 125784 549918 125836 549924
rect 125704 549766 126192 549794
rect 126164 547963 126192 549766
rect 126900 547963 126928 556038
rect 126992 552770 127020 574874
rect 128360 567996 128412 568002
rect 128360 567938 128412 567944
rect 127072 559632 127124 559638
rect 127072 559574 127124 559580
rect 127084 557534 127112 559574
rect 127084 557506 127664 557534
rect 126980 552764 127032 552770
rect 126980 552706 127032 552712
rect 127636 547963 127664 557506
rect 128268 552764 128320 552770
rect 128268 552706 128320 552712
rect 128280 547963 128308 552706
rect 128372 552684 128400 567938
rect 129016 557534 129044 604454
rect 130384 589348 130436 589354
rect 130384 589290 130436 589296
rect 129740 572144 129792 572150
rect 129740 572086 129792 572092
rect 129016 557506 129136 557534
rect 128372 552656 129044 552684
rect 129016 547963 129044 552656
rect 129108 550390 129136 557506
rect 129752 552770 129780 572086
rect 129832 565276 129884 565282
rect 129832 565218 129884 565224
rect 129740 552764 129792 552770
rect 129740 552706 129792 552712
rect 129096 550384 129148 550390
rect 129096 550326 129148 550332
rect 129844 548162 129872 565218
rect 130396 551342 130424 589290
rect 131132 557534 131160 640970
rect 145012 640960 145064 640966
rect 145012 640902 145064 640908
rect 140780 640824 140832 640830
rect 140780 640766 140832 640772
rect 133880 640348 133932 640354
rect 133880 640290 133932 640296
rect 132500 622464 132552 622470
rect 132500 622406 132552 622412
rect 131132 557506 131896 557534
rect 130476 552764 130528 552770
rect 130476 552706 130528 552712
rect 130384 551336 130436 551342
rect 130384 551278 130436 551284
rect 129768 548134 129872 548162
rect 129768 547944 129796 548134
rect 130488 547963 130516 552706
rect 131212 549296 131264 549302
rect 131212 549238 131264 549244
rect 131224 547963 131252 549238
rect 131868 547963 131896 557506
rect 132512 554146 132540 622406
rect 132592 572076 132644 572082
rect 132592 572018 132644 572024
rect 132604 557534 132632 572018
rect 133144 558204 133196 558210
rect 133144 558146 133196 558152
rect 132604 557506 133092 557534
rect 132512 554118 132632 554146
rect 132604 547963 132632 554118
rect 133064 549114 133092 557506
rect 133156 549302 133184 558146
rect 133892 552786 133920 640290
rect 136640 637900 136692 637906
rect 136640 637842 136692 637848
rect 133972 572008 134024 572014
rect 133972 571950 134024 571956
rect 133984 557534 134012 571950
rect 133984 557506 134748 557534
rect 133892 552758 134104 552786
rect 133144 549296 133196 549302
rect 133144 549238 133196 549244
rect 133064 549086 133368 549114
rect 133340 547963 133368 549086
rect 134076 547963 134104 552758
rect 134720 547963 134748 557506
rect 136652 552770 136680 637842
rect 140044 637832 140096 637838
rect 140044 637774 140096 637780
rect 139400 586560 139452 586566
rect 139400 586502 139452 586508
rect 136732 563916 136784 563922
rect 136732 563858 136784 563864
rect 136744 557534 136772 563858
rect 138020 561060 138072 561066
rect 138020 561002 138072 561008
rect 138032 557534 138060 561002
rect 139412 557534 139440 586502
rect 136744 557506 136956 557534
rect 138032 557506 139072 557534
rect 139412 557506 139808 557534
rect 136640 552764 136692 552770
rect 136640 552706 136692 552712
rect 135444 550792 135496 550798
rect 135444 550734 135496 550740
rect 135456 547963 135484 550734
rect 136180 550588 136232 550594
rect 136180 550530 136232 550536
rect 136192 547963 136220 550530
rect 136928 547963 136956 557506
rect 137652 552764 137704 552770
rect 137652 552706 137704 552712
rect 137664 547963 137692 552706
rect 138296 549432 138348 549438
rect 138296 549374 138348 549380
rect 138308 547963 138336 549374
rect 139044 547963 139072 557506
rect 139780 547963 139808 557506
rect 140056 550594 140084 637774
rect 140504 554056 140556 554062
rect 140504 553998 140556 554004
rect 140044 550588 140096 550594
rect 140044 550530 140096 550536
rect 140516 547963 140544 553998
rect 140792 552770 140820 640766
rect 142160 640620 142212 640626
rect 142160 640562 142212 640568
rect 140872 626612 140924 626618
rect 140872 626554 140924 626560
rect 140884 557534 140912 626554
rect 140884 557506 141280 557534
rect 140780 552764 140832 552770
rect 140780 552706 140832 552712
rect 141252 547963 141280 557506
rect 142172 552770 142200 640562
rect 144920 640552 144972 640558
rect 144920 640494 144972 640500
rect 144184 635248 144236 635254
rect 144184 635190 144236 635196
rect 143540 572348 143592 572354
rect 143540 572290 143592 572296
rect 142804 569288 142856 569294
rect 142804 569230 142856 569236
rect 141884 552764 141936 552770
rect 141884 552706 141936 552712
rect 142160 552764 142212 552770
rect 142160 552706 142212 552712
rect 141896 547963 141924 552706
rect 142620 551336 142672 551342
rect 142620 551278 142672 551284
rect 142632 547963 142660 551278
rect 142816 549438 142844 569230
rect 143552 552770 143580 572290
rect 143356 552764 143408 552770
rect 143356 552706 143408 552712
rect 143540 552764 143592 552770
rect 143540 552706 143592 552712
rect 142804 549432 142856 549438
rect 142804 549374 142856 549380
rect 143368 547963 143396 552706
rect 144196 550798 144224 635190
rect 144736 552764 144788 552770
rect 144932 552752 144960 640494
rect 145024 552906 145052 640902
rect 146116 637696 146168 637702
rect 146116 637638 146168 637644
rect 145564 603152 145616 603158
rect 145564 603094 145616 603100
rect 145576 575414 145604 603094
rect 145564 575408 145616 575414
rect 145564 575350 145616 575356
rect 145012 552900 145064 552906
rect 145012 552842 145064 552848
rect 144932 552724 145512 552752
rect 144736 552706 144788 552712
rect 144184 550792 144236 550798
rect 144184 550734 144236 550740
rect 144092 550588 144144 550594
rect 144092 550530 144144 550536
rect 144104 547963 144132 550530
rect 144748 547963 144776 552706
rect 145484 547963 145512 552724
rect 146128 550118 146156 637638
rect 146208 637628 146260 637634
rect 146208 637570 146260 637576
rect 146220 611153 146248 637570
rect 147126 635624 147182 635633
rect 147126 635559 147182 635568
rect 147140 635254 147168 635559
rect 147128 635248 147180 635254
rect 147128 635190 147180 635196
rect 146298 626784 146354 626793
rect 146298 626719 146354 626728
rect 146312 626618 146340 626719
rect 146300 626612 146352 626618
rect 146300 626554 146352 626560
rect 146298 623384 146354 623393
rect 146298 623319 146354 623328
rect 146312 622470 146340 623319
rect 146300 622464 146352 622470
rect 146300 622406 146352 622412
rect 147232 614553 147260 683130
rect 299492 646542 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 305644 700460 305696 700466
rect 305644 700402 305696 700408
rect 299480 646536 299532 646542
rect 299480 646478 299532 646484
rect 233240 641164 233292 641170
rect 233240 641106 233292 641112
rect 147588 641096 147640 641102
rect 147588 641038 147640 641044
rect 164516 641096 164568 641102
rect 164516 641038 164568 641044
rect 147312 640484 147364 640490
rect 147312 640426 147364 640432
rect 147218 614544 147274 614553
rect 147218 614479 147274 614488
rect 146206 611144 146262 611153
rect 146206 611079 146262 611088
rect 146298 605024 146354 605033
rect 146298 604959 146354 604968
rect 146312 604518 146340 604959
rect 146300 604512 146352 604518
rect 146300 604454 146352 604460
rect 147126 602304 147182 602313
rect 147126 602239 147182 602248
rect 146298 592784 146354 592793
rect 146298 592719 146354 592728
rect 146312 592074 146340 592719
rect 146300 592068 146352 592074
rect 146300 592010 146352 592016
rect 146298 590064 146354 590073
rect 146298 589999 146354 590008
rect 146312 589354 146340 589999
rect 146300 589348 146352 589354
rect 146300 589290 146352 589296
rect 146298 586664 146354 586673
rect 146298 586599 146354 586608
rect 146312 586566 146340 586599
rect 146300 586560 146352 586566
rect 146300 586502 146352 586508
rect 147034 583944 147090 583953
rect 147034 583879 147090 583888
rect 147048 566506 147076 583879
rect 147140 572762 147168 602239
rect 147218 596184 147274 596193
rect 147218 596119 147274 596128
rect 147128 572756 147180 572762
rect 147128 572698 147180 572704
rect 147036 566500 147088 566506
rect 147036 566442 147088 566448
rect 146944 562420 146996 562426
rect 146944 562362 146996 562368
rect 146956 557534 146984 562362
rect 147232 560998 147260 596119
rect 147324 575074 147352 640426
rect 147494 629504 147550 629513
rect 147494 629439 147550 629448
rect 147402 620664 147458 620673
rect 147402 620599 147458 620608
rect 147312 575068 147364 575074
rect 147312 575010 147364 575016
rect 147416 569226 147444 620599
rect 147404 569220 147456 569226
rect 147404 569162 147456 569168
rect 147220 560992 147272 560998
rect 147220 560934 147272 560940
rect 146864 557506 146984 557534
rect 146208 552900 146260 552906
rect 146208 552842 146260 552848
rect 146116 550112 146168 550118
rect 146116 550054 146168 550060
rect 146220 547963 146248 552842
rect 146864 550594 146892 557506
rect 147508 551410 147536 629439
rect 147496 551404 147548 551410
rect 147496 551346 147548 551352
rect 146852 550588 146904 550594
rect 146852 550530 146904 550536
rect 146944 550588 146996 550594
rect 146944 550530 146996 550536
rect 146956 547963 146984 550530
rect 147600 550186 147628 641038
rect 161572 641028 161624 641034
rect 161572 640970 161624 640976
rect 148876 640892 148928 640898
rect 148876 640834 148928 640840
rect 148784 640756 148836 640762
rect 148784 640698 148836 640704
rect 148324 638988 148376 638994
rect 148324 638930 148376 638936
rect 147680 552764 147732 552770
rect 147680 552706 147732 552712
rect 147588 550180 147640 550186
rect 147588 550122 147640 550128
rect 147692 547963 147720 552706
rect 148336 550594 148364 638930
rect 148598 632904 148654 632913
rect 148598 632839 148654 632848
rect 148414 608424 148470 608433
rect 148414 608359 148470 608368
rect 148428 576842 148456 608359
rect 148506 598904 148562 598913
rect 148506 598839 148562 598848
rect 148416 576836 148468 576842
rect 148416 576778 148468 576784
rect 148416 554124 148468 554130
rect 148416 554066 148468 554072
rect 148324 550588 148376 550594
rect 148324 550530 148376 550536
rect 148428 548162 148456 554066
rect 148520 552022 148548 598839
rect 148612 575210 148640 632839
rect 148690 617264 148746 617273
rect 148690 617199 148746 617208
rect 148600 575204 148652 575210
rect 148600 575146 148652 575152
rect 148704 555490 148732 617199
rect 148796 574870 148824 640698
rect 148784 574864 148836 574870
rect 148784 574806 148836 574812
rect 148888 574802 148916 640834
rect 149520 640688 149572 640694
rect 149520 640630 149572 640636
rect 148968 637968 149020 637974
rect 148968 637910 149020 637916
rect 148876 574796 148928 574802
rect 148876 574738 148928 574744
rect 148692 555484 148744 555490
rect 148692 555426 148744 555432
rect 148508 552016 148560 552022
rect 148508 551958 148560 551964
rect 148980 549982 149008 637910
rect 149532 634814 149560 640630
rect 149612 640416 149664 640422
rect 149612 640358 149664 640364
rect 149624 637650 149652 640358
rect 149980 640348 150032 640354
rect 149980 640290 150032 640296
rect 149888 639056 149940 639062
rect 149888 638998 149940 639004
rect 149624 637622 149836 637650
rect 149532 634786 149744 634814
rect 149716 580802 149744 634786
rect 149348 580774 149744 580802
rect 149348 575346 149376 580774
rect 149808 580666 149836 637622
rect 149716 580638 149836 580666
rect 149610 577788 149666 577797
rect 149610 577723 149666 577732
rect 149428 576836 149480 576842
rect 149428 576778 149480 576784
rect 149336 575340 149388 575346
rect 149336 575282 149388 575288
rect 149440 557534 149468 576778
rect 149624 573442 149652 577723
rect 149716 575278 149744 580638
rect 149794 580508 149850 580517
rect 149794 580443 149850 580452
rect 149704 575272 149756 575278
rect 149704 575214 149756 575220
rect 149808 575006 149836 580443
rect 149796 575000 149848 575006
rect 149796 574942 149848 574948
rect 149612 573436 149664 573442
rect 149612 573378 149664 573384
rect 149440 557506 149836 557534
rect 149060 552016 149112 552022
rect 149060 551958 149112 551964
rect 148968 549976 149020 549982
rect 148968 549918 149020 549924
rect 148352 548134 148456 548162
rect 148352 547944 148380 548134
rect 149072 547963 149100 551958
rect 149808 547963 149836 557506
rect 149900 550594 149928 638998
rect 149992 638058 150020 640290
rect 153200 638988 153252 638994
rect 153200 638930 153252 638936
rect 153212 638058 153240 638930
rect 161584 638058 161612 640970
rect 164528 638058 164556 641038
rect 207664 640960 207716 640966
rect 207664 640902 207716 640908
rect 172888 640892 172940 640898
rect 172888 640834 172940 640840
rect 167092 640824 167144 640830
rect 167092 640766 167144 640772
rect 167104 638058 167132 640766
rect 170312 639056 170364 639062
rect 170312 638998 170364 639004
rect 170324 638058 170352 638998
rect 172900 638058 172928 640834
rect 176108 640756 176160 640762
rect 176108 640698 176160 640704
rect 176120 638058 176148 640698
rect 190552 640688 190604 640694
rect 190552 640630 190604 640636
rect 184480 640620 184532 640626
rect 184480 640562 184532 640568
rect 184492 638058 184520 640562
rect 190564 638058 190592 640630
rect 196072 640552 196124 640558
rect 196072 640494 196124 640500
rect 196084 638058 196112 640494
rect 199292 640484 199344 640490
rect 199292 640426 199344 640432
rect 199304 638058 199332 640426
rect 201868 640416 201920 640422
rect 201868 640358 201920 640364
rect 205548 640416 205600 640422
rect 205548 640358 205600 640364
rect 201880 638058 201908 640358
rect 205560 638058 205588 640358
rect 149992 638030 150052 638058
rect 153212 638030 153272 638058
rect 161584 638030 161644 638058
rect 164528 638030 164864 638058
rect 167104 638030 167440 638058
rect 170324 638030 170660 638058
rect 172900 638030 173236 638058
rect 176120 638030 176456 638058
rect 184492 638030 184828 638058
rect 187712 638042 188048 638058
rect 187700 638036 188048 638042
rect 187752 638030 188048 638036
rect 190564 638030 190624 638058
rect 196084 638030 196420 638058
rect 199304 638030 199640 638058
rect 201880 638030 202216 638058
rect 205436 638030 205588 638058
rect 207676 638058 207704 640902
rect 226340 640824 226392 640830
rect 226340 640766 226392 640772
rect 217416 640620 217468 640626
rect 217416 640562 217468 640568
rect 212632 640416 212684 640422
rect 212632 640358 212684 640364
rect 207676 638030 208012 638058
rect 187700 637978 187752 637984
rect 158720 637968 158772 637974
rect 158772 637916 159068 637922
rect 158720 637910 159068 637916
rect 158732 637894 159068 637910
rect 178696 637906 179032 637922
rect 178684 637900 179032 637906
rect 178736 637894 179032 637900
rect 178684 637842 178736 637848
rect 193496 637832 193548 637838
rect 182100 637770 182252 637786
rect 193548 637780 193844 637786
rect 193496 637774 193844 637780
rect 182088 637764 182252 637770
rect 182140 637758 182252 637764
rect 193508 637758 193844 637774
rect 182088 637706 182140 637712
rect 155500 637696 155552 637702
rect 155552 637644 155848 637650
rect 155500 637638 155848 637644
rect 155512 637622 155848 637638
rect 210588 637350 210740 637378
rect 151820 575340 151872 575346
rect 151820 575282 151872 575288
rect 150532 575204 150584 575210
rect 150532 575146 150584 575152
rect 150052 575062 150388 575090
rect 150360 571402 150388 575062
rect 150348 571396 150400 571402
rect 150348 571338 150400 571344
rect 149888 550588 149940 550594
rect 149888 550530 149940 550536
rect 150544 547963 150572 575146
rect 151084 572756 151136 572762
rect 151084 572698 151136 572704
rect 151096 550322 151124 572698
rect 151176 571396 151228 571402
rect 151176 571338 151228 571344
rect 151188 552702 151216 571338
rect 151832 552786 151860 575282
rect 154764 575272 154816 575278
rect 154764 575214 154816 575220
rect 151924 575062 152628 575090
rect 151924 553738 151952 575062
rect 154672 572280 154724 572286
rect 154672 572222 154724 572228
rect 152004 563848 152056 563854
rect 152004 563790 152056 563796
rect 152016 557534 152044 563790
rect 152016 557506 152688 557534
rect 151924 553710 152044 553738
rect 151832 552758 151952 552786
rect 151176 552696 151228 552702
rect 151176 552638 151228 552644
rect 151268 550588 151320 550594
rect 151268 550530 151320 550536
rect 151084 550316 151136 550322
rect 151084 550258 151136 550264
rect 151280 547963 151308 550530
rect 151924 547963 151952 552758
rect 152016 550050 152044 553710
rect 152004 550044 152056 550050
rect 152004 549986 152056 549992
rect 152660 547963 152688 557506
rect 154120 555688 154172 555694
rect 154120 555630 154172 555636
rect 153384 550316 153436 550322
rect 153384 550258 153436 550264
rect 153396 547963 153424 550258
rect 154132 547963 154160 555630
rect 154684 552786 154712 572222
rect 154776 557534 154804 575214
rect 154868 575062 155204 575090
rect 156052 575068 156104 575074
rect 154868 569430 154896 575062
rect 156052 575010 156104 575016
rect 157352 575062 158424 575090
rect 160204 575062 161000 575090
rect 163884 575062 164220 575090
rect 166460 575062 166796 575090
rect 169772 575062 170016 575090
rect 172532 575062 172592 575090
rect 175476 575062 175812 575090
rect 178052 575062 178388 575090
rect 181272 575062 181608 575090
rect 183848 575062 184184 575090
rect 187068 575062 187404 575090
rect 189644 575062 189980 575090
rect 192864 575062 193200 575090
rect 195244 575068 195296 575074
rect 154856 569424 154908 569430
rect 154856 569366 154908 569372
rect 156064 557534 156092 575010
rect 154776 557506 155540 557534
rect 156064 557506 156276 557534
rect 154684 552758 154896 552786
rect 154868 547963 154896 552758
rect 155512 547963 155540 557506
rect 156248 547963 156276 557506
rect 157352 550322 157380 575062
rect 158720 573436 158772 573442
rect 158720 573378 158772 573384
rect 157432 569356 157484 569362
rect 157432 569298 157484 569304
rect 157444 557534 157472 569298
rect 157444 557506 158392 557534
rect 157340 550316 157392 550322
rect 157340 550258 157392 550264
rect 157708 550180 157760 550186
rect 157708 550122 157760 550128
rect 156972 550112 157024 550118
rect 156972 550054 157024 550060
rect 156984 547963 157012 550054
rect 157720 547963 157748 550122
rect 158364 547963 158392 557506
rect 158732 553394 158760 573378
rect 158812 572212 158864 572218
rect 158812 572154 158864 572160
rect 158824 557534 158852 572154
rect 158824 557506 159864 557534
rect 158732 553366 159128 553394
rect 159100 547963 159128 553366
rect 159836 547963 159864 557506
rect 160204 550186 160232 575062
rect 160284 575000 160336 575006
rect 160284 574942 160336 574948
rect 160296 557534 160324 574942
rect 161480 574864 161532 574870
rect 161480 574806 161532 574812
rect 160296 557506 161336 557534
rect 160560 555484 160612 555490
rect 160560 555426 160612 555432
rect 160192 550180 160244 550186
rect 160192 550122 160244 550128
rect 160572 547963 160600 555426
rect 161308 547963 161336 557506
rect 161492 553394 161520 574806
rect 161572 572484 161624 572490
rect 161572 572426 161624 572432
rect 161584 557534 161612 572426
rect 163044 572416 163096 572422
rect 163044 572358 163096 572364
rect 163056 557534 163084 572358
rect 163884 572150 163912 575062
rect 164332 575000 164384 575006
rect 164332 574942 164384 574948
rect 164240 574796 164292 574802
rect 164240 574738 164292 574744
rect 163872 572144 163924 572150
rect 163872 572086 163924 572092
rect 161584 557506 162716 557534
rect 163056 557506 164188 557534
rect 161492 553366 161980 553394
rect 161952 547963 161980 553366
rect 162688 547963 162716 557506
rect 163412 552696 163464 552702
rect 163412 552638 163464 552644
rect 163424 547963 163452 552638
rect 164160 547963 164188 557506
rect 164252 550610 164280 574738
rect 164344 550730 164372 574942
rect 166460 572354 166488 575062
rect 166448 572348 166500 572354
rect 166448 572290 166500 572296
rect 165620 569220 165672 569226
rect 165620 569162 165672 569168
rect 165632 557534 165660 569162
rect 168380 566500 168432 566506
rect 168380 566442 168432 566448
rect 165632 557506 166304 557534
rect 164332 550724 164384 550730
rect 164332 550666 164384 550672
rect 165528 550724 165580 550730
rect 165528 550666 165580 550672
rect 164252 550582 164924 550610
rect 164896 547963 164924 550582
rect 165540 547963 165568 550666
rect 166276 547963 166304 557506
rect 168392 552702 168420 566442
rect 168472 565208 168524 565214
rect 168472 565150 168524 565156
rect 168380 552696 168432 552702
rect 168380 552638 168432 552644
rect 167000 551404 167052 551410
rect 167000 551346 167052 551352
rect 167012 550050 167040 551346
rect 167092 550316 167144 550322
rect 167092 550258 167144 550264
rect 167000 550044 167052 550050
rect 167000 549986 167052 549992
rect 167104 548162 167132 550258
rect 167736 549976 167788 549982
rect 167736 549918 167788 549924
rect 167028 548134 167132 548162
rect 167028 547944 167056 548134
rect 167748 547963 167776 549918
rect 168484 548162 168512 565150
rect 169116 552696 169168 552702
rect 169116 552638 169168 552644
rect 168408 548134 168512 548162
rect 168408 547944 168436 548134
rect 169128 547963 169156 552638
rect 169772 549778 169800 575062
rect 169852 572348 169904 572354
rect 169852 572290 169904 572296
rect 169760 549772 169812 549778
rect 169760 549714 169812 549720
rect 169864 547963 169892 572290
rect 172532 554130 172560 575062
rect 175476 572354 175504 575062
rect 178052 572490 178080 575062
rect 179420 574796 179472 574802
rect 179420 574738 179472 574744
rect 178040 572484 178092 572490
rect 178040 572426 178092 572432
rect 175464 572348 175516 572354
rect 175464 572290 175516 572296
rect 173900 572144 173952 572150
rect 173900 572086 173952 572092
rect 172520 554124 172572 554130
rect 172520 554066 172572 554072
rect 171324 552832 171376 552838
rect 171324 552774 171376 552780
rect 170588 550112 170640 550118
rect 170588 550054 170640 550060
rect 170600 547963 170628 550054
rect 171336 547963 171364 552774
rect 173912 552684 173940 572086
rect 176660 568064 176712 568070
rect 176660 568006 176712 568012
rect 173992 560992 174044 560998
rect 173992 560934 174044 560940
rect 174004 557534 174032 560934
rect 174004 557506 174952 557534
rect 173912 552656 174216 552684
rect 172704 550180 172756 550186
rect 172704 550122 172756 550128
rect 171968 549908 172020 549914
rect 171968 549850 172020 549856
rect 171980 547963 172008 549850
rect 172716 547963 172744 550122
rect 173440 549772 173492 549778
rect 173440 549714 173492 549720
rect 173452 547963 173480 549714
rect 174188 547963 174216 552656
rect 174924 547963 174952 557506
rect 176672 552684 176700 568006
rect 176752 565344 176804 565350
rect 176752 565286 176804 565292
rect 176764 557534 176792 565286
rect 178040 561196 178092 561202
rect 178040 561138 178092 561144
rect 178052 557534 178080 561138
rect 176764 557506 177804 557534
rect 178052 557506 178540 557534
rect 176672 552656 177068 552684
rect 175556 550044 175608 550050
rect 175556 549986 175608 549992
rect 175568 547963 175596 549986
rect 176292 549976 176344 549982
rect 176292 549918 176344 549924
rect 176304 547963 176332 549918
rect 177040 547963 177068 552656
rect 177776 547963 177804 557506
rect 178512 547963 178540 557506
rect 179144 556844 179196 556850
rect 179144 556786 179196 556792
rect 179156 547963 179184 556786
rect 179432 552702 179460 574738
rect 179512 573436 179564 573442
rect 179512 573378 179564 573384
rect 179524 557534 179552 573378
rect 181272 572286 181300 575062
rect 183652 574864 183704 574870
rect 183652 574806 183704 574812
rect 181260 572280 181312 572286
rect 181260 572222 181312 572228
rect 180800 570716 180852 570722
rect 180800 570658 180852 570664
rect 179524 557506 179920 557534
rect 179420 552696 179472 552702
rect 179420 552638 179472 552644
rect 179892 547963 179920 557506
rect 180812 552702 180840 570658
rect 182180 559564 182232 559570
rect 182180 559506 182232 559512
rect 182192 557534 182220 559506
rect 183664 557534 183692 574806
rect 183848 572422 183876 575062
rect 183836 572416 183888 572422
rect 183836 572358 183888 572364
rect 187068 572082 187096 575062
rect 189644 572150 189672 575062
rect 192864 572218 192892 575062
rect 195244 575010 195296 575016
rect 195440 575062 195776 575090
rect 198844 575062 198996 575090
rect 201512 575062 201572 575090
rect 204272 575062 204792 575090
rect 207032 575062 207368 575090
rect 210252 575062 210588 575090
rect 192852 572212 192904 572218
rect 192852 572154 192904 572160
rect 189632 572144 189684 572150
rect 189632 572086 189684 572092
rect 193864 572144 193916 572150
rect 193864 572086 193916 572092
rect 187056 572076 187108 572082
rect 187056 572018 187108 572024
rect 192484 572076 192536 572082
rect 192484 572018 192536 572024
rect 191104 571396 191156 571402
rect 191104 571338 191156 571344
rect 186320 569220 186372 569226
rect 186320 569162 186372 569168
rect 184940 566568 184992 566574
rect 184940 566510 184992 566516
rect 184952 557534 184980 566510
rect 182192 557506 182772 557534
rect 183664 557506 184244 557534
rect 184952 557506 185624 557534
rect 180616 552696 180668 552702
rect 180616 552638 180668 552644
rect 180800 552696 180852 552702
rect 180800 552638 180852 552644
rect 181996 552696 182048 552702
rect 181996 552638 182048 552644
rect 180628 547963 180656 552638
rect 181352 552628 181404 552634
rect 181352 552570 181404 552576
rect 181364 547963 181392 552570
rect 182008 547963 182036 552638
rect 182744 547963 182772 557506
rect 183468 550044 183520 550050
rect 183468 549986 183520 549992
rect 183480 547963 183508 549986
rect 184216 547963 184244 557506
rect 184940 554192 184992 554198
rect 184940 554134 184992 554140
rect 184952 547963 184980 554134
rect 185596 547963 185624 557506
rect 186332 547963 186360 569162
rect 187700 566500 187752 566506
rect 187700 566442 187752 566448
rect 186412 563712 186464 563718
rect 186412 563654 186464 563660
rect 186424 557534 186452 563654
rect 186424 557506 187096 557534
rect 187068 547963 187096 557506
rect 187712 552786 187740 566442
rect 189080 562352 189132 562358
rect 189080 562294 189132 562300
rect 187792 561128 187844 561134
rect 187792 561070 187844 561076
rect 187804 557534 187832 561070
rect 189092 557534 189120 562294
rect 190460 558272 190512 558278
rect 190460 558214 190512 558220
rect 190472 557534 190500 558214
rect 187804 557506 188568 557534
rect 189092 557506 189212 557534
rect 190472 557506 190684 557534
rect 187712 552758 187832 552786
rect 187804 547963 187832 552758
rect 188540 547963 188568 557506
rect 189184 547963 189212 557506
rect 189908 551472 189960 551478
rect 189908 551414 189960 551420
rect 189920 547963 189948 551414
rect 190656 547963 190684 557506
rect 191116 552770 191144 571338
rect 191840 569424 191892 569430
rect 191840 569366 191892 569372
rect 191852 557534 191880 569366
rect 191852 557506 192156 557534
rect 191380 555552 191432 555558
rect 191380 555494 191432 555500
rect 191104 552764 191156 552770
rect 191104 552706 191156 552712
rect 191392 547963 191420 555494
rect 192128 547963 192156 557506
rect 192496 549914 192524 572018
rect 193496 555756 193548 555762
rect 193496 555698 193548 555704
rect 192760 554124 192812 554130
rect 192760 554066 192812 554072
rect 192484 549908 192536 549914
rect 192484 549850 192536 549856
rect 192772 547963 192800 554066
rect 193508 547963 193536 555698
rect 193876 554062 193904 572086
rect 194600 567860 194652 567866
rect 194600 567802 194652 567808
rect 194612 557534 194640 567802
rect 194612 557506 195008 557534
rect 193864 554056 193916 554062
rect 193864 553998 193916 554004
rect 194232 549908 194284 549914
rect 194232 549850 194284 549856
rect 194244 547963 194272 549850
rect 194980 547963 195008 557506
rect 195256 550118 195284 575010
rect 195440 571402 195468 575062
rect 198004 572348 198056 572354
rect 198004 572290 198056 572296
rect 195428 571396 195480 571402
rect 195428 571338 195480 571344
rect 195980 565140 196032 565146
rect 195980 565082 196032 565088
rect 195992 557534 196020 565082
rect 197360 559700 197412 559706
rect 197360 559642 197412 559648
rect 197372 557534 197400 559642
rect 195992 557506 196388 557534
rect 197372 557506 197860 557534
rect 195612 550248 195664 550254
rect 195612 550190 195664 550196
rect 195244 550112 195296 550118
rect 195244 550054 195296 550060
rect 195624 547963 195652 550190
rect 196360 547963 196388 557506
rect 197084 554056 197136 554062
rect 197084 553998 197136 554004
rect 197096 547963 197124 553998
rect 197832 547963 197860 557506
rect 198016 555626 198044 572290
rect 198740 566704 198792 566710
rect 198740 566646 198792 566652
rect 198004 555620 198056 555626
rect 198004 555562 198056 555568
rect 198556 555484 198608 555490
rect 198556 555426 198608 555432
rect 198568 547963 198596 555426
rect 198752 552770 198780 566646
rect 198844 558210 198872 575062
rect 201512 572354 201540 575062
rect 201684 573504 201736 573510
rect 201684 573446 201736 573452
rect 201500 572348 201552 572354
rect 201500 572290 201552 572296
rect 200120 570852 200172 570858
rect 200120 570794 200172 570800
rect 198832 558204 198884 558210
rect 198832 558146 198884 558152
rect 199200 557048 199252 557054
rect 199200 556990 199252 556996
rect 198740 552764 198792 552770
rect 198740 552706 198792 552712
rect 199212 547963 199240 556990
rect 200132 552770 200160 570794
rect 200212 560992 200264 560998
rect 200212 560934 200264 560940
rect 200224 557534 200252 560934
rect 201696 557534 201724 573446
rect 204272 559638 204300 575062
rect 207032 572014 207060 575062
rect 210252 572150 210280 575062
rect 210240 572144 210292 572150
rect 210240 572086 210292 572092
rect 207020 572008 207072 572014
rect 207020 571950 207072 571956
rect 210712 565214 210740 637350
rect 211158 635216 211214 635225
rect 211158 635151 211214 635160
rect 210790 585440 210846 585449
rect 210790 585375 210846 585384
rect 210700 565208 210752 565214
rect 210700 565150 210752 565156
rect 210804 563922 210832 585375
rect 210882 580136 210938 580145
rect 210882 580071 210938 580080
rect 210792 563916 210844 563922
rect 210792 563858 210844 563864
rect 210056 563780 210108 563786
rect 210056 563722 210108 563728
rect 204352 562488 204404 562494
rect 204352 562430 204404 562436
rect 204260 559632 204312 559638
rect 204260 559574 204312 559580
rect 204364 557534 204392 562430
rect 207020 559768 207072 559774
rect 207020 559710 207072 559716
rect 205640 558204 205692 558210
rect 205640 558146 205692 558152
rect 200224 557506 200712 557534
rect 201696 557506 202184 557534
rect 204364 557506 205036 557534
rect 199936 552764 199988 552770
rect 199936 552706 199988 552712
rect 200120 552764 200172 552770
rect 200120 552706 200172 552712
rect 199948 547963 199976 552706
rect 200684 547963 200712 557506
rect 201408 552764 201460 552770
rect 201408 552706 201460 552712
rect 201420 547963 201448 552706
rect 202156 547963 202184 557506
rect 202788 551404 202840 551410
rect 202788 551346 202840 551352
rect 202800 547963 202828 551346
rect 203524 550384 203576 550390
rect 203524 550326 203576 550332
rect 203536 547963 203564 550326
rect 204260 550316 204312 550322
rect 204260 550258 204312 550264
rect 204272 547963 204300 550258
rect 205008 547963 205036 557506
rect 205652 547963 205680 558146
rect 207032 557534 207060 559710
rect 210068 557534 210096 563722
rect 207032 557506 207888 557534
rect 210068 557506 210740 557534
rect 206376 556980 206428 556986
rect 206376 556922 206428 556928
rect 206388 547963 206416 556922
rect 207112 551540 207164 551546
rect 207112 551482 207164 551488
rect 207124 547963 207152 551482
rect 207860 547963 207888 557506
rect 208584 552764 208636 552770
rect 208584 552706 208636 552712
rect 208596 547963 208624 552706
rect 209228 550520 209280 550526
rect 209228 550462 209280 550468
rect 209240 547963 209268 550462
rect 209964 550452 210016 550458
rect 209964 550394 210016 550400
rect 209976 547963 210004 550394
rect 210712 547963 210740 557506
rect 210896 552838 210924 580071
rect 210974 576872 211030 576881
rect 210974 576807 211030 576816
rect 210988 556918 211016 576807
rect 211172 570790 211200 635151
rect 212538 628280 212594 628289
rect 212538 628215 212594 628224
rect 211250 625696 211306 625705
rect 211250 625631 211306 625640
rect 211160 570784 211212 570790
rect 211160 570726 211212 570732
rect 211264 567934 211292 625631
rect 211434 619712 211490 619721
rect 211434 619647 211490 619656
rect 211342 616040 211398 616049
rect 211342 615975 211398 615984
rect 211356 568002 211384 615975
rect 211448 573578 211476 619647
rect 211710 601080 211766 601089
rect 211710 601015 211766 601024
rect 211618 597680 211674 597689
rect 211618 597615 211674 597624
rect 211526 594960 211582 594969
rect 211526 594895 211582 594904
rect 211436 573572 211488 573578
rect 211436 573514 211488 573520
rect 211344 567996 211396 568002
rect 211344 567938 211396 567944
rect 211252 567928 211304 567934
rect 211252 567870 211304 567876
rect 211160 565208 211212 565214
rect 211160 565150 211212 565156
rect 210976 556912 211028 556918
rect 210976 556854 211028 556860
rect 211172 552838 211200 565150
rect 210884 552832 210936 552838
rect 210884 552774 210936 552780
rect 211160 552832 211212 552838
rect 211160 552774 211212 552780
rect 211436 552016 211488 552022
rect 211436 551958 211488 551964
rect 211448 547963 211476 551958
rect 211540 551342 211568 594895
rect 211632 561066 211660 597615
rect 211724 566642 211752 601015
rect 211802 592376 211858 592385
rect 211802 592311 211858 592320
rect 211816 574938 211844 592311
rect 211804 574932 211856 574938
rect 211804 574874 211856 574880
rect 211712 566636 211764 566642
rect 211712 566578 211764 566584
rect 212552 562426 212580 628215
rect 212644 575006 212672 640358
rect 215944 639056 215996 639062
rect 215944 638998 215996 639004
rect 214564 637764 214616 637770
rect 214564 637706 214616 637712
rect 213920 636880 213972 636886
rect 213920 636822 213972 636828
rect 212814 632496 212870 632505
rect 212814 632431 212870 632440
rect 212722 622432 212778 622441
rect 212722 622367 212778 622376
rect 212632 575000 212684 575006
rect 212632 574942 212684 574948
rect 212736 565282 212764 622367
rect 212828 575074 212856 632431
rect 213090 613320 213146 613329
rect 213090 613255 213146 613264
rect 212906 610056 212962 610065
rect 212906 609991 212962 610000
rect 212816 575068 212868 575074
rect 212816 575010 212868 575016
rect 212724 565276 212776 565282
rect 212724 565218 212776 565224
rect 212540 562420 212592 562426
rect 212540 562362 212592 562368
rect 211620 561060 211672 561066
rect 211620 561002 211672 561008
rect 212920 555694 212948 609991
rect 212998 607336 213054 607345
rect 212998 607271 213054 607280
rect 213012 563854 213040 607271
rect 213104 569294 213132 613255
rect 213182 589656 213238 589665
rect 213182 589591 213238 589600
rect 213196 569362 213224 589591
rect 213274 582720 213330 582729
rect 213274 582655 213330 582664
rect 213288 572082 213316 582655
rect 213276 572076 213328 572082
rect 213276 572018 213328 572024
rect 213184 569356 213236 569362
rect 213184 569298 213236 569304
rect 213092 569288 213144 569294
rect 213092 569230 213144 569236
rect 213000 563848 213052 563854
rect 213000 563790 213052 563796
rect 213932 557534 213960 636822
rect 214010 603800 214066 603809
rect 214010 603735 214066 603744
rect 214024 575414 214052 603735
rect 214012 575408 214064 575414
rect 214012 575350 214064 575356
rect 213932 557506 214328 557534
rect 212908 555688 212960 555694
rect 212908 555630 212960 555636
rect 212172 552832 212224 552838
rect 212172 552774 212224 552780
rect 213552 552832 213604 552838
rect 213552 552774 213604 552780
rect 211528 551336 211580 551342
rect 211528 551278 211580 551284
rect 212184 547963 212212 552774
rect 212816 550112 212868 550118
rect 212816 550054 212868 550060
rect 212828 547963 212856 550054
rect 213564 547963 213592 552774
rect 214300 547963 214328 557506
rect 214576 550390 214604 637706
rect 214656 601724 214708 601730
rect 214656 601666 214708 601672
rect 214668 552022 214696 601666
rect 214748 586560 214800 586566
rect 214748 586502 214800 586508
rect 214760 559706 214788 586502
rect 215300 570784 215352 570790
rect 215300 570726 215352 570732
rect 214748 559700 214800 559706
rect 214748 559642 214800 559648
rect 215312 557534 215340 570726
rect 215312 557506 215892 557534
rect 215760 556232 215812 556238
rect 215760 556174 215812 556180
rect 214656 552016 214708 552022
rect 214656 551958 214708 551964
rect 214564 550384 214616 550390
rect 214564 550326 214616 550332
rect 215024 550180 215076 550186
rect 215024 550122 215076 550128
rect 215036 547963 215064 550122
rect 215772 547963 215800 556174
rect 215864 550066 215892 557506
rect 215956 550254 215984 638998
rect 216036 637968 216088 637974
rect 216036 637910 216088 637916
rect 216048 550526 216076 637910
rect 217324 637696 217376 637702
rect 217324 637638 217376 637644
rect 216128 626612 216180 626618
rect 216128 626554 216180 626560
rect 216140 557054 216168 626554
rect 216680 576904 216732 576910
rect 216680 576846 216732 576852
rect 216128 557048 216180 557054
rect 216128 556990 216180 556996
rect 216692 552786 216720 576846
rect 216772 559632 216824 559638
rect 216772 559574 216824 559580
rect 216784 557534 216812 559574
rect 216784 557506 217272 557534
rect 216692 552758 217180 552786
rect 216036 550520 216088 550526
rect 216036 550462 216088 550468
rect 215944 550248 215996 550254
rect 215944 550190 215996 550196
rect 215864 550038 216444 550066
rect 216416 547963 216444 550038
rect 217152 547963 217180 552758
rect 217244 550202 217272 557506
rect 217336 550322 217364 637638
rect 217428 556238 217456 640562
rect 223580 639872 223632 639878
rect 223580 639814 223632 639820
rect 222200 639804 222252 639810
rect 222200 639746 222252 639752
rect 220084 637832 220136 637838
rect 220084 637774 220136 637780
rect 218060 616888 218112 616894
rect 218060 616830 218112 616836
rect 217416 556232 217468 556238
rect 217416 556174 217468 556180
rect 218072 552786 218100 616830
rect 218152 579692 218204 579698
rect 218152 579634 218204 579640
rect 218164 557534 218192 579634
rect 219440 572076 219492 572082
rect 219440 572018 219492 572024
rect 218164 557506 219296 557534
rect 218072 552758 218652 552786
rect 217324 550316 217376 550322
rect 217324 550258 217376 550264
rect 217244 550174 217916 550202
rect 217888 547963 217916 550174
rect 218624 547963 218652 552758
rect 219268 547963 219296 557506
rect 219452 552634 219480 572018
rect 219440 552628 219492 552634
rect 219440 552570 219492 552576
rect 219992 550588 220044 550594
rect 219992 550530 220044 550536
rect 220004 547963 220032 550530
rect 220096 550458 220124 637774
rect 220176 607232 220228 607238
rect 220176 607174 220228 607180
rect 220188 559774 220216 607174
rect 220820 572348 220872 572354
rect 220820 572290 220872 572296
rect 220176 559768 220228 559774
rect 220176 559710 220228 559716
rect 220832 557534 220860 572290
rect 220832 557506 221504 557534
rect 220728 552628 220780 552634
rect 220728 552570 220780 552576
rect 220084 550452 220136 550458
rect 220084 550394 220136 550400
rect 220740 547963 220768 552570
rect 221476 547963 221504 557506
rect 222212 552838 222240 639746
rect 222844 622464 222896 622470
rect 222844 622406 222896 622412
rect 222292 572008 222344 572014
rect 222292 571950 222344 571956
rect 222200 552832 222252 552838
rect 222200 552774 222252 552780
rect 222304 548162 222332 571950
rect 222856 558278 222884 622406
rect 222844 558272 222896 558278
rect 222844 558214 222896 558220
rect 222844 552832 222896 552838
rect 222844 552774 222896 552780
rect 222228 548134 222332 548162
rect 222228 547944 222256 548134
rect 222856 547963 222884 552774
rect 223592 547963 223620 639814
rect 223672 619676 223724 619682
rect 223672 619618 223724 619624
rect 223684 557534 223712 619618
rect 223684 557506 224356 557534
rect 224328 547963 224356 557506
rect 226352 552786 226380 640766
rect 231124 640552 231176 640558
rect 231124 640494 231176 640500
rect 228364 638036 228416 638042
rect 228364 637978 228416 637984
rect 226984 637900 227036 637906
rect 226984 637842 227036 637848
rect 226432 583772 226484 583778
rect 226432 583714 226484 583720
rect 226444 557534 226472 583714
rect 226444 557506 226932 557534
rect 226352 552758 226472 552786
rect 225052 550384 225104 550390
rect 225052 550326 225104 550332
rect 225064 547963 225092 550326
rect 225788 550248 225840 550254
rect 225788 550190 225840 550196
rect 225800 547963 225828 550190
rect 226444 547963 226472 552758
rect 226904 549794 226932 557506
rect 226996 549914 227024 637842
rect 227720 574932 227772 574938
rect 227720 574874 227772 574880
rect 227732 552838 227760 574874
rect 227812 572212 227864 572218
rect 227812 572154 227864 572160
rect 227824 557534 227852 572154
rect 227824 557506 227944 557534
rect 227720 552832 227772 552838
rect 227720 552774 227772 552780
rect 226984 549908 227036 549914
rect 226984 549850 227036 549856
rect 226904 549766 227208 549794
rect 227180 547963 227208 549766
rect 227916 547963 227944 557506
rect 228376 550594 228404 637978
rect 229744 597576 229796 597582
rect 229744 597518 229796 597524
rect 229100 573640 229152 573646
rect 229100 573582 229152 573588
rect 229112 557534 229140 573582
rect 229112 557506 229324 557534
rect 228640 552832 228692 552838
rect 228640 552774 228692 552780
rect 228364 550588 228416 550594
rect 228364 550530 228416 550536
rect 228652 547963 228680 552774
rect 229296 547963 229324 557506
rect 229756 551546 229784 597518
rect 230480 572280 230532 572286
rect 230480 572222 230532 572228
rect 230492 557534 230520 572222
rect 230492 557506 230980 557534
rect 229744 551540 229796 551546
rect 229744 551482 229796 551488
rect 230020 550588 230072 550594
rect 230020 550530 230072 550536
rect 230032 547963 230060 550530
rect 230756 550316 230808 550322
rect 230756 550258 230808 550264
rect 230768 547963 230796 550258
rect 230952 549930 230980 557506
rect 231136 550594 231164 640494
rect 231216 639192 231268 639198
rect 231216 639134 231268 639140
rect 231124 550588 231176 550594
rect 231124 550530 231176 550536
rect 231228 550050 231256 639134
rect 232504 635180 232556 635186
rect 232504 635122 232556 635128
rect 231860 594856 231912 594862
rect 231860 594798 231912 594804
rect 231872 552770 231900 594798
rect 231952 572144 232004 572150
rect 231952 572086 232004 572092
rect 231964 557534 231992 572086
rect 231964 557506 232268 557534
rect 231860 552764 231912 552770
rect 231860 552706 231912 552712
rect 231216 550044 231268 550050
rect 231216 549986 231268 549992
rect 230952 549902 231532 549930
rect 231504 547963 231532 549902
rect 232240 547963 232268 557506
rect 232516 555762 232544 635122
rect 232504 555756 232556 555762
rect 232504 555698 232556 555704
rect 233252 552770 233280 641106
rect 238024 641028 238076 641034
rect 238024 640970 238076 640976
rect 235264 640892 235316 640898
rect 235264 640834 235316 640840
rect 233332 629332 233384 629338
rect 233332 629274 233384 629280
rect 233344 557534 233372 629274
rect 233884 589348 233936 589354
rect 233884 589290 233936 589296
rect 233896 561202 233924 589290
rect 233884 561196 233936 561202
rect 233884 561138 233936 561144
rect 233344 557506 233648 557534
rect 232872 552764 232924 552770
rect 232872 552706 232924 552712
rect 233240 552764 233292 552770
rect 233240 552706 233292 552712
rect 232884 547963 232912 552706
rect 233620 547963 233648 557506
rect 235276 552906 235304 640834
rect 236644 640688 236696 640694
rect 236644 640630 236696 640636
rect 235448 604512 235500 604518
rect 235448 604454 235500 604460
rect 235356 592068 235408 592074
rect 235356 592010 235408 592016
rect 235368 554198 235396 592010
rect 235460 568070 235488 604454
rect 235540 572416 235592 572422
rect 235540 572358 235592 572364
rect 235448 568064 235500 568070
rect 235448 568006 235500 568012
rect 235356 554192 235408 554198
rect 235356 554134 235408 554140
rect 235264 552900 235316 552906
rect 235264 552842 235316 552848
rect 234344 552764 234396 552770
rect 234344 552706 234396 552712
rect 234356 547963 234384 552706
rect 235080 550588 235132 550594
rect 235080 550530 235132 550536
rect 235092 547963 235120 550530
rect 235552 550390 235580 572358
rect 236656 550594 236684 640630
rect 237380 640484 237432 640490
rect 237380 640426 237432 640432
rect 236736 638104 236788 638110
rect 236736 638046 236788 638052
rect 236644 550588 236696 550594
rect 236644 550530 236696 550536
rect 235540 550384 235592 550390
rect 235540 550326 235592 550332
rect 236748 550186 236776 638046
rect 237392 636886 237420 640426
rect 238036 637634 238064 640970
rect 239496 640960 239548 640966
rect 239496 640902 239548 640908
rect 257436 640960 257488 640966
rect 257436 640902 257488 640908
rect 238116 640416 238168 640422
rect 238116 640358 238168 640364
rect 238024 637628 238076 637634
rect 238024 637570 238076 637576
rect 237380 636880 237432 636886
rect 237380 636822 237432 636828
rect 237378 635760 237434 635769
rect 237378 635695 237434 635704
rect 237392 635186 237420 635695
rect 237380 635180 237432 635186
rect 237380 635122 237432 635128
rect 237378 629504 237434 629513
rect 237378 629439 237434 629448
rect 237392 629338 237420 629439
rect 237380 629332 237432 629338
rect 237380 629274 237432 629280
rect 237378 626784 237434 626793
rect 237378 626719 237434 626728
rect 237392 626618 237420 626719
rect 237380 626612 237432 626618
rect 237380 626554 237432 626560
rect 237378 623384 237434 623393
rect 237378 623319 237434 623328
rect 237392 622470 237420 623319
rect 237380 622464 237432 622470
rect 237380 622406 237432 622412
rect 237378 620664 237434 620673
rect 237378 620599 237434 620608
rect 237392 619682 237420 620599
rect 237380 619676 237432 619682
rect 237380 619618 237432 619624
rect 237378 617264 237434 617273
rect 237378 617199 237434 617208
rect 237392 616894 237420 617199
rect 237380 616888 237432 616894
rect 237380 616830 237432 616836
rect 238036 611153 238064 637570
rect 238022 611144 238078 611153
rect 238022 611079 238078 611088
rect 237378 608424 237434 608433
rect 237378 608359 237434 608368
rect 237392 607238 237420 608359
rect 237380 607232 237432 607238
rect 237380 607174 237432 607180
rect 237378 605024 237434 605033
rect 237378 604959 237434 604968
rect 237392 604518 237420 604959
rect 237380 604512 237432 604518
rect 237380 604454 237432 604460
rect 237378 602304 237434 602313
rect 237378 602239 237434 602248
rect 237392 601730 237420 602239
rect 237380 601724 237432 601730
rect 237380 601666 237432 601672
rect 237378 598904 237434 598913
rect 237378 598839 237434 598848
rect 237392 597582 237420 598839
rect 237380 597576 237432 597582
rect 237380 597518 237432 597524
rect 237378 596184 237434 596193
rect 237378 596119 237434 596128
rect 237392 594862 237420 596119
rect 237380 594856 237432 594862
rect 237380 594798 237432 594804
rect 237378 592784 237434 592793
rect 237378 592719 237434 592728
rect 237392 592074 237420 592719
rect 237380 592068 237432 592074
rect 237380 592010 237432 592016
rect 237378 590064 237434 590073
rect 237378 589999 237434 590008
rect 237392 589354 237420 589999
rect 237380 589348 237432 589354
rect 237380 589290 237432 589296
rect 237378 586664 237434 586673
rect 237378 586599 237434 586608
rect 237392 586566 237420 586599
rect 237380 586560 237432 586566
rect 237380 586502 237432 586508
rect 237378 583944 237434 583953
rect 237378 583879 237434 583888
rect 237392 583778 237420 583879
rect 237380 583772 237432 583778
rect 237380 583714 237432 583720
rect 237378 580544 237434 580553
rect 237378 580479 237434 580488
rect 237392 579698 237420 580479
rect 237380 579692 237432 579698
rect 237380 579634 237432 579640
rect 237378 577824 237434 577833
rect 237378 577759 237434 577768
rect 237392 576910 237420 577759
rect 237380 576904 237432 576910
rect 237380 576846 237432 576852
rect 237932 552084 237984 552090
rect 237932 552026 237984 552032
rect 236736 550180 236788 550186
rect 236736 550122 236788 550128
rect 237196 549908 237248 549914
rect 237196 549850 237248 549856
rect 235816 548140 235868 548146
rect 235816 548082 235868 548088
rect 236460 548140 236512 548146
rect 236460 548082 236512 548088
rect 235828 547963 235856 548082
rect 236472 547963 236500 548082
rect 237208 547963 237236 549850
rect 237944 547963 237972 552026
rect 238128 551478 238156 640358
rect 238944 639260 238996 639266
rect 238944 639202 238996 639208
rect 238208 637628 238260 637634
rect 238208 637570 238260 637576
rect 238116 551472 238168 551478
rect 238116 551414 238168 551420
rect 238220 549982 238248 637570
rect 238298 632904 238354 632913
rect 238298 632839 238354 632848
rect 238312 552838 238340 632839
rect 238852 630012 238904 630018
rect 238852 629954 238904 629960
rect 238864 569430 238892 629954
rect 238956 614553 238984 639202
rect 239036 639124 239088 639130
rect 239036 639066 239088 639072
rect 238942 614544 238998 614553
rect 238942 614479 238998 614488
rect 238852 569424 238904 569430
rect 238852 569366 238904 569372
rect 239048 557534 239076 639066
rect 239404 637560 239456 637566
rect 239404 637502 239456 637508
rect 239416 562494 239444 637502
rect 239508 566710 239536 640902
rect 239588 640756 239640 640762
rect 239588 640698 239640 640704
rect 239600 570858 239628 640698
rect 254860 640620 254912 640626
rect 254860 640562 254912 640568
rect 243544 640552 243596 640558
rect 243544 640494 243596 640500
rect 249708 640552 249760 640558
rect 249708 640494 249760 640500
rect 243556 640354 243584 640494
rect 243544 640348 243596 640354
rect 243544 640290 243596 640296
rect 249064 640348 249116 640354
rect 249064 640290 249116 640296
rect 245660 638104 245712 638110
rect 245712 638052 245870 638058
rect 245660 638046 245870 638052
rect 245672 638030 245870 638046
rect 249076 638044 249104 640290
rect 249720 639878 249748 640494
rect 251640 640416 251692 640422
rect 251640 640358 251692 640364
rect 249708 639872 249760 639878
rect 249708 639814 249760 639820
rect 251652 638044 251680 640358
rect 254872 638044 254900 640562
rect 255320 640348 255372 640354
rect 255320 640290 255372 640296
rect 255332 639810 255360 640290
rect 255320 639804 255372 639810
rect 255320 639746 255372 639752
rect 257448 638044 257476 640902
rect 292212 640892 292264 640898
rect 292212 640834 292264 640840
rect 274824 640756 274876 640762
rect 274824 640698 274876 640704
rect 263232 640348 263284 640354
rect 263232 640290 263284 640296
rect 263244 638044 263272 640290
rect 272248 639192 272300 639198
rect 272248 639134 272300 639140
rect 269028 639056 269080 639062
rect 269028 638998 269080 639004
rect 266280 638042 266478 638058
rect 269040 638044 269068 638998
rect 272260 638044 272288 639134
rect 274836 638044 274864 640698
rect 289636 640484 289688 640490
rect 289636 640426 289688 640432
rect 289648 638044 289676 640426
rect 292224 638044 292252 640834
rect 300584 640824 300636 640830
rect 300584 640766 300636 640772
rect 295432 640552 295484 640558
rect 295432 640494 295484 640500
rect 295444 638044 295472 640494
rect 300596 638044 300624 640766
rect 266268 638036 266478 638042
rect 266320 638030 266478 638036
rect 266268 637978 266320 637984
rect 260380 637968 260432 637974
rect 260432 637916 260682 637922
rect 260380 637910 260682 637916
rect 260392 637894 260682 637910
rect 283576 637906 283866 637922
rect 283564 637900 283866 637906
rect 283616 637894 283866 637900
rect 283564 637842 283616 637848
rect 280252 637832 280304 637838
rect 280304 637780 280646 637786
rect 280252 637774 280646 637780
rect 280264 637758 280646 637774
rect 286152 637770 286442 637786
rect 286140 637764 286442 637770
rect 286192 637758 286442 637764
rect 286140 637706 286192 637712
rect 297732 637696 297784 637702
rect 242912 637622 243294 637650
rect 277688 637634 278070 637650
rect 297784 637644 298034 637650
rect 297732 637638 298034 637644
rect 277676 637628 278070 637634
rect 242912 637566 242940 637622
rect 277728 637622 278070 637628
rect 297744 637622 298034 637638
rect 277676 637570 277728 637576
rect 242900 637560 242952 637566
rect 242900 637502 242952 637508
rect 239784 637350 240074 637378
rect 239784 630018 239812 637350
rect 300858 635216 300914 635225
rect 300858 635151 300914 635160
rect 239772 630012 239824 630018
rect 239772 629954 239824 629960
rect 300674 576872 300730 576881
rect 300674 576807 300730 576816
rect 289820 575340 289872 575346
rect 289820 575282 289872 575288
rect 288532 575204 288584 575210
rect 288532 575146 288584 575152
rect 288440 575136 288492 575142
rect 240060 572354 240088 575076
rect 241532 575062 242650 575090
rect 244292 575062 245226 575090
rect 240048 572348 240100 572354
rect 240048 572290 240100 572296
rect 239588 570852 239640 570858
rect 239588 570794 239640 570800
rect 240140 569288 240192 569294
rect 240140 569230 240192 569236
rect 239496 566704 239548 566710
rect 239496 566646 239548 566652
rect 239404 562488 239456 562494
rect 239404 562430 239456 562436
rect 240152 557534 240180 569230
rect 239048 557506 239444 557534
rect 240152 557506 240824 557534
rect 238300 552832 238352 552838
rect 238300 552774 238352 552780
rect 238666 550080 238722 550089
rect 238666 550015 238722 550024
rect 238208 549976 238260 549982
rect 238208 549918 238260 549924
rect 238680 547963 238708 550015
rect 239416 547963 239444 557506
rect 240048 549500 240100 549506
rect 240048 549442 240100 549448
rect 240060 547963 240088 549442
rect 240796 547963 240824 557506
rect 241532 550254 241560 575062
rect 244292 565350 244320 575062
rect 245660 573572 245712 573578
rect 245660 573514 245712 573520
rect 244464 567928 244516 567934
rect 244464 567870 244516 567876
rect 244280 565344 244332 565350
rect 244280 565286 244332 565292
rect 242900 558272 242952 558278
rect 242900 558214 242952 558220
rect 241612 552152 241664 552158
rect 241612 552094 241664 552100
rect 241520 550248 241572 550254
rect 241520 550190 241572 550196
rect 241624 548162 241652 552094
rect 242256 550180 242308 550186
rect 242256 550122 242308 550128
rect 241548 548134 241652 548162
rect 241548 547944 241576 548134
rect 242268 547963 242296 550122
rect 242912 547963 242940 558214
rect 244476 557534 244504 567870
rect 245672 557534 245700 573514
rect 248432 572422 248460 575076
rect 248420 572416 248472 572422
rect 248420 572358 248472 572364
rect 249064 572348 249116 572354
rect 249064 572290 249116 572296
rect 246304 571532 246356 571538
rect 246304 571474 246356 571480
rect 244476 557506 245148 557534
rect 245672 557506 245884 557534
rect 244372 551540 244424 551546
rect 244372 551482 244424 551488
rect 243636 548344 243688 548350
rect 243636 548286 243688 548292
rect 243648 547963 243676 548286
rect 244384 547963 244412 551482
rect 245120 547963 245148 557506
rect 245856 547963 245884 557506
rect 246316 550322 246344 571474
rect 247040 566636 247092 566642
rect 247040 566578 247092 566584
rect 247052 557534 247080 566578
rect 247052 557506 248000 557534
rect 246488 552764 246540 552770
rect 246488 552706 246540 552712
rect 246304 550316 246356 550322
rect 246304 550258 246356 550264
rect 246500 547963 246528 552706
rect 247224 548412 247276 548418
rect 247224 548354 247276 548360
rect 247236 547963 247264 548354
rect 247972 547963 248000 557506
rect 249076 550118 249104 572290
rect 251008 571538 251036 575076
rect 253952 575062 254242 575090
rect 250996 571532 251048 571538
rect 250996 571474 251048 571480
rect 253952 561134 253980 575062
rect 255320 569356 255372 569362
rect 255320 569298 255372 569304
rect 253940 561128 253992 561134
rect 253940 561070 253992 561076
rect 249800 561060 249852 561066
rect 249800 561002 249852 561008
rect 249812 557534 249840 561002
rect 249812 557506 250852 557534
rect 250076 556912 250128 556918
rect 250076 556854 250128 556860
rect 249432 551472 249484 551478
rect 249432 551414 249484 551420
rect 249064 550112 249116 550118
rect 249064 550054 249116 550060
rect 248694 549672 248750 549681
rect 248694 549607 248750 549616
rect 248708 547963 248736 549607
rect 249444 547963 249472 551414
rect 250088 547963 250116 556854
rect 250824 547963 250852 557506
rect 251548 555620 251600 555626
rect 251548 555562 251600 555568
rect 251560 547963 251588 555562
rect 253664 554192 253716 554198
rect 253664 554134 253716 554140
rect 252284 552220 252336 552226
rect 252284 552162 252336 552168
rect 252296 547963 252324 552162
rect 252928 550044 252980 550050
rect 252928 549986 252980 549992
rect 252940 547963 252968 549986
rect 253676 547963 253704 554134
rect 255332 552838 255360 569298
rect 256804 567194 256832 575076
rect 260024 572286 260052 575076
rect 262232 575062 262614 575090
rect 288440 575078 288492 575084
rect 260840 575000 260892 575006
rect 260840 574942 260892 574948
rect 260012 572280 260064 572286
rect 260012 572222 260064 572228
rect 256712 567166 256832 567194
rect 255320 552832 255372 552838
rect 255320 552774 255372 552780
rect 256516 552832 256568 552838
rect 256516 552774 256568 552780
rect 254400 551132 254452 551138
rect 254400 551074 254452 551080
rect 254412 547963 254440 551074
rect 255872 550724 255924 550730
rect 255872 550666 255924 550672
rect 255134 549808 255190 549817
rect 255134 549743 255190 549752
rect 255148 547963 255176 549743
rect 255884 547963 255912 550666
rect 256528 547963 256556 552774
rect 256712 551410 256740 567166
rect 256792 561128 256844 561134
rect 256792 561070 256844 561076
rect 256804 552838 256832 561070
rect 259460 559700 259512 559706
rect 259460 559642 259512 559648
rect 259472 557534 259500 559642
rect 260852 557534 260880 574942
rect 259472 557506 260144 557534
rect 260852 557506 261616 557534
rect 259460 554260 259512 554266
rect 259460 554202 259512 554208
rect 256792 552832 256844 552838
rect 256792 552774 256844 552780
rect 257988 552832 258040 552838
rect 257988 552774 258040 552780
rect 256700 551404 256752 551410
rect 256700 551346 256752 551352
rect 257252 549568 257304 549574
rect 257252 549510 257304 549516
rect 257264 547963 257292 549510
rect 258000 547963 258028 552774
rect 258724 552288 258776 552294
rect 258724 552230 258776 552236
rect 258736 547963 258764 552230
rect 259472 547963 259500 554202
rect 260116 547963 260144 557506
rect 260840 548208 260892 548214
rect 260840 548150 260892 548156
rect 260852 547963 260880 548150
rect 261588 547963 261616 557506
rect 262232 556986 262260 575062
rect 265820 572218 265848 575076
rect 265808 572212 265860 572218
rect 265808 572154 265860 572160
rect 268396 572082 268424 575076
rect 271616 572354 271644 575076
rect 271604 572348 271656 572354
rect 271604 572290 271656 572296
rect 273904 572212 273956 572218
rect 273904 572154 273956 572160
rect 268384 572076 268436 572082
rect 268384 572018 268436 572024
rect 269120 572076 269172 572082
rect 269120 572018 269172 572024
rect 267740 567248 267792 567254
rect 267740 567190 267792 567196
rect 263600 563916 263652 563922
rect 263600 563858 263652 563864
rect 263612 557534 263640 563858
rect 267752 557534 267780 567190
rect 263612 557506 263732 557534
rect 267752 557506 268056 557534
rect 262220 556980 262272 556986
rect 262220 556922 262272 556928
rect 262312 551268 262364 551274
rect 262312 551210 262364 551216
rect 262324 547963 262352 551210
rect 263048 548276 263100 548282
rect 263048 548218 263100 548224
rect 263060 547963 263088 548218
rect 263704 547963 263732 557506
rect 266544 556980 266596 556986
rect 266544 556922 266596 556928
rect 264428 551200 264480 551206
rect 264428 551142 264480 551148
rect 264440 547963 264468 551142
rect 265900 550860 265952 550866
rect 265900 550802 265952 550808
rect 265164 548684 265216 548690
rect 265164 548626 265216 548632
rect 265176 547963 265204 548626
rect 265912 547963 265940 550802
rect 266556 547963 266584 556922
rect 267280 552832 267332 552838
rect 267280 552774 267332 552780
rect 267292 547963 267320 552774
rect 268028 547963 268056 557506
rect 269132 552786 269160 572018
rect 269212 566704 269264 566710
rect 269212 566646 269264 566652
rect 269224 557534 269252 566646
rect 273260 563848 273312 563854
rect 273260 563790 273312 563796
rect 269224 557506 270172 557534
rect 269132 552758 269528 552786
rect 268752 548752 268804 548758
rect 268752 548694 268804 548700
rect 268764 547963 268792 548694
rect 269500 547963 269528 552758
rect 270144 547963 270172 557506
rect 273272 552634 273300 563790
rect 273916 559638 273944 572154
rect 274192 572014 274220 575076
rect 274180 572008 274232 572014
rect 274180 571950 274232 571956
rect 274640 565276 274692 565282
rect 274640 565218 274692 565224
rect 273904 559632 273956 559638
rect 273904 559574 273956 559580
rect 274652 557534 274680 565218
rect 274652 557506 275232 557534
rect 273260 552628 273312 552634
rect 273260 552570 273312 552576
rect 274456 552628 274508 552634
rect 274456 552570 274508 552576
rect 271604 551336 271656 551342
rect 271604 551278 271656 551284
rect 270868 550112 270920 550118
rect 270868 550054 270920 550060
rect 270880 547963 270908 550054
rect 271616 547963 271644 551278
rect 273720 551064 273772 551070
rect 273720 551006 273772 551012
rect 272340 550996 272392 551002
rect 272340 550938 272392 550944
rect 272352 547963 272380 550938
rect 273076 550928 273128 550934
rect 273076 550870 273128 550876
rect 273088 547963 273116 550870
rect 273260 549500 273312 549506
rect 273260 549442 273312 549448
rect 273272 548554 273300 549442
rect 273260 548548 273312 548554
rect 273260 548490 273312 548496
rect 273732 547963 273760 551006
rect 274468 547963 274496 552570
rect 275204 547963 275232 557506
rect 277412 555558 277440 575076
rect 279988 572150 280016 575076
rect 283208 572218 283236 575076
rect 283196 572212 283248 572218
rect 283196 572154 283248 572160
rect 279976 572144 280028 572150
rect 279976 572086 280028 572092
rect 280804 572144 280856 572150
rect 280804 572086 280856 572092
rect 280160 572008 280212 572014
rect 280160 571950 280212 571956
rect 277400 555552 277452 555558
rect 277400 555494 277452 555500
rect 279516 555552 279568 555558
rect 279516 555494 279568 555500
rect 275928 549704 275980 549710
rect 275928 549646 275980 549652
rect 275940 547963 275968 549646
rect 277308 549636 277360 549642
rect 277308 549578 277360 549584
rect 276572 548480 276624 548486
rect 276572 548422 276624 548428
rect 276584 547963 276612 548422
rect 277320 547963 277348 549578
rect 278044 549500 278096 549506
rect 278044 549442 278096 549448
rect 278056 547963 278084 549442
rect 278780 548616 278832 548622
rect 278780 548558 278832 548564
rect 278792 547963 278820 548558
rect 279528 547963 279556 555494
rect 280172 552786 280200 571950
rect 280816 554130 280844 572086
rect 285784 567194 285812 575076
rect 287060 575068 287112 575074
rect 287060 575010 287112 575016
rect 285692 567166 285812 567194
rect 281540 558340 281592 558346
rect 281540 558282 281592 558288
rect 281552 557534 281580 558282
rect 285692 558210 285720 567166
rect 285680 558204 285732 558210
rect 285680 558146 285732 558152
rect 281552 557506 282408 557534
rect 280804 554124 280856 554130
rect 280804 554066 280856 554072
rect 280172 552758 280936 552786
rect 280160 549772 280212 549778
rect 280160 549714 280212 549720
rect 280172 547963 280200 549714
rect 280908 547963 280936 552758
rect 281632 549296 281684 549302
rect 281632 549238 281684 549244
rect 281644 547963 281672 549238
rect 282380 547963 282408 557506
rect 283748 552900 283800 552906
rect 283748 552842 283800 552848
rect 283104 549840 283156 549846
rect 283104 549782 283156 549788
rect 283116 547963 283144 549782
rect 283760 547963 283788 552842
rect 287072 552786 287100 575010
rect 287704 572212 287756 572218
rect 287704 572154 287756 572160
rect 287716 555490 287744 572154
rect 287704 555484 287756 555490
rect 287704 555426 287756 555432
rect 288452 552786 288480 575078
rect 288544 557534 288572 575146
rect 288636 575062 289018 575090
rect 288636 562358 288664 575062
rect 288624 562352 288676 562358
rect 288624 562294 288676 562300
rect 289832 557534 289860 575282
rect 293960 575272 294012 575278
rect 293960 575214 294012 575220
rect 291304 575062 291594 575090
rect 291200 574728 291252 574734
rect 291200 574670 291252 574676
rect 288544 557506 289584 557534
rect 289832 557506 290228 557534
rect 287072 552758 288112 552786
rect 288452 552758 288848 552786
rect 286692 552560 286744 552566
rect 286692 552502 286744 552508
rect 285680 552492 285732 552498
rect 285680 552434 285732 552440
rect 285220 552356 285272 552362
rect 285220 552298 285272 552304
rect 284484 549432 284536 549438
rect 284484 549374 284536 549380
rect 284496 547963 284524 549374
rect 285232 547963 285260 552298
rect 285692 549914 285720 552434
rect 285956 552424 286008 552430
rect 285956 552366 286008 552372
rect 285680 549908 285732 549914
rect 285680 549850 285732 549856
rect 285968 547963 285996 552366
rect 286704 547963 286732 552502
rect 287336 550792 287388 550798
rect 287336 550734 287388 550740
rect 287348 547963 287376 550734
rect 288084 547963 288112 552758
rect 288820 547963 288848 552758
rect 289556 547963 289584 557506
rect 290200 547963 290228 557506
rect 290924 552968 290976 552974
rect 290924 552910 290976 552916
rect 290936 547963 290964 552910
rect 291212 552634 291240 574670
rect 291304 556850 291332 575062
rect 291292 556844 291344 556850
rect 291292 556786 291344 556792
rect 293972 552634 294000 575214
rect 294064 575062 294814 575090
rect 294064 566574 294092 575062
rect 296904 574660 296956 574666
rect 296904 574602 296956 574608
rect 294052 566568 294104 566574
rect 294052 566510 294104 566516
rect 296916 557534 296944 574602
rect 297376 572150 297404 575076
rect 300596 572218 300624 575076
rect 300584 572212 300636 572218
rect 300584 572154 300636 572160
rect 297364 572144 297416 572150
rect 297364 572086 297416 572092
rect 300688 559570 300716 576807
rect 300872 574802 300900 635151
rect 300950 632496 301006 632505
rect 300950 632431 301006 632440
rect 300964 574938 300992 632431
rect 302238 628280 302294 628289
rect 302238 628215 302294 628224
rect 301042 625696 301098 625705
rect 301042 625631 301098 625640
rect 300952 574932 301004 574938
rect 300952 574874 301004 574880
rect 301056 574870 301084 625631
rect 301134 619712 301190 619721
rect 301134 619647 301190 619656
rect 301044 574864 301096 574870
rect 301044 574806 301096 574812
rect 300860 574796 300912 574802
rect 300860 574738 300912 574744
rect 301148 570722 301176 619647
rect 301318 610056 301374 610065
rect 301318 609991 301374 610000
rect 301226 601080 301282 601089
rect 301226 601015 301282 601024
rect 301136 570716 301188 570722
rect 301136 570658 301188 570664
rect 300676 559564 300728 559570
rect 300676 559506 300728 559512
rect 296916 557506 297404 557534
rect 295340 552968 295392 552974
rect 295340 552910 295392 552916
rect 295352 552634 295380 552910
rect 291200 552628 291252 552634
rect 291200 552570 291252 552576
rect 292396 552628 292448 552634
rect 292396 552570 292448 552576
rect 293960 552628 294012 552634
rect 293960 552570 294012 552576
rect 295248 552628 295300 552634
rect 295248 552570 295300 552576
rect 295340 552628 295392 552634
rect 295340 552570 295392 552576
rect 291660 550656 291712 550662
rect 291660 550598 291712 550604
rect 291672 547963 291700 550598
rect 292408 547963 292436 552570
rect 294510 549536 294566 549545
rect 294510 549471 294566 549480
rect 293130 549400 293186 549409
rect 293130 549335 293186 549344
rect 293144 547963 293172 549335
rect 293776 548820 293828 548826
rect 293776 548762 293828 548768
rect 293788 547963 293816 548762
rect 294524 547963 294552 549471
rect 295260 547963 295288 552570
rect 295984 550248 296036 550254
rect 295984 550190 296036 550196
rect 295996 547963 296024 550190
rect 296720 549364 296772 549370
rect 296720 549306 296772 549312
rect 296732 547963 296760 549306
rect 297376 547963 297404 557506
rect 301240 552702 301268 601015
rect 301332 565214 301360 609991
rect 301410 592376 301466 592385
rect 301410 592311 301466 592320
rect 301424 569226 301452 592311
rect 301502 589656 301558 589665
rect 301502 589591 301558 589600
rect 301516 570790 301544 589591
rect 301594 582720 301650 582729
rect 301594 582655 301650 582664
rect 301608 573442 301636 582655
rect 302252 573510 302280 628215
rect 302330 622432 302386 622441
rect 302330 622367 302386 622376
rect 302240 573504 302292 573510
rect 302240 573446 302292 573452
rect 301596 573436 301648 573442
rect 301596 573378 301648 573384
rect 301504 570784 301556 570790
rect 301504 570726 301556 570732
rect 301412 569220 301464 569226
rect 301412 569162 301464 569168
rect 302344 566506 302372 622367
rect 302422 616040 302478 616049
rect 302422 615975 302478 615984
rect 302332 566500 302384 566506
rect 302332 566442 302384 566448
rect 301320 565208 301372 565214
rect 301320 565150 301372 565156
rect 302436 563718 302464 615975
rect 302514 613320 302570 613329
rect 302514 613255 302570 613264
rect 302528 565146 302556 613255
rect 302698 607336 302754 607345
rect 302698 607271 302754 607280
rect 302606 597680 302662 597689
rect 302606 597615 302662 597624
rect 302516 565140 302568 565146
rect 302516 565082 302568 565088
rect 302424 563712 302476 563718
rect 302424 563654 302476 563660
rect 302620 554062 302648 597615
rect 302712 563786 302740 607271
rect 302882 603800 302938 603809
rect 302882 603735 302938 603744
rect 303158 603800 303214 603809
rect 303158 603735 303160 603744
rect 302790 594960 302846 594969
rect 302790 594895 302846 594904
rect 302700 563780 302752 563786
rect 302700 563722 302752 563728
rect 302804 560998 302832 594895
rect 302896 575414 302924 603735
rect 303212 603735 303214 603744
rect 303160 603706 303212 603712
rect 304264 596216 304316 596222
rect 304264 596158 304316 596164
rect 302974 585440 303030 585449
rect 302974 585375 303030 585384
rect 302884 575408 302936 575414
rect 302884 575350 302936 575356
rect 302896 574122 302924 575350
rect 302884 574116 302936 574122
rect 302884 574058 302936 574064
rect 302988 567866 303016 585375
rect 303066 580136 303122 580145
rect 303066 580071 303122 580080
rect 303080 573646 303108 580071
rect 303344 574116 303396 574122
rect 303344 574058 303396 574064
rect 303068 573640 303120 573646
rect 303068 573582 303120 573588
rect 302976 567860 303028 567866
rect 302976 567802 303028 567808
rect 302792 560992 302844 560998
rect 302792 560934 302844 560940
rect 302608 554056 302660 554062
rect 302608 553998 302660 554004
rect 301228 552696 301280 552702
rect 301228 552638 301280 552644
rect 300124 551268 300176 551274
rect 300124 551210 300176 551216
rect 299572 549976 299624 549982
rect 298098 549944 298154 549953
rect 299572 549918 299624 549924
rect 298098 549879 298154 549888
rect 298836 549908 298888 549914
rect 298112 547963 298140 549879
rect 298836 549850 298888 549856
rect 298848 547963 298876 549850
rect 299584 547963 299612 549918
rect 300136 526250 300164 551210
rect 302884 551200 302936 551206
rect 302884 551142 302936 551148
rect 300676 550248 300728 550254
rect 300676 550190 300728 550196
rect 300308 549772 300360 549778
rect 300308 549714 300360 549720
rect 300216 549704 300268 549710
rect 300216 549646 300268 549652
rect 300228 527882 300256 549646
rect 300320 528222 300348 549714
rect 300398 549672 300454 549681
rect 300398 549607 300454 549616
rect 300412 528465 300440 549607
rect 300492 549432 300544 549438
rect 300492 549374 300544 549380
rect 300504 529786 300532 549374
rect 300584 549296 300636 549302
rect 300584 549238 300636 549244
rect 300596 529854 300624 549238
rect 300688 529922 300716 550190
rect 301686 550080 301742 550089
rect 301686 550015 301742 550024
rect 301596 549568 301648 549574
rect 301596 549510 301648 549516
rect 301502 549400 301558 549409
rect 301502 549335 301558 549344
rect 301044 548140 301096 548146
rect 301044 548082 301096 548088
rect 301056 543726 301084 548082
rect 301044 543720 301096 543726
rect 301044 543662 301096 543668
rect 300676 529916 300728 529922
rect 300676 529858 300728 529864
rect 300584 529848 300636 529854
rect 300584 529790 300636 529796
rect 300492 529780 300544 529786
rect 300492 529722 300544 529728
rect 300398 528456 300454 528465
rect 300398 528391 300454 528400
rect 300308 528216 300360 528222
rect 300308 528158 300360 528164
rect 300216 527876 300268 527882
rect 300216 527818 300268 527824
rect 300124 526244 300176 526250
rect 300124 526186 300176 526192
rect 301516 525774 301544 549335
rect 301608 528154 301636 549510
rect 301700 528329 301728 550015
rect 301872 549840 301924 549846
rect 301872 549782 301924 549788
rect 301780 548412 301832 548418
rect 301780 548354 301832 548360
rect 301686 528320 301742 528329
rect 301686 528255 301742 528264
rect 301596 528148 301648 528154
rect 301596 528090 301648 528096
rect 301792 526590 301820 548354
rect 301884 529718 301912 549782
rect 301964 548344 302016 548350
rect 301964 548286 302016 548292
rect 301976 539578 302004 548286
rect 302790 540424 302846 540433
rect 302790 540359 302846 540368
rect 302804 539646 302832 540359
rect 302792 539640 302844 539646
rect 302792 539582 302844 539588
rect 301964 539572 302016 539578
rect 301964 539514 302016 539520
rect 301872 529712 301924 529718
rect 301872 529654 301924 529660
rect 302896 526726 302924 551142
rect 302976 551132 303028 551138
rect 302976 551074 303028 551080
rect 302884 526720 302936 526726
rect 302884 526662 302936 526668
rect 301780 526584 301832 526590
rect 301780 526526 301832 526532
rect 302988 526522 303016 551074
rect 303160 550180 303212 550186
rect 303160 550122 303212 550128
rect 303068 548752 303120 548758
rect 303068 548694 303120 548700
rect 302976 526516 303028 526522
rect 302976 526458 303028 526464
rect 303080 526318 303108 548694
rect 303172 529650 303200 550122
rect 303160 529644 303212 529650
rect 303160 529586 303212 529592
rect 303068 526312 303120 526318
rect 303068 526254 303120 526260
rect 301504 525768 301556 525774
rect 301504 525710 301556 525716
rect 302882 525464 302938 525473
rect 302882 525399 302938 525408
rect 302896 524482 302924 525399
rect 302884 524476 302936 524482
rect 302884 524418 302936 524424
rect 57886 517984 57942 517993
rect 57886 517919 57942 517928
rect 57900 517546 57928 517919
rect 53748 517540 53800 517546
rect 53748 517482 53800 517488
rect 57888 517540 57940 517546
rect 57888 517482 57940 517488
rect 15844 486464 15896 486470
rect 15844 486406 15896 486412
rect 15856 411262 15884 486406
rect 50988 485308 51040 485314
rect 50988 485250 51040 485256
rect 42432 485172 42484 485178
rect 42432 485114 42484 485120
rect 42246 479496 42302 479505
rect 42246 479431 42302 479440
rect 42156 476876 42208 476882
rect 42156 476818 42208 476824
rect 42064 465996 42116 466002
rect 42064 465938 42116 465944
rect 15844 411256 15896 411262
rect 15844 411198 15896 411204
rect 42076 378078 42104 465938
rect 42168 379030 42196 476818
rect 42156 379024 42208 379030
rect 42156 378966 42208 378972
rect 42064 378072 42116 378078
rect 42064 378014 42116 378020
rect 42260 271561 42288 479431
rect 42338 476776 42394 476785
rect 42338 476711 42394 476720
rect 42246 271552 42302 271561
rect 42246 271487 42302 271496
rect 42352 268530 42380 476711
rect 42444 271862 42472 485114
rect 43628 485104 43680 485110
rect 43628 485046 43680 485052
rect 42614 480040 42670 480049
rect 42614 479975 42670 479984
rect 42524 467696 42576 467702
rect 42524 467638 42576 467644
rect 42432 271856 42484 271862
rect 42432 271798 42484 271804
rect 42340 268524 42392 268530
rect 42340 268466 42392 268472
rect 42536 166326 42564 467638
rect 42524 166320 42576 166326
rect 42524 166262 42576 166268
rect 42628 70378 42656 479975
rect 43534 476912 43590 476921
rect 43534 476847 43590 476856
rect 43444 467356 43496 467362
rect 43444 467298 43496 467304
rect 42706 467120 42762 467129
rect 42706 467055 42762 467064
rect 42616 70372 42668 70378
rect 42616 70314 42668 70320
rect 42720 57662 42748 467055
rect 43352 465928 43404 465934
rect 43352 465870 43404 465876
rect 43364 377466 43392 465870
rect 43352 377460 43404 377466
rect 43352 377402 43404 377408
rect 43456 270502 43484 467298
rect 43444 270496 43496 270502
rect 43444 270438 43496 270444
rect 43548 268394 43576 476847
rect 43640 273630 43668 485046
rect 50620 484968 50672 484974
rect 50620 484910 50672 484916
rect 50632 484537 50660 484910
rect 50896 484832 50948 484838
rect 50896 484774 50948 484780
rect 50908 484537 50936 484774
rect 50618 484528 50674 484537
rect 50618 484463 50674 484472
rect 50894 484528 50950 484537
rect 50894 484463 50950 484472
rect 50436 482996 50488 483002
rect 50436 482938 50488 482944
rect 48044 482928 48096 482934
rect 48044 482870 48096 482876
rect 47860 482792 47912 482798
rect 47860 482734 47912 482740
rect 46572 482724 46624 482730
rect 46572 482666 46624 482672
rect 46388 482588 46440 482594
rect 46388 482530 46440 482536
rect 45468 479936 45520 479942
rect 45468 479878 45520 479884
rect 43720 479868 43772 479874
rect 43720 479810 43772 479816
rect 43628 273624 43680 273630
rect 43628 273566 43680 273572
rect 43732 269006 43760 479810
rect 43810 479632 43866 479641
rect 43810 479567 43866 479576
rect 43720 269000 43772 269006
rect 43720 268942 43772 268948
rect 43824 268462 43852 479567
rect 45376 477420 45428 477426
rect 45376 477362 45428 477368
rect 44732 476808 44784 476814
rect 44732 476750 44784 476756
rect 43996 476604 44048 476610
rect 43996 476546 44048 476552
rect 43904 467492 43956 467498
rect 43904 467434 43956 467440
rect 43812 268456 43864 268462
rect 43812 268398 43864 268404
rect 43536 268388 43588 268394
rect 43536 268330 43588 268336
rect 43916 166394 43944 467434
rect 44008 175234 44036 476546
rect 44086 467256 44142 467265
rect 44086 467191 44142 467200
rect 43996 175228 44048 175234
rect 43996 175170 44048 175176
rect 43904 166388 43956 166394
rect 43904 166330 43956 166336
rect 42708 57656 42760 57662
rect 42708 57598 42760 57604
rect 44100 54534 44128 467191
rect 44640 416832 44692 416838
rect 44640 416774 44692 416780
rect 44652 380866 44680 416774
rect 44744 391950 44772 476750
rect 45100 467832 45152 467838
rect 45100 467774 45152 467780
rect 44824 467764 44876 467770
rect 44824 467706 44876 467712
rect 44732 391944 44784 391950
rect 44732 391886 44784 391892
rect 44640 380860 44692 380866
rect 44640 380802 44692 380808
rect 44836 273562 44864 467706
rect 45008 467424 45060 467430
rect 45008 467366 45060 467372
rect 44916 467288 44968 467294
rect 44916 467230 44968 467236
rect 44824 273556 44876 273562
rect 44824 273498 44876 273504
rect 44928 273494 44956 467230
rect 44916 273488 44968 273494
rect 44916 273430 44968 273436
rect 45020 273426 45048 467366
rect 45008 273420 45060 273426
rect 45008 273362 45060 273368
rect 45112 273358 45140 467774
rect 45284 467220 45336 467226
rect 45284 467162 45336 467168
rect 45192 467152 45244 467158
rect 45192 467094 45244 467100
rect 45100 273352 45152 273358
rect 45100 273294 45152 273300
rect 45204 273290 45232 467094
rect 45192 273284 45244 273290
rect 45192 273226 45244 273232
rect 45296 268802 45324 467162
rect 45284 268796 45336 268802
rect 45284 268738 45336 268744
rect 45388 267714 45416 477362
rect 45480 268938 45508 479878
rect 46112 479664 46164 479670
rect 46112 479606 46164 479612
rect 46020 469056 46072 469062
rect 46020 468998 46072 469004
rect 46032 383654 46060 468998
rect 46124 389094 46152 479606
rect 46296 476944 46348 476950
rect 46296 476886 46348 476892
rect 46204 471980 46256 471986
rect 46204 471922 46256 471928
rect 46112 389088 46164 389094
rect 46112 389030 46164 389036
rect 46032 383626 46152 383654
rect 46124 379273 46152 383626
rect 46110 379264 46166 379273
rect 46110 379199 46166 379208
rect 46124 270978 46152 379199
rect 46216 378622 46244 471922
rect 46308 379098 46336 476886
rect 46296 379092 46348 379098
rect 46296 379034 46348 379040
rect 46204 378616 46256 378622
rect 46204 378558 46256 378564
rect 46400 303618 46428 482530
rect 46480 482520 46532 482526
rect 46480 482462 46532 482468
rect 46388 303612 46440 303618
rect 46388 303554 46440 303560
rect 46492 300830 46520 482462
rect 46480 300824 46532 300830
rect 46480 300766 46532 300772
rect 46584 272406 46612 482666
rect 46846 482352 46902 482361
rect 46664 482316 46716 482322
rect 46846 482287 46902 482296
rect 46664 482258 46716 482264
rect 46676 273086 46704 482258
rect 46756 480140 46808 480146
rect 46756 480082 46808 480088
rect 46664 273080 46716 273086
rect 46664 273022 46716 273028
rect 46572 272400 46624 272406
rect 46572 272342 46624 272348
rect 46112 270972 46164 270978
rect 46112 270914 46164 270920
rect 45468 268932 45520 268938
rect 45468 268874 45520 268880
rect 46124 267734 46152 270914
rect 46386 268560 46442 268569
rect 46386 268495 46442 268504
rect 45376 267708 45428 267714
rect 46124 267706 46336 267734
rect 45376 267650 45428 267656
rect 46308 146266 46336 267706
rect 46400 164150 46428 268495
rect 46478 268424 46534 268433
rect 46478 268359 46534 268368
rect 46388 164144 46440 164150
rect 46388 164086 46440 164092
rect 46492 148714 46520 268359
rect 46480 148708 46532 148714
rect 46480 148650 46532 148656
rect 46296 146260 46348 146266
rect 46296 146202 46348 146208
rect 46584 145382 46612 272342
rect 46768 269074 46796 480082
rect 46756 269068 46808 269074
rect 46756 269010 46808 269016
rect 46664 268524 46716 268530
rect 46664 268466 46716 268472
rect 46676 148850 46704 268466
rect 46860 251190 46888 482287
rect 47676 479800 47728 479806
rect 47676 479742 47728 479748
rect 47584 479596 47636 479602
rect 47584 479538 47636 479544
rect 47400 471232 47452 471238
rect 47400 471174 47452 471180
rect 47412 379409 47440 471174
rect 47492 471164 47544 471170
rect 47492 471106 47544 471112
rect 47398 379400 47454 379409
rect 47398 379335 47454 379344
rect 47412 373994 47440 379335
rect 47504 378842 47532 471106
rect 47596 380186 47624 479538
rect 47584 380180 47636 380186
rect 47584 380122 47636 380128
rect 47688 379302 47716 479742
rect 47768 479732 47820 479738
rect 47768 479674 47820 479680
rect 47780 379438 47808 479674
rect 47768 379432 47820 379438
rect 47768 379374 47820 379380
rect 47676 379296 47728 379302
rect 47676 379238 47728 379244
rect 47766 378992 47822 379001
rect 47766 378927 47822 378936
rect 47780 378842 47808 378927
rect 47504 378814 47808 378842
rect 47676 378616 47728 378622
rect 47676 378558 47728 378564
rect 47688 378214 47716 378558
rect 47676 378208 47728 378214
rect 47676 378150 47728 378156
rect 47412 373966 47624 373994
rect 47596 271425 47624 373966
rect 47688 271833 47716 378150
rect 47674 271824 47730 271833
rect 47674 271759 47730 271768
rect 47780 271697 47808 378814
rect 47872 272474 47900 482734
rect 47950 482488 48006 482497
rect 47950 482423 48006 482432
rect 47860 272468 47912 272474
rect 47860 272410 47912 272416
rect 47872 271946 47900 272410
rect 47964 272066 47992 482423
rect 48056 272678 48084 482870
rect 49240 482860 49292 482866
rect 49240 482802 49292 482808
rect 49148 482452 49200 482458
rect 49148 482394 49200 482400
rect 48136 482384 48188 482390
rect 48136 482326 48188 482332
rect 48044 272672 48096 272678
rect 48044 272614 48096 272620
rect 47952 272060 48004 272066
rect 47952 272002 48004 272008
rect 47872 271918 47992 271946
rect 47766 271688 47822 271697
rect 47766 271623 47822 271632
rect 47582 271416 47638 271425
rect 47582 271351 47638 271360
rect 47780 267734 47808 271623
rect 47780 267706 47900 267734
rect 46848 251184 46900 251190
rect 46848 251126 46900 251132
rect 46664 148844 46716 148850
rect 46664 148786 46716 148792
rect 47872 145858 47900 267706
rect 47860 145852 47912 145858
rect 47860 145794 47912 145800
rect 47964 145450 47992 271918
rect 48042 271824 48098 271833
rect 48042 271759 48098 271768
rect 48056 271017 48084 271759
rect 48148 271153 48176 482326
rect 48228 480072 48280 480078
rect 48228 480014 48280 480020
rect 48134 271144 48190 271153
rect 48134 271079 48190 271088
rect 48042 271008 48098 271017
rect 48042 270943 48098 270952
rect 48056 148782 48084 270943
rect 48240 268870 48268 480014
rect 49056 477080 49108 477086
rect 49056 477022 49108 477028
rect 48964 477012 49016 477018
rect 48964 476954 49016 476960
rect 48780 468988 48832 468994
rect 48780 468930 48832 468936
rect 48228 268864 48280 268870
rect 48228 268806 48280 268812
rect 48044 148776 48096 148782
rect 48044 148718 48096 148724
rect 47952 145444 48004 145450
rect 47952 145386 48004 145392
rect 46572 145376 46624 145382
rect 46572 145318 46624 145324
rect 48792 58818 48820 468930
rect 48872 466540 48924 466546
rect 48872 466482 48924 466488
rect 48884 418130 48912 466482
rect 48872 418124 48924 418130
rect 48872 418066 48924 418072
rect 48872 409896 48924 409902
rect 48872 409838 48924 409844
rect 48884 377262 48912 409838
rect 48976 380390 49004 476954
rect 48964 380384 49016 380390
rect 48964 380326 49016 380332
rect 49068 378690 49096 477022
rect 49056 378684 49108 378690
rect 49056 378626 49108 378632
rect 48872 377256 48924 377262
rect 48872 377198 48924 377204
rect 49160 273018 49188 482394
rect 49148 273012 49200 273018
rect 49148 272954 49200 272960
rect 49252 272610 49280 482802
rect 50342 479768 50398 479777
rect 50342 479703 50398 479712
rect 50068 477148 50120 477154
rect 50068 477090 50120 477096
rect 49424 471708 49476 471714
rect 49424 471650 49476 471656
rect 49332 468512 49384 468518
rect 49332 468454 49384 468460
rect 49240 272604 49292 272610
rect 49240 272546 49292 272552
rect 49146 271416 49202 271425
rect 49146 271351 49202 271360
rect 49056 268592 49108 268598
rect 49056 268534 49108 268540
rect 49068 268394 49096 268534
rect 49056 268388 49108 268394
rect 49056 268330 49108 268336
rect 49068 164218 49096 268330
rect 49056 164212 49108 164218
rect 49056 164154 49108 164160
rect 49160 148646 49188 271351
rect 49240 268660 49292 268666
rect 49240 268602 49292 268608
rect 49252 268462 49280 268602
rect 49240 268456 49292 268462
rect 49240 268398 49292 268404
rect 49148 148640 49200 148646
rect 49148 148582 49200 148588
rect 49252 144634 49280 268398
rect 49344 165481 49372 468454
rect 49436 167006 49464 471650
rect 49516 469192 49568 469198
rect 49516 469134 49568 469140
rect 49528 467945 49556 469134
rect 49514 467936 49570 467945
rect 49514 467871 49570 467880
rect 49516 465724 49568 465730
rect 49516 465666 49568 465672
rect 49424 167000 49476 167006
rect 49424 166942 49476 166948
rect 49330 165472 49386 165481
rect 49330 165407 49386 165416
rect 49240 144628 49292 144634
rect 49240 144570 49292 144576
rect 49528 59430 49556 465666
rect 49608 411324 49660 411330
rect 49608 411266 49660 411272
rect 49620 380905 49648 411266
rect 49606 380896 49662 380905
rect 49606 380831 49662 380840
rect 50080 378758 50108 477090
rect 50252 471368 50304 471374
rect 50252 471310 50304 471316
rect 50160 412752 50212 412758
rect 50160 412694 50212 412700
rect 50172 380730 50200 412694
rect 50160 380724 50212 380730
rect 50160 380666 50212 380672
rect 50068 378752 50120 378758
rect 50068 378694 50120 378700
rect 50264 271114 50292 471310
rect 50356 272814 50384 479703
rect 50344 272808 50396 272814
rect 50344 272750 50396 272756
rect 50448 272746 50476 482938
rect 50528 482656 50580 482662
rect 50528 482598 50580 482604
rect 50436 272740 50488 272746
rect 50436 272682 50488 272688
rect 50252 271108 50304 271114
rect 50252 271050 50304 271056
rect 50540 270434 50568 482598
rect 51000 480254 51028 485250
rect 51816 485240 51868 485246
rect 51816 485182 51868 485188
rect 50908 480226 51028 480254
rect 50620 471776 50672 471782
rect 50620 471718 50672 471724
rect 50528 270428 50580 270434
rect 50528 270370 50580 270376
rect 50436 268388 50488 268394
rect 50436 268330 50488 268336
rect 50448 144770 50476 268330
rect 50436 144764 50488 144770
rect 50436 144706 50488 144712
rect 50540 144702 50568 270370
rect 50632 166258 50660 471718
rect 50804 469940 50856 469946
rect 50804 469882 50856 469888
rect 50712 469124 50764 469130
rect 50712 469066 50764 469072
rect 50724 467945 50752 469066
rect 50710 467936 50766 467945
rect 50710 467871 50766 467880
rect 50816 465882 50844 469882
rect 50724 465854 50844 465882
rect 50620 166252 50672 166258
rect 50620 166194 50672 166200
rect 50724 164898 50752 465854
rect 50804 465792 50856 465798
rect 50804 465734 50856 465740
rect 50816 166938 50844 465734
rect 50804 166932 50856 166938
rect 50804 166874 50856 166880
rect 50908 165345 50936 480226
rect 51724 479460 51776 479466
rect 51724 479402 51776 479408
rect 51632 474156 51684 474162
rect 51632 474098 51684 474104
rect 50988 471912 51040 471918
rect 50988 471854 51040 471860
rect 51000 465798 51028 471854
rect 51540 471844 51592 471850
rect 51540 471786 51592 471792
rect 51448 466064 51500 466070
rect 51448 466006 51500 466012
rect 50988 465792 51040 465798
rect 50988 465734 51040 465740
rect 50986 379536 51042 379545
rect 50986 379471 51042 379480
rect 50894 165336 50950 165345
rect 50894 165271 50950 165280
rect 50712 164892 50764 164898
rect 50712 164834 50764 164840
rect 50896 164212 50948 164218
rect 50896 164154 50948 164160
rect 50804 164144 50856 164150
rect 50804 164086 50856 164092
rect 50816 163538 50844 164086
rect 50908 163674 50936 164154
rect 50896 163668 50948 163674
rect 50896 163610 50948 163616
rect 50804 163532 50856 163538
rect 50804 163474 50856 163480
rect 50528 144696 50580 144702
rect 50528 144638 50580 144644
rect 49516 59424 49568 59430
rect 49516 59366 49568 59372
rect 48780 58812 48832 58818
rect 48780 58754 48832 58760
rect 50816 56506 50844 163474
rect 50804 56500 50856 56506
rect 50804 56442 50856 56448
rect 50908 54942 50936 163610
rect 51000 58682 51028 379471
rect 50988 58676 51040 58682
rect 50988 58618 51040 58624
rect 51460 57458 51488 466006
rect 51552 465798 51580 471786
rect 51540 465792 51592 465798
rect 51540 465734 51592 465740
rect 51540 414044 51592 414050
rect 51540 413986 51592 413992
rect 51552 380089 51580 413986
rect 51538 380080 51594 380089
rect 51538 380015 51594 380024
rect 51538 379128 51594 379137
rect 51538 379063 51594 379072
rect 51552 282198 51580 379063
rect 51540 282192 51592 282198
rect 51540 282134 51592 282140
rect 51540 273080 51592 273086
rect 51540 273022 51592 273028
rect 51552 163878 51580 273022
rect 51644 271250 51672 474098
rect 51632 271244 51684 271250
rect 51632 271186 51684 271192
rect 51736 270162 51764 479402
rect 51828 271182 51856 485182
rect 52184 485036 52236 485042
rect 52184 484978 52236 484984
rect 51908 482248 51960 482254
rect 51908 482190 51960 482196
rect 51920 272542 51948 482190
rect 52092 471096 52144 471102
rect 52092 471038 52144 471044
rect 52000 466336 52052 466342
rect 52000 466278 52052 466284
rect 52012 465905 52040 466278
rect 51998 465896 52054 465905
rect 51998 465831 52054 465840
rect 52000 465792 52052 465798
rect 52000 465734 52052 465740
rect 51908 272536 51960 272542
rect 51908 272478 51960 272484
rect 51816 271176 51868 271182
rect 51816 271118 51868 271124
rect 51814 270328 51870 270337
rect 51814 270263 51870 270272
rect 51724 270156 51776 270162
rect 51724 270098 51776 270104
rect 51724 269816 51776 269822
rect 51724 269758 51776 269764
rect 51736 269074 51764 269758
rect 51724 269068 51776 269074
rect 51724 269010 51776 269016
rect 51540 163872 51592 163878
rect 51540 163814 51592 163820
rect 51736 144906 51764 269010
rect 51724 144900 51776 144906
rect 51724 144842 51776 144848
rect 51828 144838 51856 270263
rect 52012 166870 52040 465734
rect 52000 166864 52052 166870
rect 52000 166806 52052 166812
rect 52104 164966 52132 471038
rect 52092 164960 52144 164966
rect 52092 164902 52144 164908
rect 52196 164830 52224 484978
rect 53562 471608 53618 471617
rect 53562 471543 53618 471552
rect 53288 471504 53340 471510
rect 53288 471446 53340 471452
rect 53196 471436 53248 471442
rect 53196 471378 53248 471384
rect 53104 467628 53156 467634
rect 53104 467570 53156 467576
rect 52368 467560 52420 467566
rect 52368 467502 52420 467508
rect 52276 466404 52328 466410
rect 52276 466346 52328 466352
rect 52288 465225 52316 466346
rect 52274 465216 52330 465225
rect 52274 465151 52330 465160
rect 52380 451274 52408 467502
rect 52920 464500 52972 464506
rect 52920 464442 52972 464448
rect 52288 451246 52408 451274
rect 52288 411126 52316 451246
rect 52276 411120 52328 411126
rect 52276 411062 52328 411068
rect 52368 408536 52420 408542
rect 52368 408478 52420 408484
rect 52380 380633 52408 408478
rect 52932 380798 52960 464442
rect 53012 411120 53064 411126
rect 53012 411062 53064 411068
rect 52920 380792 52972 380798
rect 52920 380734 52972 380740
rect 52366 380624 52422 380633
rect 52366 380559 52422 380568
rect 52274 379536 52330 379545
rect 52274 379471 52330 379480
rect 52184 164824 52236 164830
rect 52184 164766 52236 164772
rect 52184 148640 52236 148646
rect 52184 148582 52236 148588
rect 52092 146260 52144 146266
rect 52092 146202 52144 146208
rect 52104 145518 52132 146202
rect 52092 145512 52144 145518
rect 52092 145454 52144 145460
rect 51816 144832 51868 144838
rect 51816 144774 51868 144780
rect 51448 57452 51500 57458
rect 51448 57394 51500 57400
rect 52104 57254 52132 145454
rect 52092 57248 52144 57254
rect 52092 57190 52144 57196
rect 50896 54936 50948 54942
rect 50896 54878 50948 54884
rect 52196 54602 52224 148582
rect 52288 57730 52316 379471
rect 53024 287054 53052 411062
rect 52932 287026 53052 287054
rect 52366 282296 52422 282305
rect 52366 282231 52422 282240
rect 52380 57866 52408 282231
rect 52828 272060 52880 272066
rect 52828 272002 52880 272008
rect 52840 267734 52868 272002
rect 52932 271386 52960 287026
rect 53116 277394 53144 467570
rect 53024 277366 53144 277394
rect 52920 271380 52972 271386
rect 52920 271322 52972 271328
rect 53024 271318 53052 277366
rect 53208 274530 53236 471378
rect 53116 274502 53236 274530
rect 53116 271454 53144 274502
rect 53300 274394 53328 471446
rect 53380 468716 53432 468722
rect 53380 468658 53432 468664
rect 53208 274366 53328 274394
rect 53208 271522 53236 274366
rect 53286 271824 53342 271833
rect 53286 271759 53342 271768
rect 53196 271516 53248 271522
rect 53196 271458 53248 271464
rect 53104 271448 53156 271454
rect 53104 271390 53156 271396
rect 53012 271312 53064 271318
rect 53012 271254 53064 271260
rect 53196 270020 53248 270026
rect 53196 269962 53248 269968
rect 52840 267706 52960 267734
rect 52460 251864 52512 251870
rect 52460 251806 52512 251812
rect 52472 251190 52500 251806
rect 52460 251184 52512 251190
rect 52460 251126 52512 251132
rect 52932 163810 52960 267706
rect 53012 251184 53064 251190
rect 53012 251126 53064 251132
rect 53024 165714 53052 251126
rect 53012 165708 53064 165714
rect 53012 165650 53064 165656
rect 52920 163804 52972 163810
rect 52920 163746 52972 163752
rect 52368 57860 52420 57866
rect 52368 57802 52420 57808
rect 52276 57724 52328 57730
rect 52276 57666 52328 57672
rect 53024 55010 53052 165650
rect 53104 145852 53156 145858
rect 53104 145794 53156 145800
rect 53116 55214 53144 145794
rect 53208 144566 53236 269962
rect 53196 144560 53248 144566
rect 53196 144502 53248 144508
rect 53300 58750 53328 271759
rect 53392 165102 53420 468658
rect 53472 468580 53524 468586
rect 53472 468522 53524 468528
rect 53484 165306 53512 468522
rect 53576 166802 53604 471543
rect 53654 471336 53710 471345
rect 53654 471271 53710 471280
rect 53564 166796 53616 166802
rect 53564 166738 53616 166744
rect 53472 165300 53524 165306
rect 53472 165242 53524 165248
rect 53380 165096 53432 165102
rect 53380 165038 53432 165044
rect 53668 163946 53696 471271
rect 53760 389162 53788 517482
rect 303356 510513 303384 574058
rect 304276 558346 304304 596158
rect 304264 558340 304316 558346
rect 304264 558282 304316 558288
rect 304264 551540 304316 551546
rect 304264 551482 304316 551488
rect 304276 527105 304304 551482
rect 305656 527950 305684 700402
rect 364352 645182 364380 702406
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 434720 700460 434772 700466
rect 434720 700402 434772 700408
rect 405924 646536 405976 646542
rect 405924 646478 405976 646484
rect 364340 645176 364392 645182
rect 364340 645118 364392 645124
rect 322572 643136 322624 643142
rect 322572 643078 322624 643084
rect 322480 642728 322532 642734
rect 322480 642670 322532 642676
rect 316776 642592 316828 642598
rect 316776 642534 316828 642540
rect 309784 642524 309836 642530
rect 309784 642466 309836 642472
rect 307024 642184 307076 642190
rect 307024 642126 307076 642132
rect 305736 581052 305788 581058
rect 305736 580994 305788 581000
rect 305748 559706 305776 580994
rect 307036 563922 307064 642126
rect 307116 590708 307168 590714
rect 307116 590650 307168 590656
rect 307128 575482 307156 590650
rect 307116 575476 307168 575482
rect 307116 575418 307168 575424
rect 309796 569294 309824 642466
rect 311164 641980 311216 641986
rect 311164 641922 311216 641928
rect 309876 614168 309928 614174
rect 309876 614110 309928 614116
rect 309784 569288 309836 569294
rect 309784 569230 309836 569236
rect 307024 563916 307076 563922
rect 307024 563858 307076 563864
rect 305736 559700 305788 559706
rect 305736 559642 305788 559648
rect 309888 552906 309916 614110
rect 309968 586560 310020 586566
rect 309968 586502 310020 586508
rect 309980 572082 310008 586502
rect 309968 572076 310020 572082
rect 309968 572018 310020 572024
rect 309876 552900 309928 552906
rect 309876 552842 309928 552848
rect 311176 552838 311204 641922
rect 314108 640824 314160 640830
rect 314108 640766 314160 640772
rect 314016 640620 314068 640626
rect 314016 640562 314068 640568
rect 312544 633480 312596 633486
rect 312544 633422 312596 633428
rect 311256 619676 311308 619682
rect 311256 619618 311308 619624
rect 311164 552832 311216 552838
rect 311164 552774 311216 552780
rect 311268 552770 311296 619618
rect 311348 605872 311400 605878
rect 311348 605814 311400 605820
rect 311360 566710 311388 605814
rect 311348 566704 311400 566710
rect 311348 566646 311400 566652
rect 311256 552764 311308 552770
rect 311256 552706 311308 552712
rect 312556 551342 312584 633422
rect 313924 629332 313976 629338
rect 313924 629274 313976 629280
rect 313936 555558 313964 629274
rect 314028 575346 314056 640562
rect 314016 575340 314068 575346
rect 314016 575282 314068 575288
rect 314120 574734 314148 640766
rect 316684 640756 316736 640762
rect 316684 640698 316736 640704
rect 314200 610020 314252 610026
rect 314200 609962 314252 609968
rect 314108 574728 314160 574734
rect 314108 574670 314160 574676
rect 314212 556918 314240 609962
rect 314200 556912 314252 556918
rect 314200 556854 314252 556860
rect 313924 555552 313976 555558
rect 313924 555494 313976 555500
rect 312544 551336 312596 551342
rect 312544 551278 312596 551284
rect 316696 549982 316724 640698
rect 316788 565282 316816 642534
rect 318156 642388 318208 642394
rect 318156 642330 318208 642336
rect 316868 640348 316920 640354
rect 316868 640290 316920 640296
rect 316880 575142 316908 640290
rect 316960 639192 317012 639198
rect 316960 639134 317012 639140
rect 316972 575210 317000 639134
rect 317052 639056 317104 639062
rect 317052 638998 317104 639004
rect 316960 575204 317012 575210
rect 316960 575146 317012 575152
rect 316868 575136 316920 575142
rect 316868 575078 316920 575084
rect 317064 575074 317092 638998
rect 318064 623824 318116 623830
rect 318064 623766 318116 623772
rect 317052 575068 317104 575074
rect 317052 575010 317104 575016
rect 316776 565276 316828 565282
rect 316776 565218 316828 565224
rect 316684 549976 316736 549982
rect 316684 549918 316736 549924
rect 305736 549636 305788 549642
rect 305736 549578 305788 549584
rect 305748 529582 305776 549578
rect 307024 548684 307076 548690
rect 307024 548626 307076 548632
rect 305736 529576 305788 529582
rect 305736 529518 305788 529524
rect 305644 527944 305696 527950
rect 305644 527886 305696 527892
rect 307036 527134 307064 548626
rect 311164 539640 311216 539646
rect 311164 539582 311216 539588
rect 307024 527128 307076 527134
rect 304262 527096 304318 527105
rect 307024 527070 307076 527076
rect 304262 527031 304318 527040
rect 311176 515438 311204 539582
rect 311164 515432 311216 515438
rect 311164 515374 311216 515380
rect 303342 510504 303398 510513
rect 303342 510439 303398 510448
rect 302238 495544 302294 495553
rect 302238 495479 302240 495488
rect 302292 495479 302294 495488
rect 302240 495450 302292 495456
rect 59372 488022 60214 488050
rect 60598 488022 60688 488050
rect 56508 485648 56560 485654
rect 56508 485590 56560 485596
rect 55128 485444 55180 485450
rect 55128 485386 55180 485392
rect 54852 482180 54904 482186
rect 54852 482122 54904 482128
rect 54760 479324 54812 479330
rect 54760 479266 54812 479272
rect 54484 477216 54536 477222
rect 54484 477158 54536 477164
rect 54392 466200 54444 466206
rect 54392 466142 54444 466148
rect 54300 466132 54352 466138
rect 54300 466074 54352 466080
rect 53748 389156 53800 389162
rect 53748 389098 53800 389104
rect 53746 388512 53802 388521
rect 53746 388447 53802 388456
rect 53656 163940 53708 163946
rect 53656 163882 53708 163888
rect 53472 148504 53524 148510
rect 53472 148446 53524 148452
rect 53380 148368 53432 148374
rect 53380 148310 53432 148316
rect 53288 58744 53340 58750
rect 53288 58686 53340 58692
rect 53392 56574 53420 148310
rect 53380 56568 53432 56574
rect 53380 56510 53432 56516
rect 53484 56438 53512 148446
rect 53564 148436 53616 148442
rect 53564 148378 53616 148384
rect 53472 56432 53524 56438
rect 53472 56374 53524 56380
rect 53104 55208 53156 55214
rect 53104 55150 53156 55156
rect 53576 55078 53604 148378
rect 53656 146056 53708 146062
rect 53656 145998 53708 146004
rect 53564 55072 53616 55078
rect 53564 55014 53616 55020
rect 53012 55004 53064 55010
rect 53012 54946 53064 54952
rect 53668 54738 53696 145998
rect 53760 57798 53788 388447
rect 54312 377874 54340 466074
rect 54404 377942 54432 466142
rect 54496 380526 54524 477158
rect 54668 471640 54720 471646
rect 54668 471582 54720 471588
rect 54576 464568 54628 464574
rect 54576 464510 54628 464516
rect 54484 380520 54536 380526
rect 54484 380462 54536 380468
rect 54392 377936 54444 377942
rect 54392 377878 54444 377884
rect 54300 377868 54352 377874
rect 54300 377810 54352 377816
rect 54484 358080 54536 358086
rect 54484 358022 54536 358028
rect 54300 273012 54352 273018
rect 54300 272954 54352 272960
rect 53840 272808 53892 272814
rect 53838 272776 53840 272785
rect 53892 272776 53894 272785
rect 53838 272711 53894 272720
rect 54206 272776 54262 272785
rect 54206 272711 54262 272720
rect 54116 272264 54168 272270
rect 54116 272206 54168 272212
rect 54024 165640 54076 165646
rect 54024 165582 54076 165588
rect 53840 145716 53892 145722
rect 53840 145658 53892 145664
rect 53852 144906 53880 145658
rect 53932 145580 53984 145586
rect 53932 145522 53984 145528
rect 53840 144900 53892 144906
rect 53840 144842 53892 144848
rect 53944 144770 53972 145522
rect 53932 144764 53984 144770
rect 53932 144706 53984 144712
rect 53748 57792 53800 57798
rect 53748 57734 53800 57740
rect 54036 55146 54064 165582
rect 54128 146062 54156 272206
rect 54220 146305 54248 272711
rect 54206 146296 54262 146305
rect 54206 146231 54262 146240
rect 54116 146056 54168 146062
rect 54116 145998 54168 146004
rect 54312 145994 54340 272954
rect 54496 271726 54524 358022
rect 54484 271720 54536 271726
rect 54484 271662 54536 271668
rect 54588 271658 54616 464510
rect 54576 271652 54628 271658
rect 54576 271594 54628 271600
rect 54680 271590 54708 471582
rect 54772 272270 54800 479266
rect 54760 272264 54812 272270
rect 54760 272206 54812 272212
rect 54668 271584 54720 271590
rect 54668 271526 54720 271532
rect 54864 271046 54892 482122
rect 55034 471200 55090 471209
rect 55034 471135 55090 471144
rect 54944 468784 54996 468790
rect 54944 468726 54996 468732
rect 54852 271040 54904 271046
rect 54852 270982 54904 270988
rect 54576 270156 54628 270162
rect 54576 270098 54628 270104
rect 54392 252000 54444 252006
rect 54392 251942 54444 251948
rect 54404 165646 54432 251942
rect 54484 251932 54536 251938
rect 54484 251874 54536 251880
rect 54392 165640 54444 165646
rect 54392 165582 54444 165588
rect 54496 148578 54524 251874
rect 54484 148572 54536 148578
rect 54484 148514 54536 148520
rect 54300 145988 54352 145994
rect 54300 145930 54352 145936
rect 54392 145444 54444 145450
rect 54392 145386 54444 145392
rect 54404 59702 54432 145386
rect 54588 144906 54616 270098
rect 54956 165170 54984 468726
rect 55048 165510 55076 471135
rect 55036 165504 55088 165510
rect 55036 165446 55088 165452
rect 55140 165374 55168 485386
rect 56416 485376 56468 485382
rect 56416 485318 56468 485324
rect 55956 477284 56008 477290
rect 55956 477226 56008 477232
rect 55864 464636 55916 464642
rect 55864 464578 55916 464584
rect 55772 417172 55824 417178
rect 55772 417114 55824 417120
rect 55680 413976 55732 413982
rect 55680 413918 55732 413924
rect 55692 378962 55720 413918
rect 55680 378956 55732 378962
rect 55680 378898 55732 378904
rect 55784 378826 55812 417114
rect 55876 381750 55904 464578
rect 55864 381744 55916 381750
rect 55864 381686 55916 381692
rect 55864 380792 55916 380798
rect 55864 380734 55916 380740
rect 55772 378820 55824 378826
rect 55772 378762 55824 378768
rect 55876 282674 55904 380734
rect 55968 380458 55996 477226
rect 56322 471472 56378 471481
rect 56322 471407 56378 471416
rect 56140 468920 56192 468926
rect 56140 468862 56192 468868
rect 56048 465860 56100 465866
rect 56048 465802 56100 465808
rect 55956 380452 56008 380458
rect 55956 380394 56008 380400
rect 55864 282668 55916 282674
rect 55864 282610 55916 282616
rect 55956 269952 56008 269958
rect 55956 269894 56008 269900
rect 55968 268870 55996 269894
rect 55956 268864 56008 268870
rect 55956 268806 56008 268812
rect 55968 258074 55996 268806
rect 55876 258046 55996 258074
rect 55128 165368 55180 165374
rect 55128 165310 55180 165316
rect 54944 165164 54996 165170
rect 54944 165106 54996 165112
rect 55876 151814 55904 258046
rect 56060 165073 56088 465802
rect 56046 165064 56102 165073
rect 56152 165034 56180 468862
rect 56232 468852 56284 468858
rect 56232 468794 56284 468800
rect 56244 165238 56272 468794
rect 56336 165442 56364 471407
rect 56428 166734 56456 485318
rect 56416 166728 56468 166734
rect 56416 166670 56468 166676
rect 56520 165578 56548 485590
rect 59084 485580 59136 485586
rect 59084 485522 59136 485528
rect 58716 482112 58768 482118
rect 58716 482054 58768 482060
rect 57888 481024 57940 481030
rect 57888 480966 57940 480972
rect 57244 480208 57296 480214
rect 57244 480150 57296 480156
rect 57060 464432 57112 464438
rect 57060 464374 57112 464380
rect 57072 422294 57100 464374
rect 57152 464364 57204 464370
rect 57152 464306 57204 464312
rect 56980 422266 57100 422294
rect 56876 416220 56928 416226
rect 56876 416162 56928 416168
rect 56690 410408 56746 410417
rect 56690 410343 56746 410352
rect 56704 409902 56732 410343
rect 56692 409896 56744 409902
rect 56692 409838 56744 409844
rect 56888 380254 56916 416162
rect 56980 413982 57008 422266
rect 57060 418124 57112 418130
rect 57060 418066 57112 418072
rect 57072 417897 57100 418066
rect 57058 417888 57114 417897
rect 57058 417823 57114 417832
rect 57058 414216 57114 414225
rect 57058 414151 57114 414160
rect 57072 414050 57100 414151
rect 57060 414044 57112 414050
rect 57060 413986 57112 413992
rect 56968 413976 57020 413982
rect 56968 413918 57020 413924
rect 57164 393314 57192 464306
rect 57256 417178 57284 480150
rect 57428 477352 57480 477358
rect 57428 477294 57480 477300
rect 57336 471572 57388 471578
rect 57336 471514 57388 471520
rect 57244 417172 57296 417178
rect 57244 417114 57296 417120
rect 57242 416936 57298 416945
rect 57242 416871 57298 416880
rect 57256 416838 57284 416871
rect 57244 416832 57296 416838
rect 57244 416774 57296 416780
rect 57242 413264 57298 413273
rect 57242 413199 57298 413208
rect 57256 412758 57284 413199
rect 57244 412752 57296 412758
rect 57244 412694 57296 412700
rect 57242 411496 57298 411505
rect 57242 411431 57298 411440
rect 57256 411330 57284 411431
rect 57244 411324 57296 411330
rect 57244 411266 57296 411272
rect 57242 408640 57298 408649
rect 57242 408575 57298 408584
rect 57256 408542 57284 408575
rect 57244 408536 57296 408542
rect 57244 408478 57296 408484
rect 56980 393286 57192 393314
rect 56980 383654 57008 393286
rect 57244 391944 57296 391950
rect 57244 391886 57296 391892
rect 57256 391649 57284 391886
rect 57242 391640 57298 391649
rect 57242 391575 57298 391584
rect 57060 389564 57112 389570
rect 57060 389506 57112 389512
rect 57072 388414 57100 389506
rect 57244 389156 57296 389162
rect 57244 389098 57296 389104
rect 57152 389088 57204 389094
rect 57150 389056 57152 389065
rect 57204 389056 57206 389065
rect 57150 388991 57206 389000
rect 57060 388408 57112 388414
rect 57060 388350 57112 388356
rect 56980 383626 57100 383654
rect 56876 380248 56928 380254
rect 56876 380190 56928 380196
rect 57072 378894 57100 383626
rect 57060 378888 57112 378894
rect 57060 378830 57112 378836
rect 56968 378820 57020 378826
rect 56968 378762 57020 378768
rect 56874 309904 56930 309913
rect 56874 309839 56930 309848
rect 56782 301608 56838 301617
rect 56782 301543 56838 301552
rect 56796 300830 56824 301543
rect 56784 300824 56836 300830
rect 56784 300766 56836 300772
rect 56888 203425 56916 309839
rect 56980 300830 57008 378762
rect 57152 358692 57204 358698
rect 57152 358634 57204 358640
rect 56968 300824 57020 300830
rect 56968 300766 57020 300772
rect 57060 300756 57112 300762
rect 57060 300698 57112 300704
rect 56968 251388 57020 251394
rect 56968 251330 57020 251336
rect 56874 203416 56930 203425
rect 56874 203351 56930 203360
rect 56508 165572 56560 165578
rect 56508 165514 56560 165520
rect 56324 165436 56376 165442
rect 56324 165378 56376 165384
rect 56232 165232 56284 165238
rect 56232 165174 56284 165180
rect 56046 164999 56102 165008
rect 56140 165028 56192 165034
rect 56140 164970 56192 164976
rect 56980 164014 57008 251330
rect 57072 195265 57100 300698
rect 57164 271794 57192 358634
rect 57256 282577 57284 389098
rect 57348 381002 57376 471514
rect 57440 389570 57468 477294
rect 57612 475448 57664 475454
rect 57612 475390 57664 475396
rect 57520 469872 57572 469878
rect 57520 469814 57572 469820
rect 57428 389564 57480 389570
rect 57428 389506 57480 389512
rect 57532 389450 57560 469814
rect 57440 389422 57560 389450
rect 57440 388498 57468 389422
rect 57518 389328 57574 389337
rect 57518 389263 57574 389272
rect 57532 389162 57560 389263
rect 57520 389156 57572 389162
rect 57520 389098 57572 389104
rect 57440 388470 57560 388498
rect 57428 388408 57480 388414
rect 57428 388350 57480 388356
rect 57336 380996 57388 381002
rect 57336 380938 57388 380944
rect 57440 380322 57468 388350
rect 57428 380316 57480 380322
rect 57428 380258 57480 380264
rect 57426 309088 57482 309097
rect 57426 309023 57482 309032
rect 57440 307873 57468 309023
rect 57426 307864 57482 307873
rect 57426 307799 57482 307808
rect 57336 303612 57388 303618
rect 57336 303554 57388 303560
rect 57242 282568 57298 282577
rect 57242 282503 57298 282512
rect 57152 271788 57204 271794
rect 57152 271730 57204 271736
rect 57152 269884 57204 269890
rect 57152 269826 57204 269832
rect 57164 268938 57192 269826
rect 57152 268932 57204 268938
rect 57152 268874 57204 268880
rect 57058 195256 57114 195265
rect 57058 195191 57114 195200
rect 57060 175228 57112 175234
rect 57060 175170 57112 175176
rect 57072 175137 57100 175170
rect 57058 175128 57114 175137
rect 57058 175063 57114 175072
rect 56968 164008 57020 164014
rect 56968 163950 57020 163956
rect 56876 163872 56928 163878
rect 56876 163814 56928 163820
rect 56508 163804 56560 163810
rect 56508 163746 56560 163752
rect 55876 151786 55996 151814
rect 55036 148776 55088 148782
rect 55036 148718 55088 148724
rect 54758 146296 54814 146305
rect 54758 146231 54814 146240
rect 54484 144900 54536 144906
rect 54484 144842 54536 144848
rect 54576 144900 54628 144906
rect 54576 144842 54628 144848
rect 54392 59696 54444 59702
rect 54392 59638 54444 59644
rect 54496 56166 54524 144842
rect 54668 144764 54720 144770
rect 54668 144706 54720 144712
rect 54680 59022 54708 144706
rect 54772 59498 54800 146231
rect 54852 145988 54904 145994
rect 54852 145930 54904 145936
rect 54864 59634 54892 145930
rect 54944 145376 54996 145382
rect 54944 145318 54996 145324
rect 54852 59628 54904 59634
rect 54852 59570 54904 59576
rect 54760 59492 54812 59498
rect 54760 59434 54812 59440
rect 54668 59016 54720 59022
rect 54668 58958 54720 58964
rect 54956 57118 54984 145318
rect 54944 57112 54996 57118
rect 54944 57054 54996 57060
rect 54484 56160 54536 56166
rect 54484 56102 54536 56108
rect 55048 56030 55076 148718
rect 55968 146130 55996 151786
rect 56232 148572 56284 148578
rect 56232 148514 56284 148520
rect 56138 146160 56194 146169
rect 55956 146124 56008 146130
rect 56138 146095 56194 146104
rect 55956 146066 56008 146072
rect 55864 144696 55916 144702
rect 55864 144638 55916 144644
rect 55876 59362 55904 144638
rect 55968 144430 55996 146066
rect 55956 144424 56008 144430
rect 55956 144366 56008 144372
rect 55864 59356 55916 59362
rect 55864 59298 55916 59304
rect 56152 57526 56180 146095
rect 56244 58954 56272 148514
rect 56324 147688 56376 147694
rect 56324 147630 56376 147636
rect 56336 144514 56364 147630
rect 56416 145784 56468 145790
rect 56416 145726 56468 145732
rect 56428 144702 56456 145726
rect 56416 144696 56468 144702
rect 56416 144638 56468 144644
rect 56336 144486 56456 144514
rect 56324 144424 56376 144430
rect 56324 144366 56376 144372
rect 56232 58948 56284 58954
rect 56232 58890 56284 58896
rect 56140 57520 56192 57526
rect 56140 57462 56192 57468
rect 56336 56234 56364 144366
rect 56428 57594 56456 144486
rect 56520 59090 56548 163746
rect 56888 59158 56916 163814
rect 57164 162858 57192 268874
rect 57242 204232 57298 204241
rect 57242 204167 57298 204176
rect 57152 162852 57204 162858
rect 57152 162794 57204 162800
rect 57060 146260 57112 146266
rect 57060 146202 57112 146208
rect 56876 59152 56928 59158
rect 56876 59094 56928 59100
rect 56508 59084 56560 59090
rect 56508 59026 56560 59032
rect 56416 57588 56468 57594
rect 56416 57530 56468 57536
rect 56324 56228 56376 56234
rect 56324 56170 56376 56176
rect 55036 56024 55088 56030
rect 55036 55966 55088 55972
rect 54024 55140 54076 55146
rect 54024 55082 54076 55088
rect 57072 54806 57100 146202
rect 57256 97481 57284 204167
rect 57348 197033 57376 303554
rect 57440 209774 57468 307799
rect 57532 305017 57560 388470
rect 57624 311137 57652 475390
rect 57796 474088 57848 474094
rect 57796 474030 57848 474036
rect 57704 471300 57756 471306
rect 57704 471242 57756 471248
rect 57610 311128 57666 311137
rect 57610 311063 57666 311072
rect 57518 305008 57574 305017
rect 57518 304943 57574 304952
rect 57518 303648 57574 303657
rect 57518 303583 57520 303592
rect 57572 303583 57574 303592
rect 57520 303554 57572 303560
rect 57440 209746 57560 209774
rect 57532 203538 57560 209746
rect 57624 204241 57652 311063
rect 57716 306785 57744 471242
rect 57808 309097 57836 474030
rect 57900 309913 57928 480966
rect 58532 479392 58584 479398
rect 58532 479334 58584 479340
rect 58440 476740 58492 476746
rect 58440 476682 58492 476688
rect 58452 380934 58480 476682
rect 58544 381886 58572 479334
rect 58624 472660 58676 472666
rect 58624 472602 58676 472608
rect 58532 381880 58584 381886
rect 58532 381822 58584 381828
rect 58440 380928 58492 380934
rect 58440 380870 58492 380876
rect 58532 357400 58584 357406
rect 58532 357342 58584 357348
rect 57886 309904 57942 309913
rect 57886 309839 57942 309848
rect 57794 309088 57850 309097
rect 57794 309023 57850 309032
rect 57702 306776 57758 306785
rect 57702 306711 57758 306720
rect 57610 204232 57666 204241
rect 57610 204167 57666 204176
rect 57532 203510 57652 203538
rect 57518 203416 57574 203425
rect 57518 203351 57574 203360
rect 57426 198792 57482 198801
rect 57426 198727 57482 198736
rect 57334 197024 57390 197033
rect 57334 196959 57390 196968
rect 57242 97472 57298 97481
rect 57242 97407 57298 97416
rect 57348 90545 57376 196959
rect 57440 93401 57468 198727
rect 57532 96529 57560 203351
rect 57624 200841 57652 203510
rect 57610 200832 57666 200841
rect 57610 200767 57666 200776
rect 57518 96520 57574 96529
rect 57518 96455 57574 96464
rect 57624 93809 57652 200767
rect 57716 199889 57744 306711
rect 57794 305008 57850 305017
rect 57794 304943 57850 304952
rect 57702 199880 57758 199889
rect 57702 199815 57758 199824
rect 57716 198801 57744 199815
rect 57702 198792 57758 198801
rect 57702 198727 57758 198736
rect 57808 198234 57836 304943
rect 58440 300824 58492 300830
rect 58440 300766 58492 300772
rect 57886 282568 57942 282577
rect 57886 282503 57942 282512
rect 57716 198206 57836 198234
rect 57716 198121 57744 198206
rect 57702 198112 57758 198121
rect 57702 198047 57758 198056
rect 57610 93800 57666 93809
rect 57610 93735 57666 93744
rect 57426 93392 57482 93401
rect 57426 93327 57482 93336
rect 57716 91089 57744 198047
rect 57794 195256 57850 195265
rect 57794 195191 57850 195200
rect 57702 91080 57758 91089
rect 57702 91015 57758 91024
rect 57334 90536 57390 90545
rect 57334 90471 57390 90480
rect 57808 88233 57836 195191
rect 57900 175817 57928 282503
rect 58348 282192 58400 282198
rect 58348 282134 58400 282140
rect 58360 272202 58388 282134
rect 58452 272950 58480 300766
rect 58440 272944 58492 272950
rect 58440 272886 58492 272892
rect 58544 272513 58572 357342
rect 58636 284209 58664 472602
rect 58622 284200 58678 284209
rect 58622 284135 58678 284144
rect 58624 282668 58676 282674
rect 58624 282610 58676 282616
rect 58530 272504 58586 272513
rect 58530 272439 58586 272448
rect 58348 272196 58400 272202
rect 58348 272138 58400 272144
rect 58636 272134 58664 282610
rect 58728 282033 58756 482054
rect 58808 465792 58860 465798
rect 58808 465734 58860 465740
rect 58714 282024 58770 282033
rect 58714 281959 58770 281968
rect 58624 272128 58676 272134
rect 58624 272070 58676 272076
rect 57980 270088 58032 270094
rect 57980 270030 58032 270036
rect 57992 269006 58020 270030
rect 58636 270026 58664 272070
rect 58624 270020 58676 270026
rect 58624 269962 58676 269968
rect 57980 269000 58032 269006
rect 57980 268942 58032 268948
rect 57886 175808 57942 175817
rect 57886 175743 57942 175752
rect 57794 88224 57850 88233
rect 57794 88159 57850 88168
rect 57612 70372 57664 70378
rect 57612 70314 57664 70320
rect 57624 70145 57652 70314
rect 57610 70136 57666 70145
rect 57610 70071 57666 70080
rect 57900 68921 57928 175743
rect 57992 146266 58020 268942
rect 58716 268456 58768 268462
rect 58716 268398 58768 268404
rect 58072 267708 58124 267714
rect 58072 267650 58124 267656
rect 58084 267238 58112 267650
rect 58728 267238 58756 268398
rect 58072 267232 58124 267238
rect 58072 267174 58124 267180
rect 58716 267232 58768 267238
rect 58716 267174 58768 267180
rect 58084 149054 58112 267174
rect 58624 252136 58676 252142
rect 58624 252078 58676 252084
rect 58636 164218 58664 252078
rect 58716 251796 58768 251802
rect 58716 251738 58768 251744
rect 58624 164212 58676 164218
rect 58624 164154 58676 164160
rect 58162 164112 58218 164121
rect 58162 164047 58164 164056
rect 58216 164047 58218 164056
rect 58164 164018 58216 164024
rect 58072 149048 58124 149054
rect 58072 148990 58124 148996
rect 58084 147801 58112 148990
rect 58728 148986 58756 251738
rect 58820 177585 58848 465734
rect 58992 464772 59044 464778
rect 58992 464714 59044 464720
rect 58900 464704 58952 464710
rect 58900 464646 58952 464652
rect 58806 177576 58862 177585
rect 58806 177511 58862 177520
rect 58912 166462 58940 464646
rect 59004 166666 59032 464714
rect 58992 166660 59044 166666
rect 58992 166602 59044 166608
rect 59096 166530 59124 485522
rect 59372 474026 59400 488022
rect 60004 485716 60056 485722
rect 60004 485658 60056 485664
rect 59728 480004 59780 480010
rect 59728 479946 59780 479952
rect 59636 477488 59688 477494
rect 59636 477430 59688 477436
rect 59360 474020 59412 474026
rect 59360 473962 59412 473968
rect 59268 467084 59320 467090
rect 59268 467026 59320 467032
rect 59176 467016 59228 467022
rect 59176 466958 59228 466964
rect 59084 166524 59136 166530
rect 59084 166466 59136 166472
rect 58900 166456 58952 166462
rect 58900 166398 58952 166404
rect 59084 162852 59136 162858
rect 59084 162794 59136 162800
rect 59096 162178 59124 162794
rect 59084 162172 59136 162178
rect 59084 162114 59136 162120
rect 58716 148980 58768 148986
rect 58716 148922 58768 148928
rect 58070 147792 58126 147801
rect 58070 147727 58126 147736
rect 58728 147694 58756 148922
rect 58992 148708 59044 148714
rect 58992 148650 59044 148656
rect 58716 147688 58768 147694
rect 58716 147630 58768 147636
rect 57980 146260 58032 146266
rect 57980 146202 58032 146208
rect 58808 145920 58860 145926
rect 58808 145862 58860 145868
rect 58714 145752 58770 145761
rect 58714 145687 58770 145696
rect 58624 145648 58676 145654
rect 58624 145590 58676 145596
rect 58636 144838 58664 145590
rect 58624 144832 58676 144838
rect 58624 144774 58676 144780
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57900 57934 57928 68847
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57900 57186 57928 57870
rect 57244 57180 57296 57186
rect 57244 57122 57296 57128
rect 57888 57180 57940 57186
rect 57888 57122 57940 57128
rect 57060 54800 57112 54806
rect 57060 54742 57112 54748
rect 53656 54732 53708 54738
rect 53656 54674 53708 54680
rect 52184 54596 52236 54602
rect 52184 54538 52236 54544
rect 44088 54528 44140 54534
rect 44088 54470 44140 54476
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 10324 20664 10376 20670
rect 10324 20606 10376 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 57256 3466 57284 57122
rect 58636 54670 58664 144774
rect 58728 144634 58756 145687
rect 58820 144906 58848 145862
rect 58898 145616 58954 145625
rect 58898 145551 58954 145560
rect 58808 144900 58860 144906
rect 58808 144842 58860 144848
rect 58716 144628 58768 144634
rect 58716 144570 58768 144576
rect 58728 56302 58756 144570
rect 58716 56296 58768 56302
rect 58716 56238 58768 56244
rect 58820 56098 58848 144842
rect 58912 144566 58940 145551
rect 58900 144560 58952 144566
rect 58900 144502 58952 144508
rect 58912 59566 58940 144502
rect 58900 59560 58952 59566
rect 58900 59502 58952 59508
rect 59004 58886 59032 148650
rect 59096 59294 59124 162114
rect 59084 59288 59136 59294
rect 59084 59230 59136 59236
rect 58992 58880 59044 58886
rect 58992 58822 59044 58828
rect 59188 57322 59216 466958
rect 59280 57390 59308 467026
rect 59648 416226 59676 477430
rect 59636 416220 59688 416226
rect 59636 416162 59688 416168
rect 59542 388512 59598 388521
rect 59542 388447 59598 388456
rect 59360 381744 59412 381750
rect 59360 381686 59412 381692
rect 59372 358086 59400 381686
rect 59452 380996 59504 381002
rect 59452 380938 59504 380944
rect 59464 358698 59492 380938
rect 59556 378049 59584 388447
rect 59636 381880 59688 381886
rect 59636 381822 59688 381828
rect 59542 378040 59598 378049
rect 59542 377975 59598 377984
rect 59452 358692 59504 358698
rect 59452 358634 59504 358640
rect 59360 358080 59412 358086
rect 59360 358022 59412 358028
rect 59648 272338 59676 381822
rect 59740 379166 59768 479946
rect 59820 476672 59872 476678
rect 59820 476614 59872 476620
rect 59728 379160 59780 379166
rect 59728 379102 59780 379108
rect 59832 272649 59860 476614
rect 59912 468648 59964 468654
rect 59912 468590 59964 468596
rect 59818 272640 59874 272649
rect 59818 272575 59874 272584
rect 59636 272332 59688 272338
rect 59636 272274 59688 272280
rect 59728 272196 59780 272202
rect 59728 272138 59780 272144
rect 59360 164008 59412 164014
rect 59360 163950 59412 163956
rect 59372 163606 59400 163950
rect 59360 163600 59412 163606
rect 59360 163542 59412 163548
rect 59372 140865 59400 163542
rect 59740 146169 59768 272138
rect 59818 271144 59874 271153
rect 59818 271079 59874 271088
rect 59832 270609 59860 271079
rect 59818 270600 59874 270609
rect 59818 270535 59874 270544
rect 59832 146266 59860 270535
rect 59924 165209 59952 468590
rect 60016 166598 60044 485658
rect 60660 483682 60688 488022
rect 60844 488022 61042 488050
rect 61120 488022 61502 488050
rect 61672 488022 61962 488050
rect 62224 488022 62330 488050
rect 62408 488022 62790 488050
rect 62960 488022 63250 488050
rect 63512 488022 63710 488050
rect 60648 483676 60700 483682
rect 60648 483618 60700 483624
rect 60740 477964 60792 477970
rect 60740 477906 60792 477912
rect 60752 466002 60780 477906
rect 60844 475386 60872 488022
rect 61120 477970 61148 488022
rect 61672 478174 61700 488022
rect 62120 480888 62172 480894
rect 62120 480830 62172 480836
rect 61660 478168 61712 478174
rect 61660 478110 61712 478116
rect 61108 477964 61160 477970
rect 61108 477906 61160 477912
rect 60832 475380 60884 475386
rect 60832 475322 60884 475328
rect 62132 466206 62160 480830
rect 62120 466200 62172 466206
rect 62120 466142 62172 466148
rect 60740 465996 60792 466002
rect 60740 465938 60792 465944
rect 62224 465934 62252 488022
rect 62408 479534 62436 488022
rect 62960 480894 62988 488022
rect 63222 485344 63278 485353
rect 63222 485279 63278 485288
rect 63236 484809 63264 485279
rect 63222 484800 63278 484809
rect 63222 484735 63278 484744
rect 62948 480888 63000 480894
rect 62948 480830 63000 480836
rect 62396 479528 62448 479534
rect 62396 479470 62448 479476
rect 63512 466138 63540 488022
rect 64156 485518 64184 488036
rect 64248 488022 64538 488050
rect 65014 488022 65104 488050
rect 64144 485512 64196 485518
rect 64144 485454 64196 485460
rect 64248 470594 64276 488022
rect 64880 487076 64932 487082
rect 64880 487018 64932 487024
rect 64892 471986 64920 487018
rect 65076 485774 65104 488022
rect 65168 488022 65458 488050
rect 65536 488022 65918 488050
rect 65168 487082 65196 488022
rect 65156 487076 65208 487082
rect 65156 487018 65208 487024
rect 65076 485746 65196 485774
rect 65168 476114 65196 485746
rect 65430 485616 65486 485625
rect 65430 485551 65486 485560
rect 65444 485353 65472 485551
rect 65430 485344 65486 485353
rect 65430 485279 65486 485288
rect 64984 476086 65196 476114
rect 64880 471980 64932 471986
rect 64880 471922 64932 471928
rect 64984 471170 65012 476086
rect 65536 471238 65564 488022
rect 66364 482769 66392 488036
rect 66456 488022 66746 488050
rect 66824 488022 67206 488050
rect 67682 488022 67772 488050
rect 66350 482760 66406 482769
rect 66350 482695 66406 482704
rect 66456 476114 66484 488022
rect 66272 476086 66484 476114
rect 65524 471232 65576 471238
rect 65524 471174 65576 471180
rect 64972 471164 65024 471170
rect 64972 471106 65024 471112
rect 63604 470566 64276 470594
rect 63604 469062 63632 470566
rect 63592 469056 63644 469062
rect 63592 468998 63644 469004
rect 63500 466132 63552 466138
rect 63500 466074 63552 466080
rect 66272 466070 66300 476086
rect 66824 470594 66852 488022
rect 67744 481098 67772 488022
rect 67836 488022 68126 488050
rect 68204 488022 68494 488050
rect 67732 481092 67784 481098
rect 67732 481034 67784 481040
rect 67836 475946 67864 488022
rect 67916 481092 67968 481098
rect 67916 481034 67968 481040
rect 66364 470566 66852 470594
rect 67652 475918 67864 475946
rect 66364 467022 66392 470566
rect 66352 467016 66404 467022
rect 66352 466958 66404 466964
rect 66260 466064 66312 466070
rect 66260 466006 66312 466012
rect 62212 465928 62264 465934
rect 62212 465870 62264 465876
rect 67652 465633 67680 475918
rect 67928 473354 67956 481034
rect 67744 473326 67956 473354
rect 67744 467090 67772 473326
rect 68204 470594 68232 488022
rect 68940 484945 68968 488036
rect 69032 488022 69414 488050
rect 69492 488022 69874 488050
rect 69952 488022 70334 488050
rect 70596 488022 70702 488050
rect 70872 488022 71162 488050
rect 71240 488022 71622 488050
rect 71792 488022 72082 488050
rect 68926 484936 68982 484945
rect 68926 484871 68982 484880
rect 68284 484764 68336 484770
rect 68284 484706 68336 484712
rect 68296 471102 68324 484706
rect 68284 471096 68336 471102
rect 68284 471038 68336 471044
rect 67836 470566 68232 470594
rect 67836 468353 67864 470566
rect 67822 468344 67878 468353
rect 67822 468279 67878 468288
rect 67732 467084 67784 467090
rect 67732 467026 67784 467032
rect 69032 466449 69060 488022
rect 69112 480888 69164 480894
rect 69112 480830 69164 480836
rect 69124 469033 69152 480830
rect 69492 470594 69520 488022
rect 69952 480894 69980 488022
rect 70492 484220 70544 484226
rect 70492 484162 70544 484168
rect 70400 484152 70452 484158
rect 70400 484094 70452 484100
rect 69940 480888 69992 480894
rect 69940 480830 69992 480836
rect 69216 470566 69520 470594
rect 69110 469024 69166 469033
rect 69110 468959 69166 468968
rect 69216 468897 69244 470566
rect 69202 468888 69258 468897
rect 69202 468823 69258 468832
rect 69018 466440 69074 466449
rect 69018 466375 69074 466384
rect 70412 465730 70440 484094
rect 70504 467129 70532 484162
rect 70596 468994 70624 488022
rect 70872 484158 70900 488022
rect 71240 484226 71268 488022
rect 71228 484220 71280 484226
rect 71228 484162 71280 484168
rect 70860 484152 70912 484158
rect 70860 484094 70912 484100
rect 70584 468988 70636 468994
rect 70584 468930 70636 468936
rect 70490 467120 70546 467129
rect 70490 467055 70546 467064
rect 71792 466313 71820 488022
rect 72528 485625 72556 488036
rect 72620 488022 72910 488050
rect 73172 488022 73370 488050
rect 72514 485616 72570 485625
rect 72514 485551 72570 485560
rect 72424 485512 72476 485518
rect 72424 485454 72476 485460
rect 71872 484152 71924 484158
rect 71872 484094 71924 484100
rect 71884 467265 71912 484094
rect 71870 467256 71926 467265
rect 71870 467191 71926 467200
rect 71778 466304 71834 466313
rect 71778 466239 71834 466248
rect 72436 465730 72464 485454
rect 72620 484158 72648 488022
rect 72608 484152 72660 484158
rect 72608 484094 72660 484100
rect 73172 469169 73200 488022
rect 73342 485616 73398 485625
rect 73342 485551 73398 485560
rect 73250 485480 73306 485489
rect 73250 485415 73306 485424
rect 73264 484974 73292 485415
rect 73252 484968 73304 484974
rect 73252 484910 73304 484916
rect 73356 484838 73384 485551
rect 73816 485353 73844 488036
rect 73988 485784 74040 485790
rect 73988 485726 74040 485732
rect 73802 485344 73858 485353
rect 73802 485279 73858 485288
rect 73804 484968 73856 484974
rect 73804 484910 73856 484916
rect 73344 484832 73396 484838
rect 73344 484774 73396 484780
rect 73158 469160 73214 469169
rect 73158 469095 73214 469104
rect 73816 467838 73844 484910
rect 73896 484900 73948 484906
rect 73896 484842 73948 484848
rect 73804 467832 73856 467838
rect 73804 467774 73856 467780
rect 73908 467702 73936 484842
rect 74000 467770 74028 485726
rect 74276 484809 74304 488036
rect 74552 488022 74658 488050
rect 74736 488022 75118 488050
rect 75288 488022 75578 488050
rect 74262 484800 74318 484809
rect 74262 484735 74318 484744
rect 73988 467764 74040 467770
rect 73988 467706 74040 467712
rect 73896 467696 73948 467702
rect 73896 467638 73948 467644
rect 74552 465905 74580 488022
rect 74632 484152 74684 484158
rect 74632 484094 74684 484100
rect 74644 466177 74672 484094
rect 74630 466168 74686 466177
rect 74630 466103 74686 466112
rect 74538 465896 74594 465905
rect 74538 465831 74594 465840
rect 74736 465769 74764 488022
rect 75288 484158 75316 488022
rect 76024 485761 76052 488036
rect 76208 488022 76498 488050
rect 76576 488022 76866 488050
rect 76010 485752 76066 485761
rect 76010 485687 76066 485696
rect 75276 484152 75328 484158
rect 75276 484094 75328 484100
rect 75920 484152 75972 484158
rect 75920 484094 75972 484100
rect 75932 466342 75960 484094
rect 76208 470594 76236 488022
rect 76576 484158 76604 488022
rect 77312 485217 77340 488036
rect 77772 485489 77800 488036
rect 77864 488022 78246 488050
rect 77758 485480 77814 485489
rect 77758 485415 77814 485424
rect 77298 485208 77354 485217
rect 77298 485143 77354 485152
rect 76564 484152 76616 484158
rect 76564 484094 76616 484100
rect 77864 470594 77892 488022
rect 78692 485625 78720 488036
rect 78876 488022 79074 488050
rect 79152 488022 79534 488050
rect 79704 488022 79994 488050
rect 80072 488022 80454 488050
rect 80532 488022 80822 488050
rect 80992 488022 81282 488050
rect 78678 485616 78734 485625
rect 78678 485551 78734 485560
rect 78680 484220 78732 484226
rect 78680 484162 78732 484168
rect 76024 470566 76236 470594
rect 77312 470566 77892 470594
rect 75920 466336 75972 466342
rect 75920 466278 75972 466284
rect 76024 466041 76052 470566
rect 77312 466410 77340 470566
rect 78692 468761 78720 484162
rect 78772 484152 78824 484158
rect 78772 484094 78824 484100
rect 78784 469130 78812 484094
rect 78772 469124 78824 469130
rect 78772 469066 78824 469072
rect 78678 468752 78734 468761
rect 78678 468687 78734 468696
rect 78876 468625 78904 488022
rect 79152 484226 79180 488022
rect 79324 485512 79376 485518
rect 79324 485454 79376 485460
rect 79336 484974 79364 485454
rect 79324 484968 79376 484974
rect 79324 484910 79376 484916
rect 79140 484220 79192 484226
rect 79140 484162 79192 484168
rect 79704 484158 79732 488022
rect 79692 484152 79744 484158
rect 79692 484094 79744 484100
rect 80072 469198 80100 488022
rect 80532 480049 80560 488022
rect 80704 483676 80756 483682
rect 80704 483618 80756 483624
rect 80518 480040 80574 480049
rect 80518 479975 80574 479984
rect 80060 469192 80112 469198
rect 80060 469134 80112 469140
rect 78862 468616 78918 468625
rect 78862 468551 78918 468560
rect 80716 467838 80744 483618
rect 80992 476610 81020 488022
rect 81728 485042 81756 488036
rect 81912 488022 82202 488050
rect 82280 488022 82662 488050
rect 82924 488022 83030 488050
rect 83200 488022 83490 488050
rect 83568 488022 83950 488050
rect 81716 485036 81768 485042
rect 81716 484978 81768 484984
rect 81532 480888 81584 480894
rect 81532 480830 81584 480836
rect 80980 476604 81032 476610
rect 80980 476546 81032 476552
rect 81544 469849 81572 480830
rect 81912 470594 81940 488022
rect 82280 480894 82308 488022
rect 82268 480888 82320 480894
rect 82268 480830 82320 480836
rect 82820 480888 82872 480894
rect 82820 480830 82872 480836
rect 82832 471918 82860 480830
rect 82820 471912 82872 471918
rect 82820 471854 82872 471860
rect 82924 471782 82952 488022
rect 82912 471776 82964 471782
rect 82912 471718 82964 471724
rect 83200 471714 83228 488022
rect 83568 480894 83596 488022
rect 84396 484770 84424 488036
rect 84488 488022 84870 488050
rect 84948 488022 85238 488050
rect 85714 488022 85804 488050
rect 84384 484764 84436 484770
rect 84384 484706 84436 484712
rect 83556 480888 83608 480894
rect 83556 480830 83608 480836
rect 84292 480888 84344 480894
rect 84292 480830 84344 480836
rect 83188 471708 83240 471714
rect 83188 471650 83240 471656
rect 84304 471617 84332 480830
rect 84488 471850 84516 488022
rect 84948 480894 84976 488022
rect 85776 483014 85804 488022
rect 85684 482986 85804 483014
rect 85868 488022 86158 488050
rect 86328 488022 86618 488050
rect 86972 488022 87078 488050
rect 87156 488022 87446 488050
rect 87524 488022 87906 488050
rect 84936 480888 84988 480894
rect 84936 480830 84988 480836
rect 85580 480888 85632 480894
rect 85580 480830 85632 480836
rect 84476 471844 84528 471850
rect 84476 471786 84528 471792
rect 84290 471608 84346 471617
rect 84290 471543 84346 471552
rect 81636 470566 81940 470594
rect 81636 469946 81664 470566
rect 81624 469940 81676 469946
rect 81624 469882 81676 469888
rect 81530 469840 81586 469849
rect 81530 469775 81586 469784
rect 85592 468926 85620 480830
rect 85684 478122 85712 482986
rect 85684 478094 85804 478122
rect 85672 474632 85724 474638
rect 85672 474574 85724 474580
rect 85580 468920 85632 468926
rect 85580 468862 85632 468868
rect 85684 468722 85712 474574
rect 85776 471345 85804 478094
rect 85868 474638 85896 488022
rect 86328 480894 86356 488022
rect 86316 480888 86368 480894
rect 86316 480830 86368 480836
rect 85856 474632 85908 474638
rect 85856 474574 85908 474580
rect 85762 471336 85818 471345
rect 85762 471271 85818 471280
rect 86972 468790 87000 488022
rect 87156 476114 87184 488022
rect 87064 476086 87184 476114
rect 86960 468784 87012 468790
rect 86960 468726 87012 468732
rect 85672 468716 85724 468722
rect 85672 468658 85724 468664
rect 87064 468586 87092 476086
rect 87524 470594 87552 488022
rect 88352 485450 88380 488036
rect 88536 488022 88826 488050
rect 88904 488022 89194 488050
rect 88340 485444 88392 485450
rect 88340 485386 88392 485392
rect 88432 476468 88484 476474
rect 88432 476410 88484 476416
rect 88444 471209 88472 476410
rect 88536 471481 88564 488022
rect 88904 476474 88932 488022
rect 89640 485654 89668 488036
rect 89824 488022 90114 488050
rect 89628 485648 89680 485654
rect 89628 485590 89680 485596
rect 88892 476468 88944 476474
rect 88892 476410 88944 476416
rect 88522 471472 88578 471481
rect 88522 471407 88578 471416
rect 88430 471200 88486 471209
rect 88430 471135 88486 471144
rect 87156 470566 87552 470594
rect 87156 468858 87184 470566
rect 87144 468852 87196 468858
rect 87144 468794 87196 468800
rect 87052 468580 87104 468586
rect 87052 468522 87104 468528
rect 80704 467832 80756 467838
rect 80704 467774 80756 467780
rect 77300 466404 77352 466410
rect 77300 466346 77352 466352
rect 76010 466032 76066 466041
rect 76010 465967 76066 465976
rect 89824 465866 89852 488022
rect 90560 485382 90588 488036
rect 90744 488022 91034 488050
rect 90548 485376 90600 485382
rect 90548 485318 90600 485324
rect 90744 470594 90772 488022
rect 91388 485081 91416 488036
rect 91848 485722 91876 488036
rect 91836 485716 91888 485722
rect 91836 485658 91888 485664
rect 92308 485586 92336 488036
rect 92584 488022 92782 488050
rect 92860 488022 93242 488050
rect 92296 485580 92348 485586
rect 92296 485522 92348 485528
rect 91374 485072 91430 485081
rect 91374 485007 91430 485016
rect 89916 470566 90772 470594
rect 89812 465860 89864 465866
rect 89812 465802 89864 465808
rect 74722 465760 74778 465769
rect 70400 465724 70452 465730
rect 70400 465666 70452 465672
rect 72424 465724 72476 465730
rect 74722 465695 74778 465704
rect 72424 465666 72476 465672
rect 67638 465624 67694 465633
rect 67638 465559 67694 465568
rect 89916 464778 89944 470566
rect 92584 468654 92612 488022
rect 92860 470594 92888 488022
rect 93596 485314 93624 488036
rect 93964 488022 94070 488050
rect 94240 488022 94530 488050
rect 94608 488022 94990 488050
rect 93584 485308 93636 485314
rect 93584 485250 93636 485256
rect 93860 484152 93912 484158
rect 93860 484094 93912 484100
rect 92676 470566 92888 470594
rect 92572 468648 92624 468654
rect 92572 468590 92624 468596
rect 89904 464772 89956 464778
rect 89904 464714 89956 464720
rect 92676 464710 92704 470566
rect 93872 467498 93900 484094
rect 93964 468518 93992 488022
rect 94240 470594 94268 488022
rect 94608 484158 94636 488022
rect 95344 484906 95372 488036
rect 95436 488022 95818 488050
rect 95332 484900 95384 484906
rect 95332 484842 95384 484848
rect 94596 484152 94648 484158
rect 94596 484094 94648 484100
rect 94056 470566 94268 470594
rect 93952 468512 94004 468518
rect 94056 468489 94084 470566
rect 93952 468454 94004 468460
rect 94042 468480 94098 468489
rect 94042 468415 94098 468424
rect 93860 467492 93912 467498
rect 93860 467434 93912 467440
rect 95436 465798 95464 488022
rect 96264 482118 96292 488036
rect 96724 482186 96752 488036
rect 97184 483002 97212 488036
rect 97172 482996 97224 483002
rect 97172 482938 97224 482944
rect 97552 482934 97580 488036
rect 97540 482928 97592 482934
rect 97540 482870 97592 482876
rect 98012 482866 98040 488036
rect 98000 482860 98052 482866
rect 98000 482802 98052 482808
rect 98472 482254 98500 488036
rect 98656 488022 98946 488050
rect 98460 482248 98512 482254
rect 98460 482190 98512 482196
rect 96712 482180 96764 482186
rect 96712 482122 96764 482128
rect 96252 482112 96304 482118
rect 96252 482054 96304 482060
rect 98656 471374 98684 488022
rect 99392 485246 99420 488036
rect 99576 488022 99774 488050
rect 99944 488022 100234 488050
rect 100312 488022 100694 488050
rect 100956 488022 101154 488050
rect 101232 488022 101522 488050
rect 101600 488022 101982 488050
rect 102244 488022 102442 488050
rect 99380 485240 99432 485246
rect 99380 485182 99432 485188
rect 99472 480888 99524 480894
rect 99472 480830 99524 480836
rect 98644 471368 98696 471374
rect 98644 471310 98696 471316
rect 99484 467566 99512 480830
rect 99576 474162 99604 488022
rect 99564 474156 99616 474162
rect 99564 474098 99616 474104
rect 99944 470594 99972 488022
rect 100312 480894 100340 488022
rect 100300 480888 100352 480894
rect 100300 480830 100352 480836
rect 100760 480888 100812 480894
rect 100760 480830 100812 480836
rect 100772 471646 100800 480830
rect 100852 476536 100904 476542
rect 100852 476478 100904 476484
rect 100760 471640 100812 471646
rect 100760 471582 100812 471588
rect 100864 471510 100892 476478
rect 100852 471504 100904 471510
rect 100852 471446 100904 471452
rect 100956 471442 100984 488022
rect 101232 476542 101260 488022
rect 101600 480894 101628 488022
rect 101588 480888 101640 480894
rect 101588 480830 101640 480836
rect 101220 476536 101272 476542
rect 101220 476478 101272 476484
rect 100944 471436 100996 471442
rect 100944 471378 100996 471384
rect 99668 470566 99972 470594
rect 99668 467634 99696 470566
rect 99656 467628 99708 467634
rect 99656 467570 99708 467576
rect 99472 467560 99524 467566
rect 99472 467502 99524 467508
rect 95424 465792 95476 465798
rect 95424 465734 95476 465740
rect 92664 464704 92716 464710
rect 92664 464646 92716 464652
rect 102244 464574 102272 488022
rect 102888 485178 102916 488036
rect 103072 488022 103362 488050
rect 103624 488022 103730 488050
rect 103808 488022 104190 488050
rect 102876 485172 102928 485178
rect 102876 485114 102928 485120
rect 103072 470594 103100 488022
rect 103624 471578 103652 488022
rect 103612 471572 103664 471578
rect 103612 471514 103664 471520
rect 103808 470594 103836 488022
rect 104636 485110 104664 488036
rect 105096 485790 105124 488036
rect 105188 488022 105570 488050
rect 105648 488022 105938 488050
rect 105084 485784 105136 485790
rect 105084 485726 105136 485732
rect 104624 485104 104676 485110
rect 104624 485046 104676 485052
rect 105188 476114 105216 488022
rect 102336 470566 103100 470594
rect 103716 470566 103836 470594
rect 105004 476086 105216 476114
rect 102336 464642 102364 470566
rect 103716 467362 103744 470566
rect 103704 467356 103756 467362
rect 103704 467298 103756 467304
rect 105004 467294 105032 476086
rect 105648 470594 105676 488022
rect 106384 485518 106412 488036
rect 106476 488022 106858 488050
rect 106936 488022 107318 488050
rect 107794 488022 107884 488050
rect 106372 485512 106424 485518
rect 106372 485454 106424 485460
rect 106372 480888 106424 480894
rect 106372 480830 106424 480836
rect 105096 470566 105676 470594
rect 105096 467430 105124 470566
rect 105084 467424 105136 467430
rect 105084 467366 105136 467372
rect 104992 467288 105044 467294
rect 104992 467230 105044 467236
rect 106384 467226 106412 480830
rect 106372 467220 106424 467226
rect 106372 467162 106424 467168
rect 106476 467158 106504 488022
rect 106936 480894 106964 488022
rect 107856 485790 107884 488022
rect 107948 488022 108146 488050
rect 108224 488022 108606 488050
rect 109082 488022 109448 488050
rect 107844 485784 107896 485790
rect 107844 485726 107896 485732
rect 106924 480888 106976 480894
rect 107948 480842 107976 488022
rect 108028 485784 108080 485790
rect 108028 485726 108080 485732
rect 106924 480830 106976 480836
rect 107672 480814 107976 480842
rect 106464 467152 106516 467158
rect 106464 467094 106516 467100
rect 107672 465798 107700 480814
rect 107752 478576 107804 478582
rect 107752 478518 107804 478524
rect 107764 468518 107792 478518
rect 108040 470594 108068 485726
rect 108224 478582 108252 488022
rect 109420 486606 109448 488022
rect 109408 486600 109460 486606
rect 109408 486542 109460 486548
rect 109512 486538 109540 488036
rect 109604 488022 109894 488050
rect 109500 486532 109552 486538
rect 109500 486474 109552 486480
rect 108212 478576 108264 478582
rect 108212 478518 108264 478524
rect 109604 470594 109632 488022
rect 110340 485110 110368 488036
rect 110616 488022 110814 488050
rect 110328 485104 110380 485110
rect 110328 485046 110380 485052
rect 110616 472666 110644 488022
rect 111260 482730 111288 488036
rect 111720 482798 111748 488036
rect 111708 482792 111760 482798
rect 111708 482734 111760 482740
rect 111248 482724 111300 482730
rect 111248 482666 111300 482672
rect 112088 482526 112116 488036
rect 112548 482594 112576 488036
rect 112640 488022 113022 488050
rect 112536 482588 112588 482594
rect 112536 482530 112588 482536
rect 112076 482520 112128 482526
rect 112076 482462 112128 482468
rect 110604 472660 110656 472666
rect 110604 472602 110656 472608
rect 112640 470594 112668 488022
rect 113272 480888 113324 480894
rect 113272 480830 113324 480836
rect 113284 474094 113312 480830
rect 113468 476114 113496 488036
rect 113560 488022 113942 488050
rect 113560 480894 113588 488022
rect 114296 481030 114324 488036
rect 114284 481024 114336 481030
rect 114284 480966 114336 480972
rect 113548 480888 113600 480894
rect 113548 480830 113600 480836
rect 113376 476086 113496 476114
rect 113272 474088 113324 474094
rect 113272 474030 113324 474036
rect 113376 471306 113404 476086
rect 114756 475454 114784 488036
rect 115216 482458 115244 488036
rect 115676 482662 115704 488036
rect 116074 488022 116164 488050
rect 115664 482656 115716 482662
rect 115664 482598 115716 482604
rect 115204 482452 115256 482458
rect 115204 482394 115256 482400
rect 116136 479466 116164 488022
rect 116228 488022 116518 488050
rect 116688 488022 116978 488050
rect 117454 488022 117544 488050
rect 116228 480146 116256 488022
rect 116216 480140 116268 480146
rect 116216 480082 116268 480088
rect 116124 479460 116176 479466
rect 116124 479402 116176 479408
rect 116688 479330 116716 488022
rect 117516 480078 117544 488022
rect 117608 488022 117898 488050
rect 117976 488022 118266 488050
rect 117504 480072 117556 480078
rect 117504 480014 117556 480020
rect 117608 479942 117636 488022
rect 117596 479936 117648 479942
rect 117596 479878 117648 479884
rect 117976 479874 118004 488022
rect 118712 479913 118740 488036
rect 118804 488022 119186 488050
rect 118698 479904 118754 479913
rect 117964 479868 118016 479874
rect 118698 479839 118754 479848
rect 117964 479810 118016 479816
rect 118804 479641 118832 488022
rect 119632 482390 119660 488036
rect 119620 482384 119672 482390
rect 119620 482326 119672 482332
rect 120092 482322 120120 488036
rect 120460 482497 120488 488036
rect 120950 488022 121224 488050
rect 121196 486674 121224 488022
rect 121184 486668 121236 486674
rect 121184 486610 121236 486616
rect 121380 482633 121408 488036
rect 121472 488022 121854 488050
rect 121932 488022 122222 488050
rect 122392 488022 122682 488050
rect 123036 488022 123142 488050
rect 123312 488022 123602 488050
rect 123680 488022 124062 488050
rect 124232 488022 124430 488050
rect 124508 488022 124890 488050
rect 124968 488022 125350 488050
rect 121366 482624 121422 482633
rect 121366 482559 121422 482568
rect 120446 482488 120502 482497
rect 120446 482423 120502 482432
rect 120080 482316 120132 482322
rect 120080 482258 120132 482264
rect 118790 479632 118846 479641
rect 118790 479567 118846 479576
rect 116676 479324 116728 479330
rect 116676 479266 116728 479272
rect 114744 475448 114796 475454
rect 114744 475390 114796 475396
rect 113364 471300 113416 471306
rect 113364 471242 113416 471248
rect 107856 470566 108068 470594
rect 109052 470566 109632 470594
rect 111996 470566 112668 470594
rect 107856 468586 107884 470566
rect 109052 468654 109080 470566
rect 111996 469878 112024 470566
rect 111984 469872 112036 469878
rect 111984 469814 112036 469820
rect 109040 468648 109092 468654
rect 109040 468590 109092 468596
rect 107844 468580 107896 468586
rect 107844 468522 107896 468528
rect 107752 468512 107804 468518
rect 107752 468454 107804 468460
rect 107660 465792 107712 465798
rect 107660 465734 107712 465740
rect 102324 464636 102376 464642
rect 102324 464578 102376 464584
rect 102232 464568 102284 464574
rect 102232 464510 102284 464516
rect 121472 464506 121500 488022
rect 121932 479777 121960 488022
rect 121918 479768 121974 479777
rect 121918 479703 121974 479712
rect 122392 479505 122420 488022
rect 123036 480214 123064 488022
rect 123024 480208 123076 480214
rect 123024 480150 123076 480156
rect 122378 479496 122434 479505
rect 122378 479431 122434 479440
rect 123312 477426 123340 488022
rect 123680 479398 123708 488022
rect 123668 479392 123720 479398
rect 123668 479334 123720 479340
rect 123300 477420 123352 477426
rect 123300 477362 123352 477368
rect 124232 477193 124260 488022
rect 124218 477184 124274 477193
rect 124218 477119 124274 477128
rect 124508 476785 124536 488022
rect 124968 476921 124996 488022
rect 125600 480888 125652 480894
rect 125600 480830 125652 480836
rect 124954 476912 125010 476921
rect 124954 476847 125010 476856
rect 124494 476776 124550 476785
rect 124494 476711 124550 476720
rect 125612 464506 125640 480830
rect 125796 477057 125824 488036
rect 125888 488022 126270 488050
rect 126348 488022 126638 488050
rect 125782 477048 125838 477057
rect 125782 476983 125838 476992
rect 125888 476114 125916 488022
rect 126348 480894 126376 488022
rect 127084 482361 127112 488036
rect 127176 488022 127558 488050
rect 127636 488022 128018 488050
rect 128494 488022 128584 488050
rect 127070 482352 127126 482361
rect 127070 482287 127126 482296
rect 126336 480888 126388 480894
rect 126336 480830 126388 480836
rect 127176 476114 127204 488022
rect 127636 476678 127664 488022
rect 128360 487076 128412 487082
rect 128360 487018 128412 487024
rect 128372 477329 128400 487018
rect 128556 485774 128584 488022
rect 128648 488022 128846 488050
rect 128924 488022 129306 488050
rect 129782 488022 129872 488050
rect 128648 487082 128676 488022
rect 128636 487076 128688 487082
rect 128636 487018 128688 487024
rect 128556 485746 128676 485774
rect 128648 483970 128676 485746
rect 128464 483942 128676 483970
rect 128358 477320 128414 477329
rect 128358 477255 128414 477264
rect 128464 476746 128492 483942
rect 128924 479670 128952 488022
rect 129844 484362 129872 488022
rect 129936 488022 130226 488050
rect 130304 488022 130594 488050
rect 130672 488022 131054 488050
rect 131224 488022 131514 488050
rect 131592 488022 131974 488050
rect 132144 488022 132434 488050
rect 132512 488022 132802 488050
rect 132880 488022 133262 488050
rect 133432 488022 133722 488050
rect 133984 488022 134182 488050
rect 134352 488022 134642 488050
rect 134720 488022 135010 488050
rect 135486 488022 135668 488050
rect 129832 484356 129884 484362
rect 129832 484298 129884 484304
rect 129936 484294 129964 488022
rect 130016 484356 130068 484362
rect 130016 484298 130068 484304
rect 129740 484288 129792 484294
rect 129740 484230 129792 484236
rect 129924 484288 129976 484294
rect 129924 484230 129976 484236
rect 129752 479806 129780 484230
rect 130028 484106 130056 484298
rect 129936 484078 130056 484106
rect 129832 484016 129884 484022
rect 129832 483958 129884 483964
rect 129844 480010 129872 483958
rect 129832 480004 129884 480010
rect 129832 479946 129884 479952
rect 129740 479800 129792 479806
rect 129740 479742 129792 479748
rect 129936 479738 129964 484078
rect 130304 484022 130332 488022
rect 130292 484016 130344 484022
rect 130292 483958 130344 483964
rect 129924 479732 129976 479738
rect 129924 479674 129976 479680
rect 128912 479664 128964 479670
rect 128912 479606 128964 479612
rect 130672 477086 130700 488022
rect 131120 484152 131172 484158
rect 131120 484094 131172 484100
rect 130660 477080 130712 477086
rect 130660 477022 130712 477028
rect 128452 476740 128504 476746
rect 128452 476682 128504 476688
rect 127624 476672 127676 476678
rect 127624 476614 127676 476620
rect 125704 476086 125916 476114
rect 126992 476086 127204 476114
rect 125704 471306 125732 476086
rect 126992 474094 127020 476086
rect 126980 474088 127032 474094
rect 126980 474030 127032 474036
rect 125692 471300 125744 471306
rect 125692 471242 125744 471248
rect 121460 464500 121512 464506
rect 121460 464442 121512 464448
rect 125600 464500 125652 464506
rect 125600 464442 125652 464448
rect 131132 464438 131160 484094
rect 131224 477154 131252 488022
rect 131212 477148 131264 477154
rect 131212 477090 131264 477096
rect 131592 476882 131620 488022
rect 132144 484158 132172 488022
rect 132132 484152 132184 484158
rect 132132 484094 132184 484100
rect 131580 476876 131632 476882
rect 131580 476818 131632 476824
rect 131120 464432 131172 464438
rect 131120 464374 131172 464380
rect 132512 464370 132540 488022
rect 132592 484152 132644 484158
rect 132592 484094 132644 484100
rect 132604 477018 132632 484094
rect 132592 477012 132644 477018
rect 132592 476954 132644 476960
rect 132880 476950 132908 488022
rect 133432 484158 133460 488022
rect 133420 484152 133472 484158
rect 133420 484094 133472 484100
rect 133880 484152 133932 484158
rect 133880 484094 133932 484100
rect 133892 477290 133920 484094
rect 133880 477284 133932 477290
rect 133880 477226 133932 477232
rect 133984 477222 134012 488022
rect 134352 479602 134380 488022
rect 134720 484158 134748 488022
rect 134708 484152 134760 484158
rect 134708 484094 134760 484100
rect 135640 482662 135668 488022
rect 135732 488022 135930 488050
rect 136008 488022 136390 488050
rect 136774 488022 136864 488050
rect 135628 482656 135680 482662
rect 135628 482598 135680 482604
rect 135732 482474 135760 488022
rect 135272 482446 135760 482474
rect 134340 479596 134392 479602
rect 134340 479538 134392 479544
rect 135272 477358 135300 482446
rect 136008 477494 136036 488022
rect 136836 482526 136864 488022
rect 136928 488022 137218 488050
rect 137694 488022 137968 488050
rect 138154 488022 138520 488050
rect 136824 482520 136876 482526
rect 136824 482462 136876 482468
rect 135996 477488 136048 477494
rect 135996 477430 136048 477436
rect 135260 477352 135312 477358
rect 135260 477294 135312 477300
rect 133972 477216 134024 477222
rect 133972 477158 134024 477164
rect 132868 476944 132920 476950
rect 132868 476886 132920 476892
rect 136928 470594 136956 488022
rect 137940 482390 137968 488022
rect 138492 482594 138520 488022
rect 138480 482588 138532 482594
rect 138480 482530 138532 482536
rect 137928 482384 137980 482390
rect 137928 482326 137980 482332
rect 138584 482322 138612 488036
rect 138676 488022 138966 488050
rect 138572 482316 138624 482322
rect 138572 482258 138624 482264
rect 138676 470594 138704 488022
rect 139412 484974 139440 488036
rect 139504 488022 139886 488050
rect 140056 488022 140346 488050
rect 140822 488022 140912 488050
rect 139400 484968 139452 484974
rect 139400 484910 139452 484916
rect 139400 484152 139452 484158
rect 139400 484094 139452 484100
rect 136652 470566 136956 470594
rect 138032 470566 138704 470594
rect 136652 464370 136680 470566
rect 138032 464438 138060 470566
rect 139412 468790 139440 484094
rect 139504 474162 139532 488022
rect 140056 484158 140084 488022
rect 140884 486742 140912 488022
rect 140976 488022 141174 488050
rect 141344 488022 141634 488050
rect 141712 488022 142094 488050
rect 142264 488022 142554 488050
rect 142632 488022 142922 488050
rect 143000 488022 143382 488050
rect 143644 488022 143842 488050
rect 144318 488022 144408 488050
rect 140872 486736 140924 486742
rect 140872 486678 140924 486684
rect 140044 484152 140096 484158
rect 140044 484094 140096 484100
rect 140872 484152 140924 484158
rect 140872 484094 140924 484100
rect 140780 482452 140832 482458
rect 140780 482394 140832 482400
rect 139492 474156 139544 474162
rect 139492 474098 139544 474104
rect 140792 471374 140820 482394
rect 140884 471442 140912 484094
rect 140976 471510 141004 488022
rect 141344 484158 141372 488022
rect 141332 484152 141384 484158
rect 141332 484094 141384 484100
rect 141712 482458 141740 488022
rect 142160 484152 142212 484158
rect 142160 484094 142212 484100
rect 141792 482656 141844 482662
rect 141792 482598 141844 482604
rect 141804 482458 141832 482598
rect 141700 482452 141752 482458
rect 141700 482394 141752 482400
rect 141792 482452 141844 482458
rect 141792 482394 141844 482400
rect 140964 471504 141016 471510
rect 140964 471446 141016 471452
rect 140872 471436 140924 471442
rect 140872 471378 140924 471384
rect 140780 471368 140832 471374
rect 140780 471310 140832 471316
rect 139400 468784 139452 468790
rect 139400 468726 139452 468732
rect 142172 464574 142200 484094
rect 142264 465866 142292 488022
rect 142632 484158 142660 488022
rect 142620 484152 142672 484158
rect 142620 484094 142672 484100
rect 143000 470594 143028 488022
rect 143540 484152 143592 484158
rect 143540 484094 143592 484100
rect 142356 470566 143028 470594
rect 142356 468722 142384 470566
rect 143552 469878 143580 484094
rect 143644 476814 143672 488022
rect 144380 483721 144408 488022
rect 144472 488022 144762 488050
rect 145146 488022 145512 488050
rect 145606 488022 145696 488050
rect 144472 484158 144500 488022
rect 145484 485081 145512 488022
rect 145668 485353 145696 488022
rect 145760 488022 146050 488050
rect 146312 488022 146510 488050
rect 146680 488022 146970 488050
rect 147354 488022 147628 488050
rect 145654 485344 145710 485353
rect 145654 485279 145710 485288
rect 145470 485072 145526 485081
rect 145470 485007 145526 485016
rect 144460 484152 144512 484158
rect 144460 484094 144512 484100
rect 144366 483712 144422 483721
rect 144366 483647 144422 483656
rect 143632 476808 143684 476814
rect 143632 476750 143684 476756
rect 145760 472569 145788 488022
rect 145746 472560 145802 472569
rect 145746 472495 145802 472504
rect 143540 469872 143592 469878
rect 143540 469814 143592 469820
rect 142344 468716 142396 468722
rect 142344 468658 142396 468664
rect 146312 467158 146340 488022
rect 146680 479641 146708 488022
rect 147600 485217 147628 488022
rect 147586 485208 147642 485217
rect 147586 485143 147642 485152
rect 147680 484152 147732 484158
rect 147680 484094 147732 484100
rect 146666 479632 146722 479641
rect 146666 479567 146722 479576
rect 147692 472705 147720 484094
rect 147784 478145 147812 488036
rect 148244 485382 148272 488036
rect 148336 488022 148718 488050
rect 149194 488022 149468 488050
rect 148232 485376 148284 485382
rect 148232 485318 148284 485324
rect 148336 484158 148364 488022
rect 149440 485450 149468 488022
rect 149532 485722 149560 488036
rect 149624 488022 150006 488050
rect 149520 485716 149572 485722
rect 149520 485658 149572 485664
rect 149428 485444 149480 485450
rect 149428 485386 149480 485392
rect 148324 484152 148376 484158
rect 148324 484094 148376 484100
rect 147770 478136 147826 478145
rect 147770 478071 147826 478080
rect 147678 472696 147734 472705
rect 147678 472631 147734 472640
rect 149624 470594 149652 488022
rect 150452 485246 150480 488036
rect 150544 488022 150926 488050
rect 150440 485240 150492 485246
rect 150440 485182 150492 485188
rect 150544 484106 150572 488022
rect 151280 485790 151308 488036
rect 151372 488022 151754 488050
rect 151268 485784 151320 485790
rect 151268 485726 151320 485732
rect 150452 484078 150572 484106
rect 150452 474065 150480 484078
rect 151372 476785 151400 488022
rect 152200 485518 152228 488036
rect 152292 488022 152674 488050
rect 152752 488022 153134 488050
rect 153212 488022 153502 488050
rect 153978 488022 154344 488050
rect 154438 488022 154528 488050
rect 154898 488022 155264 488050
rect 155358 488022 155632 488050
rect 155726 488022 155908 488050
rect 152188 485512 152240 485518
rect 152188 485454 152240 485460
rect 152292 484106 152320 488022
rect 151832 484078 152320 484106
rect 151832 478281 151860 484078
rect 152752 479505 152780 488022
rect 152738 479496 152794 479505
rect 152738 479431 152794 479440
rect 151818 478272 151874 478281
rect 151818 478207 151874 478216
rect 151358 476776 151414 476785
rect 151358 476711 151414 476720
rect 150438 474056 150494 474065
rect 150438 473991 150494 474000
rect 149072 470566 149652 470594
rect 149072 467226 149100 470566
rect 149060 467220 149112 467226
rect 149060 467162 149112 467168
rect 146300 467152 146352 467158
rect 153212 467129 153240 488022
rect 154316 485654 154344 488022
rect 154304 485648 154356 485654
rect 154304 485590 154356 485596
rect 154500 480865 154528 488022
rect 155236 482361 155264 488022
rect 155604 484906 155632 488022
rect 155592 484900 155644 484906
rect 155592 484842 155644 484848
rect 155880 483857 155908 488022
rect 155972 488022 156170 488050
rect 156646 488022 156736 488050
rect 155866 483848 155922 483857
rect 155866 483783 155922 483792
rect 155222 482352 155278 482361
rect 155222 482287 155278 482296
rect 154486 480856 154542 480865
rect 154486 480791 154542 480800
rect 155972 474201 156000 488022
rect 156708 485314 156736 488022
rect 156800 488022 157090 488050
rect 156696 485308 156748 485314
rect 156696 485250 156748 485256
rect 156800 475561 156828 488022
rect 157444 485042 157472 488036
rect 157536 488022 157918 488050
rect 158394 488022 158760 488050
rect 158854 488022 159128 488050
rect 157432 485036 157484 485042
rect 157432 484978 157484 484984
rect 157536 476921 157564 488022
rect 158732 484974 158760 488022
rect 158720 484968 158772 484974
rect 158720 484910 158772 484916
rect 159100 481030 159128 488022
rect 159284 482730 159312 488036
rect 159376 488022 159666 488050
rect 160142 488022 160232 488050
rect 159272 482724 159324 482730
rect 159272 482666 159324 482672
rect 159088 481024 159140 481030
rect 159088 480966 159140 480972
rect 157522 476912 157578 476921
rect 157522 476847 157578 476856
rect 156786 475552 156842 475561
rect 156786 475487 156842 475496
rect 159376 474230 159404 488022
rect 160204 479602 160232 488022
rect 160572 482662 160600 488036
rect 160664 488022 161046 488050
rect 160560 482656 160612 482662
rect 160560 482598 160612 482604
rect 160192 479596 160244 479602
rect 160192 479538 160244 479544
rect 160664 476114 160692 488022
rect 161492 485330 161520 488036
rect 161584 488022 161874 488050
rect 161952 488022 162334 488050
rect 162504 488022 162794 488050
rect 162964 488022 163254 488050
rect 163638 488022 163728 488050
rect 161584 485466 161612 488022
rect 161584 485438 161796 485466
rect 161492 485302 161612 485330
rect 161480 485172 161532 485178
rect 161480 485114 161532 485120
rect 161492 484906 161520 485114
rect 161480 484900 161532 484906
rect 161480 484842 161532 484848
rect 161584 483682 161612 485302
rect 161572 483676 161624 483682
rect 161572 483618 161624 483624
rect 161480 480888 161532 480894
rect 161480 480830 161532 480836
rect 160112 476086 160692 476114
rect 159364 474224 159416 474230
rect 155958 474192 156014 474201
rect 159364 474166 159416 474172
rect 155958 474127 156014 474136
rect 160112 468761 160140 476086
rect 160098 468752 160154 468761
rect 160098 468687 160154 468696
rect 161492 468625 161520 480830
rect 161768 476114 161796 485438
rect 161952 480894 161980 488022
rect 162124 485580 162176 485586
rect 162124 485522 162176 485528
rect 162136 485314 162164 485522
rect 162124 485308 162176 485314
rect 162124 485250 162176 485256
rect 162216 485308 162268 485314
rect 162216 485250 162268 485256
rect 162228 485042 162256 485250
rect 162216 485036 162268 485042
rect 162216 484978 162268 484984
rect 161940 480888 161992 480894
rect 161940 480830 161992 480836
rect 161584 476086 161796 476114
rect 161584 471578 161612 476086
rect 161572 471572 161624 471578
rect 161572 471514 161624 471520
rect 162504 471209 162532 488022
rect 162964 476882 162992 488022
rect 163700 485489 163728 488022
rect 163792 488022 164082 488050
rect 164252 488022 164542 488050
rect 164620 488022 165002 488050
rect 165478 488022 165568 488050
rect 163686 485480 163742 485489
rect 163686 485415 163742 485424
rect 162952 476876 163004 476882
rect 162952 476818 163004 476824
rect 163792 476114 163820 488022
rect 162872 476086 163820 476114
rect 162490 471200 162546 471209
rect 162490 471135 162546 471144
rect 161478 468616 161534 468625
rect 161478 468551 161534 468560
rect 146300 467094 146352 467100
rect 153198 467120 153254 467129
rect 153198 467055 153254 467064
rect 142252 465860 142304 465866
rect 142252 465802 142304 465808
rect 162872 465769 162900 476086
rect 164252 469946 164280 488022
rect 164620 475454 164648 488022
rect 165540 483750 165568 488022
rect 165724 488022 165830 488050
rect 165528 483744 165580 483750
rect 165528 483686 165580 483692
rect 165724 476814 165752 488022
rect 166276 484838 166304 488036
rect 166368 488022 166750 488050
rect 167012 488022 167210 488050
rect 167288 488022 167670 488050
rect 167748 488022 168038 488050
rect 168392 488022 168498 488050
rect 168576 488022 168958 488050
rect 169036 488022 169418 488050
rect 169772 488022 169878 488050
rect 169956 488022 170246 488050
rect 170324 488022 170706 488050
rect 166264 484832 166316 484838
rect 166264 484774 166316 484780
rect 165712 476808 165764 476814
rect 165712 476750 165764 476756
rect 166368 476114 166396 488022
rect 165632 476086 166396 476114
rect 164608 475448 164660 475454
rect 164608 475390 164660 475396
rect 164240 469940 164292 469946
rect 164240 469882 164292 469888
rect 165632 466041 165660 476086
rect 165618 466032 165674 466041
rect 165618 465967 165674 465976
rect 167012 465905 167040 488022
rect 167092 484152 167144 484158
rect 167092 484094 167144 484100
rect 167104 468994 167132 484094
rect 167288 470594 167316 488022
rect 167748 484158 167776 488022
rect 167736 484152 167788 484158
rect 167736 484094 167788 484100
rect 167196 470566 167316 470594
rect 167092 468988 167144 468994
rect 167092 468930 167144 468936
rect 167196 468926 167224 470566
rect 167184 468920 167236 468926
rect 167184 468862 167236 468868
rect 168392 468489 168420 488022
rect 168576 484140 168604 488022
rect 168484 484112 168604 484140
rect 168484 468858 168512 484112
rect 169036 470594 169064 488022
rect 168576 470566 169064 470594
rect 168576 469062 168604 470566
rect 168564 469056 168616 469062
rect 168564 468998 168616 469004
rect 169772 468897 169800 488022
rect 169956 484140 169984 488022
rect 169864 484112 169984 484140
rect 169864 472841 169892 484112
rect 170324 478417 170352 488022
rect 171152 485625 171180 488036
rect 171244 488022 171626 488050
rect 171704 488022 171994 488050
rect 171138 485616 171194 485625
rect 171138 485551 171194 485560
rect 170404 485104 170456 485110
rect 170404 485046 170456 485052
rect 170310 478408 170366 478417
rect 170310 478343 170366 478352
rect 169850 472832 169906 472841
rect 169850 472767 169906 472776
rect 169758 468888 169814 468897
rect 168472 468852 168524 468858
rect 169758 468823 169814 468832
rect 168472 468794 168524 468800
rect 168378 468480 168434 468489
rect 168378 468415 168434 468424
rect 170416 466177 170444 485046
rect 171140 484152 171192 484158
rect 171140 484094 171192 484100
rect 171152 469033 171180 484094
rect 171244 471617 171272 488022
rect 171704 484158 171732 488022
rect 171692 484152 171744 484158
rect 171692 484094 171744 484100
rect 172440 481001 172468 488036
rect 172716 488022 172914 488050
rect 172992 488022 173374 488050
rect 173544 488022 173834 488050
rect 173912 488022 174202 488050
rect 174280 488022 174662 488050
rect 174832 488022 175122 488050
rect 175384 488022 175582 488050
rect 175752 488022 176042 488050
rect 176426 488022 176608 488050
rect 172520 484220 172572 484226
rect 172520 484162 172572 484168
rect 172426 480992 172482 481001
rect 172426 480927 172482 480936
rect 171230 471608 171286 471617
rect 171230 471543 171286 471552
rect 171138 469024 171194 469033
rect 171138 468959 171194 468968
rect 170402 466168 170458 466177
rect 170402 466103 170458 466112
rect 172532 466070 172560 484162
rect 172612 484152 172664 484158
rect 172612 484094 172664 484100
rect 172624 467265 172652 484094
rect 172716 471345 172744 488022
rect 172992 484158 173020 488022
rect 173544 484226 173572 488022
rect 173532 484220 173584 484226
rect 173532 484162 173584 484168
rect 172980 484152 173032 484158
rect 172980 484094 173032 484100
rect 172702 471336 172758 471345
rect 172702 471271 172758 471280
rect 172610 467256 172666 467265
rect 172610 467191 172666 467200
rect 173912 466206 173940 488022
rect 174280 484106 174308 488022
rect 174004 484078 174308 484106
rect 173900 466200 173952 466206
rect 173900 466142 173952 466148
rect 172520 466064 172572 466070
rect 172520 466006 172572 466012
rect 174004 465934 174032 484078
rect 174832 471753 174860 488022
rect 175280 484152 175332 484158
rect 175280 484094 175332 484100
rect 174818 471744 174874 471753
rect 174818 471679 174874 471688
rect 175292 467362 175320 484094
rect 175384 472734 175412 488022
rect 175752 484158 175780 488022
rect 175740 484152 175792 484158
rect 175740 484094 175792 484100
rect 176580 483818 176608 488022
rect 176764 488022 176870 488050
rect 177040 488022 177330 488050
rect 177408 488022 177790 488050
rect 178052 488022 178158 488050
rect 178236 488022 178618 488050
rect 178696 488022 179078 488050
rect 179554 488022 179644 488050
rect 176568 483812 176620 483818
rect 176568 483754 176620 483760
rect 176660 480888 176712 480894
rect 176660 480830 176712 480836
rect 176672 474366 176700 480830
rect 176764 475522 176792 488022
rect 177040 478242 177068 488022
rect 177408 480894 177436 488022
rect 177396 480888 177448 480894
rect 177396 480830 177448 480836
rect 177028 478236 177080 478242
rect 177028 478178 177080 478184
rect 176752 475516 176804 475522
rect 176752 475458 176804 475464
rect 176660 474360 176712 474366
rect 176660 474302 176712 474308
rect 175372 472728 175424 472734
rect 175372 472670 175424 472676
rect 178052 469130 178080 488022
rect 178236 476114 178264 488022
rect 178696 479777 178724 488022
rect 179616 481098 179644 488022
rect 179708 488022 179998 488050
rect 180076 488022 180366 488050
rect 180842 488022 180932 488050
rect 179604 481092 179656 481098
rect 179604 481034 179656 481040
rect 179708 480842 179736 488022
rect 179788 481092 179840 481098
rect 179788 481034 179840 481040
rect 179432 480814 179736 480842
rect 178682 479768 178738 479777
rect 178682 479703 178738 479712
rect 178144 476086 178264 476114
rect 178144 470082 178172 476086
rect 178132 470076 178184 470082
rect 178132 470018 178184 470024
rect 178040 469124 178092 469130
rect 178040 469066 178092 469072
rect 178040 467832 178092 467838
rect 178040 467774 178092 467780
rect 175280 467356 175332 467362
rect 175280 467298 175332 467304
rect 178052 466614 178080 467774
rect 178040 466608 178092 466614
rect 178038 466576 178040 466585
rect 178092 466576 178094 466585
rect 178038 466511 178094 466520
rect 179432 466002 179460 480814
rect 179512 480752 179564 480758
rect 179512 480694 179564 480700
rect 179524 470014 179552 480694
rect 179800 474298 179828 481034
rect 180076 480758 180104 488022
rect 180800 480888 180852 480894
rect 180800 480830 180852 480836
rect 180064 480752 180116 480758
rect 180064 480694 180116 480700
rect 179788 474292 179840 474298
rect 179788 474234 179840 474240
rect 180156 474020 180208 474026
rect 180156 473962 180208 473968
rect 179512 470008 179564 470014
rect 179512 469950 179564 469956
rect 180168 467294 180196 473962
rect 180156 467288 180208 467294
rect 180156 467230 180208 467236
rect 180168 466993 180196 467230
rect 180154 466984 180210 466993
rect 180154 466919 180210 466928
rect 179420 465996 179472 466002
rect 179420 465938 179472 465944
rect 173992 465928 174044 465934
rect 166998 465896 167054 465905
rect 173992 465870 174044 465876
rect 166998 465831 167054 465840
rect 162858 465760 162914 465769
rect 162858 465695 162914 465704
rect 180812 464642 180840 480830
rect 180904 466138 180932 488022
rect 180996 488022 181286 488050
rect 181456 488022 181746 488050
rect 182222 488022 182404 488050
rect 180996 466342 181024 488022
rect 181456 480894 181484 488022
rect 182376 481098 182404 488022
rect 182468 488022 182574 488050
rect 182744 488022 183034 488050
rect 183112 488022 183494 488050
rect 183756 488022 183954 488050
rect 184032 488022 184322 488050
rect 184400 488022 184782 488050
rect 184952 488022 185242 488050
rect 182364 481092 182416 481098
rect 182364 481034 182416 481040
rect 181444 480888 181496 480894
rect 181444 480830 181496 480836
rect 182180 480888 182232 480894
rect 182180 480830 182232 480836
rect 182192 467430 182220 480830
rect 182468 478224 182496 488022
rect 182548 481092 182600 481098
rect 182548 481034 182600 481040
rect 182284 478196 182496 478224
rect 182284 471481 182312 478196
rect 182560 473354 182588 481034
rect 182744 480894 182772 488022
rect 182732 480888 182784 480894
rect 182732 480830 182784 480836
rect 182376 473326 182588 473354
rect 182270 471472 182326 471481
rect 182270 471407 182326 471416
rect 182376 471170 182404 473326
rect 183112 471918 183140 488022
rect 183560 480888 183612 480894
rect 183560 480830 183612 480836
rect 183100 471912 183152 471918
rect 183100 471854 183152 471860
rect 183572 471238 183600 480830
rect 183652 477692 183704 477698
rect 183652 477634 183704 477640
rect 183664 471646 183692 477634
rect 183652 471640 183704 471646
rect 183652 471582 183704 471588
rect 183560 471232 183612 471238
rect 183560 471174 183612 471180
rect 182364 471164 182416 471170
rect 182364 471106 182416 471112
rect 183756 471102 183784 488022
rect 184032 477698 184060 488022
rect 184400 480894 184428 488022
rect 184388 480888 184440 480894
rect 184388 480830 184440 480836
rect 184020 477692 184072 477698
rect 184020 477634 184072 477640
rect 184952 472666 184980 488022
rect 185584 484968 185636 484974
rect 185688 484945 185716 488036
rect 185872 488022 186162 488050
rect 186424 488022 186530 488050
rect 187006 488022 187096 488050
rect 185584 484910 185636 484916
rect 185674 484936 185730 484945
rect 185032 477692 185084 477698
rect 185032 477634 185084 477640
rect 185044 475590 185072 477634
rect 185032 475584 185084 475590
rect 185032 475526 185084 475532
rect 184940 472660 184992 472666
rect 184940 472602 184992 472608
rect 183744 471096 183796 471102
rect 183744 471038 183796 471044
rect 182180 467424 182232 467430
rect 182180 467366 182232 467372
rect 180984 466336 181036 466342
rect 180984 466278 181036 466284
rect 180892 466132 180944 466138
rect 180892 466074 180944 466080
rect 185596 464778 185624 484910
rect 185674 484871 185730 484880
rect 185872 477698 185900 488022
rect 186320 484152 186372 484158
rect 186320 484094 186372 484100
rect 185860 477692 185912 477698
rect 185860 477634 185912 477640
rect 186332 465662 186360 484094
rect 186424 474026 186452 488022
rect 187068 485761 187096 488022
rect 187160 488022 187450 488050
rect 187712 488022 187910 488050
rect 188080 488022 188370 488050
rect 188448 488022 188738 488050
rect 189214 488022 189304 488050
rect 187054 485752 187110 485761
rect 187054 485687 187110 485696
rect 187160 484158 187188 488022
rect 187148 484152 187200 484158
rect 187148 484094 187200 484100
rect 186412 474020 186464 474026
rect 186412 473962 186464 473968
rect 186320 465656 186372 465662
rect 186320 465598 186372 465604
rect 185584 464772 185636 464778
rect 185584 464714 185636 464720
rect 180800 464636 180852 464642
rect 180800 464578 180852 464584
rect 142160 464568 142212 464574
rect 142160 464510 142212 464516
rect 138020 464432 138072 464438
rect 187712 464409 187740 488022
rect 187792 484152 187844 484158
rect 187792 484094 187844 484100
rect 187804 465594 187832 484094
rect 188080 472802 188108 488022
rect 188448 484158 188476 488022
rect 188436 484152 188488 484158
rect 188436 484094 188488 484100
rect 189080 483404 189132 483410
rect 189080 483346 189132 483352
rect 188068 472796 188120 472802
rect 188068 472738 188120 472744
rect 189092 466274 189120 483346
rect 189172 481772 189224 481778
rect 189172 481714 189224 481720
rect 189184 468314 189212 481714
rect 189276 479670 189304 488022
rect 189368 488022 189658 488050
rect 189736 488022 190118 488050
rect 190502 488022 190592 488050
rect 189368 483410 189396 488022
rect 189356 483404 189408 483410
rect 189356 483346 189408 483352
rect 189736 481778 189764 488022
rect 190460 484152 190512 484158
rect 190460 484094 190512 484100
rect 189724 481772 189776 481778
rect 189724 481714 189776 481720
rect 189264 479664 189316 479670
rect 189264 479606 189316 479612
rect 189172 468308 189224 468314
rect 189172 468250 189224 468256
rect 189080 466268 189132 466274
rect 189080 466210 189132 466216
rect 187792 465588 187844 465594
rect 187792 465530 187844 465536
rect 190472 464846 190500 484094
rect 190564 471714 190592 488022
rect 190656 488022 190946 488050
rect 191024 488022 191406 488050
rect 191882 488022 192064 488050
rect 190656 471782 190684 488022
rect 191024 484158 191052 488022
rect 191840 484220 191892 484226
rect 191840 484162 191892 484168
rect 191012 484152 191064 484158
rect 191012 484094 191064 484100
rect 190644 471776 190696 471782
rect 190644 471718 190696 471724
rect 190552 471708 190604 471714
rect 190552 471650 190604 471656
rect 191852 468382 191880 484162
rect 191932 484152 191984 484158
rect 191932 484094 191984 484100
rect 191944 468450 191972 484094
rect 192036 471850 192064 488022
rect 192128 488022 192326 488050
rect 192404 488022 192694 488050
rect 192772 488022 193154 488050
rect 193416 488022 193614 488050
rect 193784 488022 194074 488050
rect 194152 488022 194534 488050
rect 194918 488022 195192 488050
rect 192128 484158 192156 488022
rect 192404 484226 192432 488022
rect 192392 484220 192444 484226
rect 192392 484162 192444 484168
rect 192116 484152 192168 484158
rect 192116 484094 192168 484100
rect 192772 471986 192800 488022
rect 193220 484220 193272 484226
rect 193220 484162 193272 484168
rect 192760 471980 192812 471986
rect 192760 471922 192812 471928
rect 192024 471844 192076 471850
rect 192024 471786 192076 471792
rect 191932 468444 191984 468450
rect 191932 468386 191984 468392
rect 191840 468376 191892 468382
rect 191840 468318 191892 468324
rect 190918 466576 190974 466585
rect 190918 466511 190974 466520
rect 190932 466478 190960 466511
rect 190920 466472 190972 466478
rect 190920 466414 190972 466420
rect 190460 464840 190512 464846
rect 190460 464782 190512 464788
rect 193232 464710 193260 484162
rect 193312 484152 193364 484158
rect 193312 484094 193364 484100
rect 193324 466410 193352 484094
rect 193416 469198 193444 488022
rect 193784 484158 193812 488022
rect 194152 484226 194180 488022
rect 195164 484430 195192 488022
rect 195348 484974 195376 488036
rect 195440 488022 195822 488050
rect 196298 488022 196664 488050
rect 195336 484968 195388 484974
rect 195336 484910 195388 484916
rect 195152 484424 195204 484430
rect 195152 484366 195204 484372
rect 194140 484220 194192 484226
rect 194140 484162 194192 484168
rect 193772 484152 193824 484158
rect 193772 484094 193824 484100
rect 195440 470594 195468 488022
rect 194612 470566 195468 470594
rect 193404 469192 193456 469198
rect 193404 469134 193456 469140
rect 193312 466404 193364 466410
rect 193312 466346 193364 466352
rect 194612 465526 194640 470566
rect 194600 465520 194652 465526
rect 194600 465462 194652 465468
rect 193220 464704 193272 464710
rect 193220 464646 193272 464652
rect 138020 464374 138072 464380
rect 187698 464400 187754 464409
rect 132500 464364 132552 464370
rect 132500 464306 132552 464312
rect 136640 464364 136692 464370
rect 187698 464335 187754 464344
rect 136640 464306 136692 464312
rect 195888 380996 195940 381002
rect 195888 380938 195940 380944
rect 60740 380928 60792 380934
rect 60740 380870 60792 380876
rect 60752 357406 60780 380870
rect 110970 380760 111026 380769
rect 110970 380695 111026 380704
rect 113546 380760 113602 380769
rect 113546 380695 113602 380704
rect 116030 380760 116086 380769
rect 116030 380695 116086 380704
rect 118422 380760 118478 380769
rect 118422 380695 118478 380704
rect 120998 380760 121054 380769
rect 120998 380695 121054 380704
rect 123482 380760 123538 380769
rect 123482 380695 123538 380704
rect 125966 380760 126022 380769
rect 125966 380695 126022 380704
rect 131026 380760 131082 380769
rect 131026 380695 131082 380704
rect 133510 380760 133566 380769
rect 133510 380695 133566 380704
rect 140962 380760 141018 380769
rect 140962 380695 141018 380704
rect 143538 380760 143594 380769
rect 143538 380695 143594 380704
rect 146022 380760 146078 380769
rect 146022 380695 146078 380704
rect 155958 380760 156014 380769
rect 155958 380695 155960 380704
rect 110984 380390 111012 380695
rect 113560 380526 113588 380695
rect 113548 380520 113600 380526
rect 113548 380462 113600 380468
rect 110972 380384 111024 380390
rect 110972 380326 111024 380332
rect 116044 380186 116072 380695
rect 118436 380458 118464 380695
rect 118424 380452 118476 380458
rect 118424 380394 118476 380400
rect 121012 380186 121040 380695
rect 123496 380322 123524 380695
rect 123484 380316 123536 380322
rect 123484 380258 123536 380264
rect 125980 380254 126008 380695
rect 131040 380322 131068 380695
rect 133524 380390 133552 380695
rect 140976 380594 141004 380695
rect 140964 380588 141016 380594
rect 140964 380530 141016 380536
rect 143552 380458 143580 380695
rect 146036 380526 146064 380695
rect 156012 380695 156014 380704
rect 158534 380760 158590 380769
rect 158534 380695 158590 380704
rect 160926 380760 160982 380769
rect 160926 380695 160982 380704
rect 163410 380760 163466 380769
rect 163410 380695 163466 380704
rect 165986 380760 166042 380769
rect 165986 380695 166042 380704
rect 155960 380666 156012 380672
rect 158548 380662 158576 380695
rect 158536 380656 158588 380662
rect 158536 380598 158588 380604
rect 146024 380520 146076 380526
rect 146024 380462 146076 380468
rect 143540 380452 143592 380458
rect 143540 380394 143592 380400
rect 133512 380384 133564 380390
rect 133512 380326 133564 380332
rect 131028 380316 131080 380322
rect 131028 380258 131080 380264
rect 125968 380248 126020 380254
rect 128360 380248 128412 380254
rect 125968 380190 126020 380196
rect 128358 380216 128360 380225
rect 128412 380216 128414 380225
rect 116032 380180 116084 380186
rect 116032 380122 116084 380128
rect 121000 380180 121052 380186
rect 128358 380151 128414 380160
rect 121000 380122 121052 380128
rect 160940 380118 160968 380695
rect 160928 380112 160980 380118
rect 160928 380054 160980 380060
rect 163424 380050 163452 380695
rect 163412 380044 163464 380050
rect 163412 379986 163464 379992
rect 166000 379982 166028 380695
rect 165988 379976 166040 379982
rect 165988 379918 166040 379924
rect 86592 379500 86644 379506
rect 86592 379442 86644 379448
rect 86604 379409 86632 379442
rect 88340 379432 88392 379438
rect 85486 379400 85542 379409
rect 85486 379335 85542 379344
rect 86590 379400 86646 379409
rect 86590 379335 86646 379344
rect 87878 379400 87934 379409
rect 87878 379335 87934 379344
rect 88338 379400 88340 379409
rect 92388 379432 92440 379438
rect 88392 379400 88394 379409
rect 88338 379335 88394 379344
rect 88798 379400 88854 379409
rect 88798 379335 88800 379344
rect 80426 379264 80482 379273
rect 80426 379199 80482 379208
rect 77206 378992 77262 379001
rect 77206 378927 77262 378936
rect 77220 376718 77248 378927
rect 80440 378321 80468 379199
rect 83278 378856 83334 378865
rect 83278 378791 83334 378800
rect 80426 378312 80482 378321
rect 80426 378247 80482 378256
rect 80440 378214 80468 378247
rect 80428 378208 80480 378214
rect 80428 378150 80480 378156
rect 77208 376712 77260 376718
rect 77208 376654 77260 376660
rect 83292 376446 83320 378791
rect 85500 378282 85528 379335
rect 85488 378276 85540 378282
rect 85488 378218 85540 378224
rect 87892 378214 87920 379335
rect 88852 379335 88854 379344
rect 90086 379400 90142 379409
rect 90086 379335 90142 379344
rect 90638 379400 90694 379409
rect 90638 379335 90694 379344
rect 91374 379400 91430 379409
rect 91374 379335 91430 379344
rect 92386 379400 92388 379409
rect 92440 379400 92442 379409
rect 92386 379335 92442 379344
rect 93582 379400 93638 379409
rect 93582 379335 93638 379344
rect 96066 379400 96122 379409
rect 96066 379335 96122 379344
rect 98274 379400 98330 379409
rect 98274 379335 98330 379344
rect 98458 379400 98514 379409
rect 98458 379335 98514 379344
rect 101034 379400 101090 379409
rect 101034 379335 101090 379344
rect 103518 379400 103574 379409
rect 103518 379335 103574 379344
rect 104898 379400 104954 379409
rect 104898 379335 104954 379344
rect 108210 379400 108266 379409
rect 108210 379335 108266 379344
rect 108854 379400 108910 379409
rect 108854 379335 108910 379344
rect 111338 379400 111394 379409
rect 111338 379335 111394 379344
rect 112350 379400 112406 379409
rect 112350 379335 112406 379344
rect 113454 379400 113510 379409
rect 113454 379335 113510 379344
rect 114466 379400 114522 379409
rect 114466 379335 114522 379344
rect 115846 379400 115902 379409
rect 115846 379335 115902 379344
rect 135902 379400 135958 379409
rect 135902 379335 135958 379344
rect 138478 379400 138534 379409
rect 138478 379335 138534 379344
rect 150990 379400 151046 379409
rect 150990 379335 151046 379344
rect 154026 379400 154082 379409
rect 154026 379335 154082 379344
rect 88800 379306 88852 379312
rect 90100 378350 90128 379335
rect 90652 379302 90680 379335
rect 90640 379296 90692 379302
rect 90640 379238 90692 379244
rect 91388 379234 91416 379335
rect 93490 379264 93546 379273
rect 91376 379228 91428 379234
rect 93490 379199 93546 379208
rect 91376 379170 91428 379176
rect 93504 379166 93532 379199
rect 93596 379166 93624 379335
rect 95974 379264 96030 379273
rect 95974 379199 96030 379208
rect 93492 379160 93544 379166
rect 93492 379102 93544 379108
rect 93584 379160 93636 379166
rect 93584 379102 93636 379108
rect 94686 378992 94742 379001
rect 94686 378927 94742 378936
rect 90088 378344 90140 378350
rect 90088 378286 90140 378292
rect 87880 378208 87932 378214
rect 84382 378176 84438 378185
rect 87880 378150 87932 378156
rect 84382 378111 84438 378120
rect 83280 376440 83332 376446
rect 83280 376382 83332 376388
rect 84396 375358 84424 378111
rect 94700 376514 94728 378927
rect 95988 377806 96016 379199
rect 96080 378690 96108 379335
rect 96068 378684 96120 378690
rect 96068 378626 96120 378632
rect 97814 378584 97870 378593
rect 97814 378519 97870 378528
rect 95976 377800 96028 377806
rect 95976 377742 96028 377748
rect 94688 376508 94740 376514
rect 94688 376450 94740 376456
rect 97828 376038 97856 378519
rect 98288 377738 98316 379335
rect 98472 378758 98500 379335
rect 99470 379264 99526 379273
rect 99470 379199 99526 379208
rect 98460 378752 98512 378758
rect 98460 378694 98512 378700
rect 98276 377732 98328 377738
rect 98276 377674 98328 377680
rect 99484 376378 99512 379199
rect 101048 379030 101076 379335
rect 102966 379264 103022 379273
rect 102966 379199 103022 379208
rect 101036 379024 101088 379030
rect 101036 378966 101088 378972
rect 100850 378584 100906 378593
rect 100850 378519 100906 378528
rect 99472 376372 99524 376378
rect 99472 376314 99524 376320
rect 97816 376032 97868 376038
rect 97816 375974 97868 375980
rect 100864 375902 100892 378519
rect 101862 378176 101918 378185
rect 101862 378111 101918 378120
rect 100852 375896 100904 375902
rect 100852 375838 100904 375844
rect 84384 375352 84436 375358
rect 84384 375294 84436 375300
rect 101876 375222 101904 378111
rect 102980 375290 103008 379199
rect 103532 378962 103560 379335
rect 103520 378956 103572 378962
rect 103520 378898 103572 378904
rect 104912 378894 104940 379335
rect 108224 379098 108252 379335
rect 108868 379098 108896 379335
rect 108212 379092 108264 379098
rect 108212 379034 108264 379040
rect 108856 379092 108908 379098
rect 108856 379034 108908 379040
rect 104900 378888 104952 378894
rect 104900 378830 104952 378836
rect 105726 378448 105782 378457
rect 111352 378418 111380 379335
rect 112364 379030 112392 379335
rect 112352 379024 112404 379030
rect 112352 378966 112404 378972
rect 113468 378622 113496 379335
rect 113456 378616 113508 378622
rect 113456 378558 113508 378564
rect 114480 378554 114508 379335
rect 114468 378548 114520 378554
rect 114468 378490 114520 378496
rect 115860 378486 115888 379335
rect 115848 378480 115900 378486
rect 115848 378422 115900 378428
rect 105726 378383 105782 378392
rect 111340 378412 111392 378418
rect 105740 375698 105768 378383
rect 111340 378354 111392 378360
rect 106462 378176 106518 378185
rect 106462 378111 106518 378120
rect 107566 378176 107622 378185
rect 107566 378111 107622 378120
rect 105728 375692 105780 375698
rect 105728 375634 105780 375640
rect 102968 375284 103020 375290
rect 102968 375226 103020 375232
rect 101864 375216 101916 375222
rect 101864 375158 101916 375164
rect 106476 375086 106504 378111
rect 107580 375154 107608 378111
rect 135916 376582 135944 379335
rect 138492 377330 138520 379335
rect 148690 378992 148746 379001
rect 148690 378927 148746 378936
rect 138480 377324 138532 377330
rect 138480 377266 138532 377272
rect 135904 376576 135956 376582
rect 135904 376518 135956 376524
rect 148704 376310 148732 378927
rect 151004 377398 151032 379335
rect 150992 377392 151044 377398
rect 150992 377334 151044 377340
rect 154040 377194 154068 379335
rect 183466 378992 183522 379001
rect 183466 378927 183522 378936
rect 182270 378448 182326 378457
rect 182270 378383 182326 378392
rect 182284 377874 182312 378383
rect 183480 377942 183508 378927
rect 183468 377936 183520 377942
rect 183468 377878 183520 377884
rect 182272 377868 182324 377874
rect 182272 377810 182324 377816
rect 182824 377868 182876 377874
rect 182824 377810 182876 377816
rect 154028 377188 154080 377194
rect 154028 377130 154080 377136
rect 148692 376304 148744 376310
rect 148692 376246 148744 376252
rect 107568 375148 107620 375154
rect 107568 375090 107620 375096
rect 106464 375080 106516 375086
rect 106464 375022 106516 375028
rect 180156 360188 180208 360194
rect 180156 360130 180208 360136
rect 180168 358873 180196 360130
rect 178590 358864 178646 358873
rect 178590 358799 178592 358808
rect 178644 358799 178646 358808
rect 180154 358864 180210 358873
rect 180154 358799 180210 358808
rect 178592 358770 178644 358776
rect 182836 358086 182864 377810
rect 183480 374678 183508 377878
rect 183468 374672 183520 374678
rect 183468 374614 183520 374620
rect 195900 360194 195928 380938
rect 196636 377602 196664 488022
rect 196728 378146 196756 488036
rect 196820 488022 197110 488050
rect 196716 378140 196768 378146
rect 196716 378082 196768 378088
rect 196820 377670 196848 488022
rect 197452 485376 197504 485382
rect 197452 485318 197504 485324
rect 197360 485172 197412 485178
rect 197360 485114 197412 485120
rect 197372 484945 197400 485114
rect 197358 484936 197414 484945
rect 197358 484871 197414 484880
rect 197464 484809 197492 485318
rect 197450 484800 197506 484809
rect 197450 484735 197506 484744
rect 197084 484424 197136 484430
rect 197084 484366 197136 484372
rect 196900 471300 196952 471306
rect 196900 471242 196952 471248
rect 196808 377664 196860 377670
rect 196808 377606 196860 377612
rect 196624 377596 196676 377602
rect 196624 377538 196676 377544
rect 195888 360188 195940 360194
rect 195888 360130 195940 360136
rect 195900 359718 195928 360130
rect 195888 359712 195940 359718
rect 195888 359654 195940 359660
rect 190920 359508 190972 359514
rect 190920 359450 190972 359456
rect 190932 358873 190960 359450
rect 190918 358864 190974 358873
rect 190918 358799 190974 358808
rect 182824 358080 182876 358086
rect 182824 358022 182876 358028
rect 60740 357400 60792 357406
rect 60740 357342 60792 357348
rect 196912 277394 196940 471242
rect 196992 468784 197044 468790
rect 196992 468726 197044 468732
rect 197004 376310 197032 468726
rect 197096 377534 197124 484366
rect 197452 484152 197504 484158
rect 197452 484094 197504 484100
rect 197176 382220 197228 382226
rect 197176 382162 197228 382168
rect 197084 377528 197136 377534
rect 197084 377470 197136 377476
rect 196992 376304 197044 376310
rect 196992 376246 197044 376252
rect 196636 277366 196940 277394
rect 113362 273864 113418 273873
rect 113362 273799 113418 273808
rect 61566 273320 61622 273329
rect 61566 273255 61622 273264
rect 61106 273048 61162 273057
rect 61106 272983 61162 272992
rect 61016 272944 61068 272950
rect 61016 272886 61068 272892
rect 60922 272640 60978 272649
rect 60922 272575 60978 272584
rect 60738 272504 60794 272513
rect 60738 272439 60794 272448
rect 60752 252521 60780 272439
rect 60832 272332 60884 272338
rect 60832 272274 60884 272280
rect 60844 271930 60872 272274
rect 60832 271924 60884 271930
rect 60832 271866 60884 271872
rect 60738 252512 60794 252521
rect 60738 252447 60794 252456
rect 60844 252142 60872 271866
rect 60832 252136 60884 252142
rect 60832 252078 60884 252084
rect 60936 252006 60964 272575
rect 60924 252000 60976 252006
rect 60924 251942 60976 251948
rect 61028 251802 61056 272886
rect 61120 271561 61148 272983
rect 61476 272944 61528 272950
rect 61474 272912 61476 272921
rect 61528 272912 61530 272921
rect 61474 272847 61530 272856
rect 61106 271552 61162 271561
rect 61106 271487 61162 271496
rect 61120 251938 61148 271487
rect 61580 271153 61608 273255
rect 76010 273184 76066 273193
rect 76010 273119 76066 273128
rect 77114 273184 77170 273193
rect 77114 273119 77170 273128
rect 83002 273184 83058 273193
rect 83002 273119 83058 273128
rect 90730 273184 90786 273193
rect 90730 273119 90786 273128
rect 93674 273184 93730 273193
rect 93674 273119 93730 273128
rect 95882 273184 95938 273193
rect 96066 273184 96122 273193
rect 95882 273119 95938 273128
rect 95988 273142 96066 273170
rect 76024 272406 76052 273119
rect 77128 272474 77156 273119
rect 83016 273018 83044 273119
rect 83004 273012 83056 273018
rect 83004 272954 83056 272960
rect 90744 272746 90772 273119
rect 90732 272740 90784 272746
rect 90732 272682 90784 272688
rect 93688 272678 93716 273119
rect 95896 273086 95924 273119
rect 95884 273080 95936 273086
rect 95884 273022 95936 273028
rect 95882 272776 95938 272785
rect 95988 272762 96016 273142
rect 96066 273119 96122 273128
rect 95938 272734 96016 272762
rect 96066 272776 96122 272785
rect 95882 272711 95938 272720
rect 96066 272711 96122 272720
rect 98458 272776 98514 272785
rect 98458 272711 98514 272720
rect 93676 272672 93728 272678
rect 93676 272614 93728 272620
rect 96080 272610 96108 272711
rect 96068 272604 96120 272610
rect 96068 272546 96120 272552
rect 98472 272542 98500 272711
rect 98460 272536 98512 272542
rect 98460 272478 98512 272484
rect 77116 272468 77168 272474
rect 77116 272410 77168 272416
rect 98092 272468 98144 272474
rect 98092 272410 98144 272416
rect 76012 272400 76064 272406
rect 76012 272342 76064 272348
rect 87602 272368 87658 272377
rect 62212 272332 62264 272338
rect 87602 272303 87658 272312
rect 94410 272368 94466 272377
rect 94410 272303 94412 272312
rect 62212 272274 62264 272280
rect 61566 271144 61622 271153
rect 61566 271079 61622 271088
rect 62118 271144 62174 271153
rect 62118 271079 62174 271088
rect 61108 251932 61160 251938
rect 61108 251874 61160 251880
rect 61016 251796 61068 251802
rect 61016 251738 61068 251744
rect 62132 251394 62160 271079
rect 62224 270609 62252 272274
rect 87616 272270 87644 272303
rect 94464 272303 94466 272312
rect 94412 272274 94464 272280
rect 87604 272264 87656 272270
rect 87604 272206 87656 272212
rect 96620 272060 96672 272066
rect 96620 272002 96672 272008
rect 85764 271992 85816 271998
rect 85764 271934 85816 271940
rect 84198 271824 84254 271833
rect 84198 271759 84254 271768
rect 77298 271008 77354 271017
rect 77298 270943 77300 270952
rect 77352 270943 77354 270952
rect 77300 270914 77352 270920
rect 62210 270600 62266 270609
rect 62210 270535 62266 270544
rect 84212 270434 84240 271759
rect 84658 271688 84714 271697
rect 84658 271623 84714 271632
rect 84200 270428 84252 270434
rect 84200 270370 84252 270376
rect 81440 270360 81492 270366
rect 81440 270302 81492 270308
rect 80060 270292 80112 270298
rect 80060 270234 80112 270240
rect 63500 270224 63552 270230
rect 63500 270166 63552 270172
rect 63512 268666 63540 270166
rect 77392 270020 77444 270026
rect 77392 269962 77444 269968
rect 63500 268660 63552 268666
rect 63500 268602 63552 268608
rect 77404 268569 77432 269962
rect 80072 268598 80100 270234
rect 80060 268592 80112 268598
rect 77390 268560 77446 268569
rect 80060 268534 80112 268540
rect 81452 268530 81480 270302
rect 84672 270162 84700 271623
rect 85578 270600 85634 270609
rect 85578 270535 85634 270544
rect 84660 270156 84712 270162
rect 84660 270098 84712 270104
rect 85592 269822 85620 270535
rect 85580 269816 85632 269822
rect 85580 269758 85632 269764
rect 77390 268495 77446 268504
rect 81440 268524 81492 268530
rect 81440 268466 81492 268472
rect 85776 268433 85804 271934
rect 96632 271833 96660 272002
rect 96618 271824 96674 271833
rect 96618 271759 96674 271768
rect 98104 271697 98132 272410
rect 99378 272232 99434 272241
rect 99378 272167 99380 272176
rect 99432 272167 99434 272176
rect 99380 272138 99432 272144
rect 100760 272128 100812 272134
rect 100760 272070 100812 272076
rect 100772 271833 100800 272070
rect 106556 271992 106608 271998
rect 106556 271934 106608 271940
rect 106280 271924 106332 271930
rect 106280 271866 106332 271872
rect 106292 271833 106320 271866
rect 106568 271833 106596 271934
rect 112352 271924 112404 271930
rect 112352 271866 112404 271872
rect 112364 271833 112392 271866
rect 100758 271824 100814 271833
rect 100758 271759 100814 271768
rect 106278 271824 106334 271833
rect 106278 271759 106334 271768
rect 106554 271824 106610 271833
rect 106554 271759 106610 271768
rect 112350 271824 112406 271833
rect 112350 271759 112406 271768
rect 98090 271688 98146 271697
rect 98090 271623 98146 271632
rect 107658 271688 107714 271697
rect 107658 271623 107714 271632
rect 88338 271280 88394 271289
rect 88338 271215 88394 271224
rect 88352 271046 88380 271215
rect 88340 271040 88392 271046
rect 88340 270982 88392 270988
rect 88338 270872 88394 270881
rect 88338 270807 88394 270816
rect 88352 269958 88380 270807
rect 89718 270736 89774 270745
rect 89718 270671 89774 270680
rect 92478 270736 92534 270745
rect 92478 270671 92534 270680
rect 88340 269952 88392 269958
rect 88340 269894 88392 269900
rect 89732 269890 89760 270671
rect 91098 270600 91154 270609
rect 91098 270535 91154 270544
rect 91112 270094 91140 270535
rect 92492 270230 92520 270671
rect 92480 270224 92532 270230
rect 92480 270166 92532 270172
rect 91100 270088 91152 270094
rect 91100 270030 91152 270036
rect 89720 269884 89772 269890
rect 89720 269826 89772 269832
rect 85762 268424 85818 268433
rect 98104 268394 98132 271623
rect 100758 271552 100814 271561
rect 100758 271487 100814 271496
rect 100772 271114 100800 271487
rect 104898 271416 104954 271425
rect 104898 271351 104954 271360
rect 103518 271280 103574 271289
rect 104912 271250 104940 271351
rect 103518 271215 103574 271224
rect 104900 271244 104952 271250
rect 103532 271182 103560 271215
rect 104900 271186 104952 271192
rect 103520 271176 103572 271182
rect 103520 271118 103572 271124
rect 107672 271114 107700 271623
rect 109222 271416 109278 271425
rect 109222 271351 109278 271360
rect 113270 271416 113326 271425
rect 113270 271351 113326 271360
rect 100760 271108 100812 271114
rect 100760 271050 100812 271056
rect 107660 271108 107712 271114
rect 107660 271050 107712 271056
rect 106924 271040 106976 271046
rect 106924 270982 106976 270988
rect 104898 270736 104954 270745
rect 104898 270671 104954 270680
rect 104912 268462 104940 270671
rect 104900 268456 104952 268462
rect 104900 268398 104952 268404
rect 85762 268359 85818 268368
rect 98092 268388 98144 268394
rect 98092 268330 98144 268336
rect 106936 251870 106964 270982
rect 107658 270600 107714 270609
rect 107658 270535 107714 270544
rect 107672 270366 107700 270535
rect 107660 270360 107712 270366
rect 107660 270302 107712 270308
rect 109236 270298 109264 271351
rect 110418 271280 110474 271289
rect 110418 271215 110474 271224
rect 113178 271280 113234 271289
rect 113178 271215 113180 271224
rect 110432 271182 110460 271215
rect 113232 271215 113234 271224
rect 113180 271186 113232 271192
rect 110420 271176 110472 271182
rect 110420 271118 110472 271124
rect 113284 271046 113312 271351
rect 113272 271040 113324 271046
rect 113272 270982 113324 270988
rect 110418 270600 110474 270609
rect 110418 270535 110474 270544
rect 109224 270292 109276 270298
rect 109224 270234 109276 270240
rect 110432 270026 110460 270535
rect 110420 270020 110472 270026
rect 110420 269962 110472 269968
rect 113376 269822 113404 273799
rect 133418 273728 133474 273737
rect 133418 273663 133474 273672
rect 133432 273630 133460 273663
rect 133420 273624 133472 273630
rect 133420 273566 133472 273572
rect 135902 273592 135958 273601
rect 135902 273527 135904 273536
rect 135956 273527 135958 273536
rect 138478 273592 138534 273601
rect 138478 273527 138534 273536
rect 140870 273592 140926 273601
rect 140870 273527 140926 273536
rect 143538 273592 143594 273601
rect 143538 273527 143594 273536
rect 145930 273592 145986 273601
rect 145930 273527 145986 273536
rect 135904 273498 135956 273504
rect 138492 273494 138520 273527
rect 138480 273488 138532 273494
rect 138480 273430 138532 273436
rect 140884 273426 140912 273527
rect 140872 273420 140924 273426
rect 140872 273362 140924 273368
rect 143552 273358 143580 273527
rect 143540 273352 143592 273358
rect 143540 273294 143592 273300
rect 145944 273290 145972 273527
rect 145932 273284 145984 273290
rect 145932 273226 145984 273232
rect 196636 271930 196664 277366
rect 197188 272542 197216 382162
rect 197464 378010 197492 484094
rect 197452 378004 197504 378010
rect 197452 377946 197504 377952
rect 197556 377874 197584 488036
rect 197648 488022 198030 488050
rect 198200 488022 198490 488050
rect 198874 488022 199240 488050
rect 199334 488022 199424 488050
rect 197648 377942 197676 488022
rect 197912 486668 197964 486674
rect 197912 486610 197964 486616
rect 197728 468648 197780 468654
rect 197728 468590 197780 468596
rect 197636 377936 197688 377942
rect 197636 377878 197688 377884
rect 197544 377868 197596 377874
rect 197544 377810 197596 377816
rect 197636 374672 197688 374678
rect 197636 374614 197688 374620
rect 197544 359712 197596 359718
rect 197544 359654 197596 359660
rect 197360 359576 197412 359582
rect 197360 359518 197412 359524
rect 197372 358834 197400 359518
rect 197360 358828 197412 358834
rect 197360 358770 197412 358776
rect 197372 354674 197400 358770
rect 197372 354646 197492 354674
rect 197176 272536 197228 272542
rect 197176 272478 197228 272484
rect 196624 271924 196676 271930
rect 196624 271866 196676 271872
rect 123116 271856 123168 271862
rect 123114 271824 123116 271833
rect 154488 271856 154540 271862
rect 123168 271824 123170 271833
rect 123114 271759 123170 271768
rect 125598 271824 125654 271833
rect 125598 271759 125654 271768
rect 128358 271824 128414 271833
rect 128358 271759 128360 271768
rect 125612 271726 125640 271759
rect 128412 271759 128414 271768
rect 151358 271824 151414 271833
rect 151358 271759 151360 271768
rect 128360 271730 128412 271736
rect 151412 271759 151414 271768
rect 154486 271824 154488 271833
rect 154540 271824 154542 271833
rect 154486 271759 154542 271768
rect 157246 271824 157302 271833
rect 157246 271759 157302 271768
rect 151360 271730 151412 271736
rect 157260 271726 157288 271759
rect 125600 271720 125652 271726
rect 115938 271688 115994 271697
rect 115938 271623 115994 271632
rect 117318 271688 117374 271697
rect 117318 271623 117374 271632
rect 120078 271688 120134 271697
rect 125600 271662 125652 271668
rect 157248 271720 157300 271726
rect 157248 271662 157300 271668
rect 158626 271688 158682 271697
rect 120078 271623 120080 271632
rect 115846 271552 115902 271561
rect 115952 271522 115980 271623
rect 117332 271590 117360 271623
rect 120132 271623 120134 271632
rect 158626 271623 158628 271632
rect 120080 271594 120132 271600
rect 158680 271623 158682 271632
rect 161294 271688 161350 271697
rect 161294 271623 161350 271632
rect 164146 271688 164202 271697
rect 164146 271623 164202 271632
rect 158628 271594 158680 271600
rect 161308 271590 161336 271623
rect 117320 271584 117372 271590
rect 117320 271526 117372 271532
rect 161296 271584 161348 271590
rect 161296 271526 161348 271532
rect 164160 271522 164188 271623
rect 115846 271487 115902 271496
rect 115940 271516 115992 271522
rect 115860 269890 115888 271487
rect 115940 271458 115992 271464
rect 164148 271516 164200 271522
rect 164148 271458 164200 271464
rect 183466 271416 183522 271425
rect 183466 271351 183522 271360
rect 183480 271318 183508 271351
rect 183468 271312 183520 271318
rect 183468 271254 183520 271260
rect 183468 271176 183520 271182
rect 183466 271144 183468 271153
rect 183520 271144 183522 271153
rect 183466 271079 183522 271088
rect 129738 271008 129794 271017
rect 129738 270943 129794 270952
rect 129752 270502 129780 270943
rect 147678 270736 147734 270745
rect 147678 270671 147734 270680
rect 129740 270496 129792 270502
rect 129740 270438 129792 270444
rect 115848 269884 115900 269890
rect 115848 269826 115900 269832
rect 113364 269816 113416 269822
rect 113364 269758 113416 269764
rect 147692 268802 147720 270671
rect 147680 268796 147732 268802
rect 147680 268738 147732 268744
rect 191748 253904 191800 253910
rect 191748 253846 191800 253852
rect 191760 253745 191788 253846
rect 191746 253736 191802 253745
rect 191746 253671 191802 253680
rect 180524 253292 180576 253298
rect 180524 253234 180576 253240
rect 179328 253224 179380 253230
rect 179326 253192 179328 253201
rect 180536 253201 180564 253234
rect 179380 253192 179382 253201
rect 179326 253127 179382 253136
rect 180522 253192 180578 253201
rect 180522 253127 180578 253136
rect 106924 251864 106976 251870
rect 106924 251806 106976 251812
rect 62120 251388 62172 251394
rect 62120 251330 62172 251336
rect 98460 167000 98512 167006
rect 98460 166942 98512 166948
rect 98472 166841 98500 166942
rect 101036 166932 101088 166938
rect 101036 166874 101088 166880
rect 101048 166841 101076 166874
rect 105820 166864 105872 166870
rect 98458 166832 98514 166841
rect 98458 166767 98514 166776
rect 101034 166832 101090 166841
rect 101034 166767 101090 166776
rect 105818 166832 105820 166841
rect 105872 166832 105874 166841
rect 105818 166767 105874 166776
rect 108210 166832 108266 166841
rect 108210 166767 108212 166776
rect 108264 166767 108266 166776
rect 138478 166832 138534 166841
rect 138478 166767 138534 166776
rect 140870 166832 140926 166841
rect 140870 166767 140926 166776
rect 145930 166832 145986 166841
rect 145930 166767 145986 166776
rect 108212 166738 108264 166744
rect 138492 166734 138520 166767
rect 138480 166728 138532 166734
rect 138480 166670 138532 166676
rect 140884 166666 140912 166767
rect 140872 166660 140924 166666
rect 140872 166602 140924 166608
rect 145944 166598 145972 166767
rect 163318 166696 163374 166705
rect 163318 166631 163374 166640
rect 165894 166696 165950 166705
rect 165894 166631 165950 166640
rect 60004 166592 60056 166598
rect 145932 166592 145984 166598
rect 60004 166534 60056 166540
rect 114374 166560 114430 166569
rect 114374 166495 114430 166504
rect 116950 166560 117006 166569
rect 145932 166534 145984 166540
rect 148506 166560 148562 166569
rect 116950 166495 117006 166504
rect 148506 166495 148508 166504
rect 96066 166288 96122 166297
rect 96066 166223 96068 166232
rect 96120 166223 96122 166232
rect 96068 166194 96120 166200
rect 114388 165714 114416 166495
rect 114376 165708 114428 165714
rect 114376 165650 114428 165656
rect 116964 165646 116992 166495
rect 148560 166495 148562 166504
rect 153290 166560 153346 166569
rect 153290 166495 153346 166504
rect 148508 166466 148560 166472
rect 153304 166462 153332 166495
rect 153292 166456 153344 166462
rect 153292 166398 153344 166404
rect 163332 166394 163360 166631
rect 163320 166388 163372 166394
rect 163320 166330 163372 166336
rect 165908 166326 165936 166631
rect 183282 166560 183338 166569
rect 183282 166495 183338 166504
rect 165896 166320 165948 166326
rect 165896 166262 165948 166268
rect 116952 165640 117004 165646
rect 81438 165608 81494 165617
rect 81438 165543 81494 165552
rect 84198 165608 84254 165617
rect 84198 165543 84254 165552
rect 89994 165608 90050 165617
rect 89994 165543 90050 165552
rect 91098 165608 91154 165617
rect 91098 165543 91154 165552
rect 95238 165608 95294 165617
rect 95238 165543 95294 165552
rect 99378 165608 99434 165617
rect 99378 165543 99434 165552
rect 103518 165608 103574 165617
rect 103518 165543 103574 165552
rect 109498 165608 109554 165617
rect 109498 165543 109554 165552
rect 110878 165608 110934 165617
rect 110878 165543 110934 165552
rect 111154 165608 111210 165617
rect 111154 165543 111210 165552
rect 113178 165608 113234 165617
rect 113178 165543 113234 165552
rect 113546 165608 113602 165617
rect 113546 165543 113602 165552
rect 115938 165608 115994 165617
rect 116952 165582 117004 165588
rect 117962 165608 118018 165617
rect 115938 165543 115994 165552
rect 117962 165543 118018 165552
rect 118330 165608 118386 165617
rect 118330 165543 118386 165552
rect 118974 165608 119030 165617
rect 118974 165543 119030 165552
rect 120906 165608 120962 165617
rect 120906 165543 120962 165552
rect 123482 165608 123538 165617
rect 123482 165543 123538 165552
rect 125874 165608 125930 165617
rect 125874 165543 125930 165552
rect 128358 165608 128414 165617
rect 128358 165543 128414 165552
rect 129738 165608 129794 165617
rect 129738 165543 129794 165552
rect 132498 165608 132554 165617
rect 132498 165543 132500 165552
rect 59910 165200 59966 165209
rect 59910 165135 59966 165144
rect 76010 164384 76066 164393
rect 76010 164319 76066 164328
rect 75918 164248 75974 164257
rect 60004 164212 60056 164218
rect 75918 164183 75974 164192
rect 60004 164154 60056 164160
rect 60016 163742 60044 164154
rect 60004 163736 60056 163742
rect 60004 163678 60056 163684
rect 59912 148844 59964 148850
rect 59912 148786 59964 148792
rect 59820 146260 59872 146266
rect 59820 146202 59872 146208
rect 59726 146160 59782 146169
rect 59726 146095 59782 146104
rect 59358 140856 59414 140865
rect 59358 140791 59414 140800
rect 59832 59226 59860 146202
rect 59820 59220 59872 59226
rect 59820 59162 59872 59168
rect 59268 57384 59320 57390
rect 59268 57326 59320 57332
rect 59176 57316 59228 57322
rect 59176 57258 59228 57264
rect 59924 56370 59952 148786
rect 59912 56364 59964 56370
rect 59912 56306 59964 56312
rect 58808 56092 58860 56098
rect 58808 56034 58860 56040
rect 60016 54874 60044 163678
rect 75932 145382 75960 164183
rect 76024 145450 76052 164319
rect 77298 164248 77354 164257
rect 77298 164183 77354 164192
rect 78678 164248 78734 164257
rect 78678 164183 78734 164192
rect 80058 164248 80114 164257
rect 80058 164183 80114 164192
rect 77312 145518 77340 164183
rect 78692 145858 78720 164183
rect 80072 148782 80100 164183
rect 80060 148776 80112 148782
rect 80060 148718 80112 148724
rect 81452 148646 81480 165543
rect 83464 164416 83516 164422
rect 83464 164358 83516 164364
rect 82818 164248 82874 164257
rect 82818 164183 82874 164192
rect 81440 148640 81492 148646
rect 81440 148582 81492 148588
rect 82832 145994 82860 164183
rect 83476 148850 83504 164358
rect 83464 148844 83516 148850
rect 83464 148786 83516 148792
rect 82820 145988 82872 145994
rect 82820 145930 82872 145936
rect 84212 145926 84240 165543
rect 88338 164928 88394 164937
rect 90008 164898 90036 165543
rect 88338 164863 88394 164872
rect 89996 164892 90048 164898
rect 88352 164830 88380 164863
rect 89996 164834 90048 164840
rect 88340 164824 88392 164830
rect 88340 164766 88392 164772
rect 89902 164384 89958 164393
rect 87604 164348 87656 164354
rect 89902 164319 89958 164328
rect 87604 164290 87656 164296
rect 84290 164248 84346 164257
rect 84290 164183 84346 164192
rect 85578 164248 85634 164257
rect 85578 164183 85634 164192
rect 86958 164248 87014 164257
rect 86958 164183 87014 164192
rect 84200 145920 84252 145926
rect 84200 145862 84252 145868
rect 78680 145852 78732 145858
rect 78680 145794 78732 145800
rect 84304 145790 84332 164183
rect 84292 145784 84344 145790
rect 84292 145726 84344 145732
rect 85592 145722 85620 164183
rect 86972 146062 87000 164183
rect 87616 148714 87644 164290
rect 88430 164248 88486 164257
rect 88430 164183 88486 164192
rect 87604 148708 87656 148714
rect 87604 148650 87656 148656
rect 88444 146130 88472 164183
rect 89916 162178 89944 164319
rect 89904 162172 89956 162178
rect 89904 162114 89956 162120
rect 88432 146124 88484 146130
rect 88432 146066 88484 146072
rect 86960 146056 87012 146062
rect 86960 145998 87012 146004
rect 85580 145716 85632 145722
rect 85580 145658 85632 145664
rect 91112 145654 91140 165543
rect 91190 164248 91246 164257
rect 91190 164183 91246 164192
rect 92478 164248 92534 164257
rect 92478 164183 92534 164192
rect 93858 164248 93914 164257
rect 93858 164183 93914 164192
rect 91204 146198 91232 164183
rect 91192 146192 91244 146198
rect 91192 146134 91244 146140
rect 92492 145761 92520 164183
rect 93872 146266 93900 164183
rect 95252 163878 95280 165543
rect 98644 164484 98696 164490
rect 98644 164426 98696 164432
rect 96618 164248 96674 164257
rect 96618 164183 96674 164192
rect 97998 164248 98054 164257
rect 97998 164183 98054 164192
rect 95240 163872 95292 163878
rect 95240 163814 95292 163820
rect 96632 163810 96660 164183
rect 96620 163804 96672 163810
rect 96620 163746 96672 163752
rect 93860 146260 93912 146266
rect 93860 146202 93912 146208
rect 92478 145752 92534 145761
rect 92478 145687 92534 145696
rect 91100 145648 91152 145654
rect 91100 145590 91152 145596
rect 98012 145586 98040 164183
rect 98656 145625 98684 164426
rect 99392 146169 99420 165543
rect 103532 164966 103560 165543
rect 103520 164960 103572 164966
rect 103520 164902 103572 164908
rect 107658 164928 107714 164937
rect 107658 164863 107714 164872
rect 106278 164792 106334 164801
rect 106278 164727 106334 164736
rect 100758 164520 100814 164529
rect 100758 164455 100760 164464
rect 100812 164455 100814 164464
rect 100760 164426 100812 164432
rect 106292 164354 106320 164727
rect 107672 164422 107700 164863
rect 107660 164416 107712 164422
rect 107660 164358 107712 164364
rect 106280 164348 106332 164354
rect 106280 164290 106332 164296
rect 100022 164248 100078 164257
rect 100022 164183 100078 164192
rect 102138 164248 102194 164257
rect 102138 164183 102194 164192
rect 103518 164248 103574 164257
rect 103518 164183 103574 164192
rect 106186 164248 106242 164257
rect 106370 164248 106426 164257
rect 106242 164206 106320 164234
rect 106186 164183 106242 164192
rect 100036 146305 100064 164183
rect 102152 148578 102180 164183
rect 103532 148986 103560 164183
rect 106292 149054 106320 164206
rect 106370 164183 106426 164192
rect 106384 163742 106412 164183
rect 106372 163736 106424 163742
rect 106372 163678 106424 163684
rect 109512 163674 109540 165543
rect 110892 164150 110920 165543
rect 110880 164144 110932 164150
rect 110880 164086 110932 164092
rect 109500 163668 109552 163674
rect 109500 163610 109552 163616
rect 111168 163538 111196 165543
rect 113192 164898 113220 165543
rect 113560 165102 113588 165543
rect 113548 165096 113600 165102
rect 113548 165038 113600 165044
rect 115952 165034 115980 165543
rect 115940 165028 115992 165034
rect 115940 164970 115992 164976
rect 114560 164960 114612 164966
rect 114560 164902 114612 164908
rect 113180 164892 113232 164898
rect 113180 164834 113232 164840
rect 111156 163532 111208 163538
rect 111156 163474 111208 163480
rect 106280 149048 106332 149054
rect 106280 148990 106332 148996
rect 103520 148980 103572 148986
rect 103520 148922 103572 148928
rect 102140 148572 102192 148578
rect 102140 148514 102192 148520
rect 113192 148510 113220 164834
rect 114572 164529 114600 164902
rect 115940 164824 115992 164830
rect 115940 164766 115992 164772
rect 115952 164529 115980 164766
rect 114558 164520 114614 164529
rect 114558 164455 114614 164464
rect 115938 164520 115994 164529
rect 115938 164455 115994 164464
rect 113180 148504 113232 148510
rect 113180 148446 113232 148452
rect 114572 148442 114600 164455
rect 114560 148436 114612 148442
rect 114560 148378 114612 148384
rect 115952 148374 115980 164455
rect 117976 164218 118004 165543
rect 118344 165170 118372 165543
rect 118332 165164 118384 165170
rect 118332 165106 118384 165112
rect 117964 164212 118016 164218
rect 117964 164154 118016 164160
rect 118988 163606 119016 165543
rect 120920 165306 120948 165543
rect 120908 165300 120960 165306
rect 120908 165242 120960 165248
rect 123496 165238 123524 165543
rect 125888 165374 125916 165543
rect 128372 165442 128400 165543
rect 129752 165510 129780 165543
rect 132552 165543 132554 165552
rect 132500 165514 132552 165520
rect 129740 165504 129792 165510
rect 129740 165446 129792 165452
rect 128360 165436 128412 165442
rect 128360 165378 128412 165384
rect 125876 165368 125928 165374
rect 125876 165310 125928 165316
rect 183296 165238 183324 166495
rect 183374 165608 183430 165617
rect 183374 165543 183430 165552
rect 123484 165232 123536 165238
rect 123484 165174 123536 165180
rect 183284 165232 183336 165238
rect 183284 165174 183336 165180
rect 183388 165102 183416 165543
rect 183376 165096 183428 165102
rect 183376 165038 183428 165044
rect 196636 164898 196664 271866
rect 197360 271448 197412 271454
rect 197360 271390 197412 271396
rect 197372 271318 197400 271390
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 196716 270496 196768 270502
rect 196716 270438 196768 270444
rect 196728 269822 196756 270438
rect 196716 269816 196768 269822
rect 196716 269758 196768 269764
rect 196728 164966 196756 269758
rect 197372 165238 197400 271254
rect 197464 253230 197492 354646
rect 197556 253298 197584 359654
rect 197648 271454 197676 374614
rect 197740 271522 197768 468590
rect 197820 464500 197872 464506
rect 197820 464442 197872 464448
rect 197728 271516 197780 271522
rect 197728 271458 197780 271464
rect 197636 271448 197688 271454
rect 197636 271390 197688 271396
rect 197832 270502 197860 464442
rect 197924 382226 197952 486610
rect 198200 484158 198228 488022
rect 199108 486736 199160 486742
rect 199108 486678 199160 486684
rect 198372 486600 198424 486606
rect 198372 486542 198424 486548
rect 198188 484152 198240 484158
rect 198188 484094 198240 484100
rect 198004 482452 198056 482458
rect 198004 482394 198056 482400
rect 198016 396030 198044 482394
rect 198096 464568 198148 464574
rect 198096 464510 198148 464516
rect 198004 396024 198056 396030
rect 198004 395966 198056 395972
rect 197912 382220 197964 382226
rect 197912 382162 197964 382168
rect 198108 380050 198136 464510
rect 198188 396364 198240 396370
rect 198188 396306 198240 396312
rect 198096 380044 198148 380050
rect 198096 379986 198148 379992
rect 198200 377398 198228 396306
rect 198280 395548 198332 395554
rect 198280 395490 198332 395496
rect 198292 380322 198320 395490
rect 198280 380316 198332 380322
rect 198280 380258 198332 380264
rect 198188 377392 198240 377398
rect 198188 377334 198240 377340
rect 198384 271658 198412 486542
rect 198740 484220 198792 484226
rect 198740 484162 198792 484168
rect 198752 377398 198780 484162
rect 199120 483970 199148 486678
rect 199212 484106 199240 488022
rect 199396 485178 199424 488022
rect 199488 488022 199778 488050
rect 199384 485172 199436 485178
rect 199384 485114 199436 485120
rect 199488 484226 199516 488022
rect 200224 485110 200252 488036
rect 200316 488022 200698 488050
rect 200776 488022 201066 488050
rect 201542 488022 201724 488050
rect 200212 485104 200264 485110
rect 200212 485046 200264 485052
rect 199476 484220 199528 484226
rect 199476 484162 199528 484168
rect 200316 484140 200344 488022
rect 200488 485444 200540 485450
rect 200488 485386 200540 485392
rect 200500 485353 200528 485386
rect 200486 485344 200542 485353
rect 200486 485279 200542 485288
rect 200132 484112 200344 484140
rect 199212 484078 199792 484106
rect 199120 483942 199240 483970
rect 199108 482520 199160 482526
rect 199108 482462 199160 482468
rect 198924 468580 198976 468586
rect 198924 468522 198976 468528
rect 198832 465724 198884 465730
rect 198832 465666 198884 465672
rect 198844 465118 198872 465666
rect 198832 465112 198884 465118
rect 198832 465054 198884 465060
rect 198832 400920 198884 400926
rect 198830 400888 198832 400897
rect 198884 400888 198886 400897
rect 198830 400823 198886 400832
rect 198832 396024 198884 396030
rect 198832 395966 198884 395972
rect 198844 380186 198872 395966
rect 198832 380180 198884 380186
rect 198832 380122 198884 380128
rect 198740 377392 198792 377398
rect 198740 377334 198792 377340
rect 198830 351928 198886 351937
rect 198830 351863 198886 351872
rect 198738 289776 198794 289785
rect 198738 289711 198794 289720
rect 198752 288833 198780 289711
rect 198738 288824 198794 288833
rect 198738 288759 198794 288768
rect 198372 271652 198424 271658
rect 198372 271594 198424 271600
rect 197820 270496 197872 270502
rect 197820 270438 197872 270444
rect 197728 269884 197780 269890
rect 197728 269826 197780 269832
rect 197544 253292 197596 253298
rect 197544 253234 197596 253240
rect 197452 253224 197504 253230
rect 197452 253166 197504 253172
rect 197452 167000 197504 167006
rect 197452 166942 197504 166948
rect 197360 165232 197412 165238
rect 197360 165174 197412 165180
rect 196716 164960 196768 164966
rect 196716 164902 196768 164908
rect 196624 164892 196676 164898
rect 196624 164834 196676 164840
rect 118976 163600 119028 163606
rect 118976 163542 119028 163548
rect 115940 148368 115992 148374
rect 115940 148310 115992 148316
rect 100022 146296 100078 146305
rect 100022 146231 100078 146240
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 99378 146160 99434 146169
rect 99378 146095 99434 146104
rect 98642 145616 98698 145625
rect 98000 145580 98052 145586
rect 98642 145551 98698 145560
rect 98000 145522 98052 145528
rect 77300 145512 77352 145518
rect 77300 145454 77352 145460
rect 76012 145444 76064 145450
rect 76012 145386 76064 145392
rect 75920 145376 75972 145382
rect 75920 145318 75972 145324
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 191288 145580 191340 145586
rect 191288 145522 191340 145528
rect 191300 144945 191328 145522
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 191286 144936 191342 144945
rect 191286 144871 191342 144880
rect 77114 59800 77170 59809
rect 77114 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 94502 59800 94558 59809
rect 94502 59735 94558 59744
rect 101770 59800 101826 59809
rect 101770 59735 101826 59744
rect 102782 59800 102838 59809
rect 102782 59735 102838 59744
rect 113546 59800 113602 59809
rect 113546 59735 113602 59744
rect 77128 59702 77156 59735
rect 77116 59696 77168 59702
rect 77116 59638 77168 59644
rect 83108 59634 83136 59735
rect 83096 59628 83148 59634
rect 83096 59570 83148 59576
rect 89994 59528 90050 59537
rect 89994 59463 90050 59472
rect 84200 59356 84252 59362
rect 84200 59298 84252 59304
rect 84212 58041 84240 59298
rect 90008 59294 90036 59463
rect 89996 59288 90048 59294
rect 89996 59230 90048 59236
rect 94516 59226 94544 59735
rect 100760 59560 100812 59566
rect 95882 59528 95938 59537
rect 95882 59463 95938 59472
rect 96986 59528 97042 59537
rect 96986 59463 97042 59472
rect 98090 59528 98146 59537
rect 98090 59463 98146 59472
rect 100758 59528 100760 59537
rect 100812 59528 100814 59537
rect 101784 59498 101812 59735
rect 100758 59463 100814 59472
rect 101772 59492 101824 59498
rect 94504 59220 94556 59226
rect 94504 59162 94556 59168
rect 95896 59158 95924 59463
rect 95884 59152 95936 59158
rect 95884 59094 95936 59100
rect 97000 59090 97028 59463
rect 96988 59084 97040 59090
rect 96988 59026 97040 59032
rect 98104 59022 98132 59463
rect 101772 59434 101824 59440
rect 98092 59016 98144 59022
rect 98092 58958 98144 58964
rect 102796 58954 102824 59735
rect 107566 59664 107622 59673
rect 107566 59599 107622 59608
rect 102784 58948 102836 58954
rect 102784 58890 102836 58896
rect 107580 58886 107608 59599
rect 113560 59430 113588 59735
rect 113548 59424 113600 59430
rect 110970 59392 111026 59401
rect 113548 59366 113600 59372
rect 110970 59327 111026 59336
rect 107568 58880 107620 58886
rect 107568 58822 107620 58828
rect 110984 58818 111012 59327
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 110972 58812 111024 58818
rect 110972 58754 111024 58760
rect 148520 58750 148548 59191
rect 148508 58744 148560 58750
rect 148508 58686 148560 58692
rect 150912 58682 150940 59191
rect 150900 58676 150952 58682
rect 150900 58618 150952 58624
rect 84198 58032 84254 58041
rect 84198 57967 84254 57976
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 78678 57896 78734 57905
rect 78678 57831 78734 57840
rect 80426 57896 80482 57905
rect 80426 57831 80482 57840
rect 81438 57896 81494 57905
rect 81438 57831 81494 57840
rect 85394 57896 85450 57905
rect 85394 57831 85450 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88338 57896 88394 57905
rect 88338 57831 88394 57840
rect 88706 57896 88762 57905
rect 88706 57831 88762 57840
rect 90730 57896 90786 57905
rect 90730 57831 90786 57840
rect 91098 57896 91154 57905
rect 91098 57831 91154 57840
rect 91466 57896 91522 57905
rect 91466 57831 91522 57840
rect 93306 57896 93362 57905
rect 93306 57831 93362 57840
rect 93674 57896 93730 57905
rect 93674 57831 93730 57840
rect 99378 57896 99434 57905
rect 99378 57831 99434 57840
rect 103794 57896 103850 57905
rect 103794 57831 103850 57840
rect 106278 57896 106334 57905
rect 106278 57831 106334 57840
rect 108210 57896 108266 57905
rect 108210 57831 108266 57840
rect 109038 57896 109094 57905
rect 109038 57831 109094 57840
rect 111154 57896 111210 57905
rect 111154 57831 111210 57840
rect 112074 57896 112130 57905
rect 112074 57831 112130 57840
rect 113178 57896 113234 57905
rect 113178 57831 113234 57840
rect 115754 57896 115810 57905
rect 115754 57831 115810 57840
rect 115938 57896 115994 57905
rect 115938 57831 115994 57840
rect 119066 57896 119122 57905
rect 119066 57831 119122 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 133418 57896 133474 57905
rect 133418 57831 133474 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 76024 57186 76052 57831
rect 78232 57254 78260 57831
rect 78220 57248 78272 57254
rect 78220 57190 78272 57196
rect 76012 57180 76064 57186
rect 76012 57122 76064 57128
rect 78692 55214 78720 57831
rect 80440 56030 80468 57831
rect 80428 56024 80480 56030
rect 80428 55966 80480 55972
rect 78680 55208 78732 55214
rect 78680 55150 78732 55156
rect 60004 54868 60056 54874
rect 60004 54810 60056 54816
rect 58624 54664 58676 54670
rect 58624 54606 58676 54612
rect 81452 54602 81480 57831
rect 85408 56098 85436 57831
rect 86512 56166 86540 57831
rect 86500 56160 86552 56166
rect 86500 56102 86552 56108
rect 85396 56092 85448 56098
rect 85396 56034 85448 56040
rect 86972 54738 87000 57831
rect 88352 57458 88380 57831
rect 88340 57452 88392 57458
rect 88340 57394 88392 57400
rect 88720 56234 88748 57831
rect 90744 57322 90772 57831
rect 90732 57316 90784 57322
rect 90732 57258 90784 57264
rect 88708 56228 88760 56234
rect 88708 56170 88760 56176
rect 91112 54806 91140 57831
rect 91100 54800 91152 54806
rect 91100 54742 91152 54748
rect 86960 54732 87012 54738
rect 86960 54674 87012 54680
rect 91480 54670 91508 57831
rect 93320 56302 93348 57831
rect 93688 57390 93716 57831
rect 99392 57526 99420 57831
rect 103808 57594 103836 57831
rect 103796 57588 103848 57594
rect 103796 57530 103848 57536
rect 99380 57520 99432 57526
rect 99380 57462 99432 57468
rect 93676 57384 93728 57390
rect 93676 57326 93728 57332
rect 93308 56296 93360 56302
rect 93308 56238 93360 56244
rect 106292 54874 106320 57831
rect 108224 56370 108252 57831
rect 108212 56364 108264 56370
rect 108212 56306 108264 56312
rect 109052 54942 109080 57831
rect 111168 56506 111196 57831
rect 111156 56500 111208 56506
rect 111156 56442 111208 56448
rect 112088 56438 112116 57831
rect 112076 56432 112128 56438
rect 112076 56374 112128 56380
rect 113192 55078 113220 57831
rect 113270 57352 113326 57361
rect 113270 57287 113326 57296
rect 113180 55072 113232 55078
rect 113180 55014 113232 55020
rect 113284 55010 113312 57287
rect 115768 56574 115796 57831
rect 115952 57662 115980 57831
rect 115940 57656 115992 57662
rect 115846 57624 115902 57633
rect 115940 57598 115992 57604
rect 116122 57624 116178 57633
rect 115846 57559 115902 57568
rect 116122 57559 116178 57568
rect 115860 57361 115888 57559
rect 115846 57352 115902 57361
rect 115846 57287 115902 57296
rect 115756 56568 115808 56574
rect 115756 56510 115808 56516
rect 116136 55146 116164 57559
rect 119080 56137 119108 57831
rect 130856 57730 130884 57831
rect 133432 57798 133460 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 183466 57896 183522 57905
rect 183466 57831 183468 57840
rect 145564 57802 145616 57808
rect 133420 57792 133472 57798
rect 133420 57734 133472 57740
rect 130844 57724 130896 57730
rect 130844 57666 130896 57672
rect 122838 57624 122894 57633
rect 122838 57559 122894 57568
rect 119066 56128 119122 56137
rect 119066 56063 119122 56072
rect 116124 55140 116176 55146
rect 116124 55082 116176 55088
rect 113272 55004 113324 55010
rect 113272 54946 113324 54952
rect 109040 54936 109092 54942
rect 109040 54878 109092 54884
rect 106280 54868 106332 54874
rect 106280 54810 106332 54816
rect 91468 54664 91520 54670
rect 91468 54606 91520 54612
rect 81440 54596 81492 54602
rect 81440 54538 81492 54544
rect 122852 54534 122880 57559
rect 153304 56273 153332 57831
rect 183520 57831 183522 57840
rect 183468 57802 183520 57808
rect 197372 57798 197400 165174
rect 197464 165102 197492 166942
rect 197452 165096 197504 165102
rect 197452 165038 197504 165044
rect 197464 57866 197492 165038
rect 197556 146198 197584 253234
rect 197636 253224 197688 253230
rect 197636 253166 197688 253172
rect 197648 146266 197676 253166
rect 197740 164830 197768 269826
rect 198752 181937 198780 288759
rect 198844 246265 198872 351863
rect 198936 271794 198964 468522
rect 199016 465112 199068 465118
rect 199016 465054 199068 465060
rect 199028 460193 199056 465054
rect 199014 460184 199070 460193
rect 199014 460119 199070 460128
rect 199028 353161 199056 460119
rect 199120 380254 199148 482462
rect 199212 396370 199240 483942
rect 199292 479528 199344 479534
rect 199292 479470 199344 479476
rect 199200 396364 199252 396370
rect 199200 396306 199252 396312
rect 199304 394641 199332 479470
rect 199384 478168 199436 478174
rect 199384 478110 199436 478116
rect 199396 397361 199424 478110
rect 199476 475380 199528 475386
rect 199476 475322 199528 475328
rect 199488 400926 199516 475322
rect 199568 464364 199620 464370
rect 199568 464306 199620 464312
rect 199476 400920 199528 400926
rect 199476 400862 199528 400868
rect 199474 398168 199530 398177
rect 199474 398103 199530 398112
rect 199382 397352 199438 397361
rect 199382 397287 199438 397296
rect 199290 394632 199346 394641
rect 199290 394567 199346 394576
rect 199304 384334 199332 394567
rect 199292 384328 199344 384334
rect 199292 384270 199344 384276
rect 199108 380248 199160 380254
rect 199108 380190 199160 380196
rect 199488 378078 199516 398103
rect 199580 395554 199608 464306
rect 199568 395548 199620 395554
rect 199568 395490 199620 395496
rect 199566 395312 199622 395321
rect 199566 395247 199622 395256
rect 199476 378072 199528 378078
rect 199476 378014 199528 378020
rect 199384 371884 199436 371890
rect 199384 371826 199436 371832
rect 199014 353152 199070 353161
rect 199014 353087 199070 353096
rect 199028 351937 199056 353087
rect 199014 351928 199070 351937
rect 199014 351863 199070 351872
rect 199290 292768 199346 292777
rect 199290 292703 199346 292712
rect 199014 291680 199070 291689
rect 199014 291615 199070 291624
rect 198924 271788 198976 271794
rect 198924 271730 198976 271736
rect 198830 246256 198886 246265
rect 198830 246191 198886 246200
rect 198738 181928 198794 181937
rect 198738 181863 198794 181872
rect 197728 164824 197780 164830
rect 197728 164766 197780 164772
rect 197636 146260 197688 146266
rect 197636 146202 197688 146208
rect 197544 146192 197596 146198
rect 197544 146134 197596 146140
rect 198752 74905 198780 181863
rect 198844 139233 198872 246191
rect 199028 184929 199056 291615
rect 199198 291000 199254 291009
rect 199198 290935 199254 290944
rect 199106 288416 199162 288425
rect 199106 288351 199162 288360
rect 199120 287609 199148 288351
rect 199106 287600 199162 287609
rect 199106 287535 199162 287544
rect 199014 184920 199070 184929
rect 198936 184878 199014 184906
rect 198830 139224 198886 139233
rect 198830 139159 198886 139168
rect 198936 77761 198964 184878
rect 199014 184855 199070 184864
rect 199014 183560 199070 183569
rect 199014 183495 199070 183504
rect 198922 77752 198978 77761
rect 198922 77687 198978 77696
rect 199028 76401 199056 183495
rect 199120 180794 199148 287535
rect 199212 183569 199240 290935
rect 199304 186425 199332 292703
rect 199396 289785 199424 371826
rect 199488 370530 199516 378014
rect 199580 377466 199608 395247
rect 199660 384328 199712 384334
rect 199660 384270 199712 384276
rect 199568 377460 199620 377466
rect 199568 377402 199620 377408
rect 199580 371890 199608 377402
rect 199568 371884 199620 371890
rect 199568 371826 199620 371832
rect 199476 370524 199528 370530
rect 199476 370466 199528 370472
rect 199488 291689 199516 370466
rect 199568 369164 199620 369170
rect 199568 369106 199620 369112
rect 199580 292777 199608 369106
rect 199672 362234 199700 384270
rect 199764 377466 199792 484078
rect 199842 397352 199898 397361
rect 199842 397287 199898 397296
rect 199752 377460 199804 377466
rect 199752 377402 199804 377408
rect 199856 364334 199884 397287
rect 200132 380322 200160 484112
rect 200776 483970 200804 488022
rect 201316 485716 201368 485722
rect 201316 485658 201368 485664
rect 201408 485716 201460 485722
rect 201408 485658 201460 485664
rect 201328 485450 201356 485658
rect 201316 485444 201368 485450
rect 201316 485386 201368 485392
rect 200224 483942 200804 483970
rect 200120 380316 200172 380322
rect 200120 380258 200172 380264
rect 200224 380254 200252 483942
rect 200304 482588 200356 482594
rect 200304 482530 200356 482536
rect 200212 380248 200264 380254
rect 200212 380190 200264 380196
rect 200316 376582 200344 482530
rect 200764 479664 200816 479670
rect 200764 479606 200816 479612
rect 200396 471504 200448 471510
rect 200396 471446 200448 471452
rect 200408 377194 200436 471446
rect 200488 468716 200540 468722
rect 200488 468658 200540 468664
rect 200500 379982 200528 468658
rect 200580 464432 200632 464438
rect 200580 464374 200632 464380
rect 200592 380594 200620 464374
rect 200776 389162 200804 479606
rect 200856 471096 200908 471102
rect 200856 471038 200908 471044
rect 200764 389156 200816 389162
rect 200764 389098 200816 389104
rect 200580 380588 200632 380594
rect 200580 380530 200632 380536
rect 200488 379976 200540 379982
rect 200488 379918 200540 379924
rect 200396 377188 200448 377194
rect 200396 377130 200448 377136
rect 200304 376576 200356 376582
rect 200304 376518 200356 376524
rect 199764 364306 199884 364334
rect 199764 363662 199792 364306
rect 199752 363656 199804 363662
rect 199752 363598 199804 363604
rect 199660 362228 199712 362234
rect 199660 362170 199712 362176
rect 199566 292768 199622 292777
rect 199566 292703 199622 292712
rect 199474 291680 199530 291689
rect 199474 291615 199530 291624
rect 199382 289776 199438 289785
rect 199382 289711 199438 289720
rect 199672 288425 199700 362170
rect 199764 291009 199792 363598
rect 200764 359508 200816 359514
rect 200764 359450 200816 359456
rect 199750 291000 199806 291009
rect 199750 290935 199806 290944
rect 199658 288416 199714 288425
rect 199658 288351 199714 288360
rect 200776 282198 200804 359450
rect 200764 282192 200816 282198
rect 200764 282134 200816 282140
rect 200868 272678 200896 471038
rect 200948 465588 201000 465594
rect 200948 465530 201000 465536
rect 200960 284306 200988 465530
rect 201420 379166 201448 485658
rect 201500 485240 201552 485246
rect 201498 485208 201500 485217
rect 201552 485208 201554 485217
rect 201498 485143 201554 485152
rect 201592 484152 201644 484158
rect 201592 484094 201644 484100
rect 201500 474088 201552 474094
rect 201500 474030 201552 474036
rect 201408 379160 201460 379166
rect 201408 379102 201460 379108
rect 201420 378962 201448 379102
rect 201408 378956 201460 378962
rect 201408 378898 201460 378904
rect 201408 360256 201460 360262
rect 201408 360198 201460 360204
rect 201420 359514 201448 360198
rect 201408 359508 201460 359514
rect 201408 359450 201460 359456
rect 200948 284300 201000 284306
rect 200948 284242 201000 284248
rect 201408 282192 201460 282198
rect 201408 282134 201460 282140
rect 200856 272672 200908 272678
rect 200856 272614 200908 272620
rect 201420 253910 201448 282134
rect 201512 269890 201540 474030
rect 201604 376582 201632 484094
rect 201696 380186 201724 488022
rect 201972 484430 202000 488036
rect 202064 488022 202446 488050
rect 201960 484424 202012 484430
rect 201960 484366 202012 484372
rect 202064 484158 202092 488022
rect 202892 485081 202920 488036
rect 202984 488022 203274 488050
rect 202878 485072 202934 485081
rect 202878 485007 202934 485016
rect 202052 484152 202104 484158
rect 202984 484140 203012 488022
rect 203524 484900 203576 484906
rect 203524 484842 203576 484848
rect 202052 484094 202104 484100
rect 202892 484112 203012 484140
rect 201868 482384 201920 482390
rect 201868 482326 201920 482332
rect 201776 465792 201828 465798
rect 201776 465734 201828 465740
rect 201684 380180 201736 380186
rect 201684 380122 201736 380128
rect 201592 376576 201644 376582
rect 201592 376518 201644 376524
rect 201592 358080 201644 358086
rect 201592 358022 201644 358028
rect 201604 271182 201632 358022
rect 201788 271862 201816 465734
rect 201880 380390 201908 482326
rect 202144 472728 202196 472734
rect 202144 472670 202196 472676
rect 201868 380384 201920 380390
rect 201868 380326 201920 380332
rect 201776 271856 201828 271862
rect 201776 271798 201828 271804
rect 201592 271176 201644 271182
rect 201592 271118 201644 271124
rect 201500 269884 201552 269890
rect 201500 269826 201552 269832
rect 201408 253904 201460 253910
rect 201408 253846 201460 253852
rect 199290 186416 199346 186425
rect 199290 186351 199346 186360
rect 199198 183560 199254 183569
rect 199198 183495 199254 183504
rect 199120 180766 199240 180794
rect 199212 180713 199240 180766
rect 199198 180704 199254 180713
rect 199198 180639 199254 180648
rect 199014 76392 199070 76401
rect 199014 76327 199070 76336
rect 198738 74896 198794 74905
rect 198738 74831 198794 74840
rect 199212 73681 199240 180639
rect 199304 79393 199332 186351
rect 201604 167006 201632 271118
rect 202156 271114 202184 472670
rect 202420 471164 202472 471170
rect 202420 471106 202472 471112
rect 202328 470076 202380 470082
rect 202328 470018 202380 470024
rect 202236 469056 202288 469062
rect 202236 468998 202288 469004
rect 202144 271108 202196 271114
rect 202144 271050 202196 271056
rect 202144 176180 202196 176186
rect 202144 176122 202196 176128
rect 201592 167000 201644 167006
rect 201592 166942 201644 166948
rect 202156 145586 202184 176122
rect 202248 166326 202276 468998
rect 202340 271658 202368 470018
rect 202432 272882 202460 471106
rect 202512 465656 202564 465662
rect 202512 465598 202564 465604
rect 202420 272876 202472 272882
rect 202420 272818 202472 272824
rect 202524 272542 202552 465598
rect 202786 380760 202842 380769
rect 202786 380695 202842 380704
rect 202512 272536 202564 272542
rect 202512 272478 202564 272484
rect 202328 271652 202380 271658
rect 202328 271594 202380 271600
rect 202236 166320 202288 166326
rect 202236 166262 202288 166268
rect 202144 145580 202196 145586
rect 202144 145522 202196 145528
rect 199290 79384 199346 79393
rect 199290 79319 199346 79328
rect 199198 73672 199254 73681
rect 199198 73607 199254 73616
rect 202800 58886 202828 380695
rect 202892 375766 202920 484112
rect 202972 484016 203024 484022
rect 202972 483958 203024 483964
rect 202984 380497 203012 483958
rect 203156 471436 203208 471442
rect 203156 471378 203208 471384
rect 203064 468512 203116 468518
rect 203064 468454 203116 468460
rect 202970 380488 203026 380497
rect 202970 380423 203026 380432
rect 202970 379264 203026 379273
rect 202970 379199 203026 379208
rect 202984 378593 203012 379199
rect 202970 378584 203026 378593
rect 202970 378519 203026 378528
rect 202880 375760 202932 375766
rect 202880 375702 202932 375708
rect 203076 271726 203104 468454
rect 203168 380730 203196 471378
rect 203156 380724 203208 380730
rect 203156 380666 203208 380672
rect 203064 271720 203116 271726
rect 203064 271662 203116 271668
rect 202880 253904 202932 253910
rect 202880 253846 202932 253852
rect 202892 176662 202920 253846
rect 202880 176656 202932 176662
rect 202880 176598 202932 176604
rect 202892 176186 202920 176598
rect 202880 176180 202932 176186
rect 202880 176122 202932 176128
rect 203536 166530 203564 484842
rect 203720 482866 203748 488036
rect 203904 488022 204194 488050
rect 204364 488022 204654 488050
rect 204732 488022 205022 488050
rect 205192 488022 205482 488050
rect 205836 488022 205942 488050
rect 206112 488022 206402 488050
rect 206480 488022 206862 488050
rect 207246 488022 207336 488050
rect 203904 484022 203932 488022
rect 204260 485512 204312 485518
rect 204260 485454 204312 485460
rect 204272 485217 204300 485454
rect 204258 485208 204314 485217
rect 204258 485143 204314 485152
rect 204260 485036 204312 485042
rect 204260 484978 204312 484984
rect 204272 484945 204300 484978
rect 204258 484936 204314 484945
rect 204258 484871 204314 484880
rect 203984 484424 204036 484430
rect 203984 484366 204036 484372
rect 203892 484016 203944 484022
rect 203892 483958 203944 483964
rect 203708 482860 203760 482866
rect 203708 482802 203760 482808
rect 203800 471232 203852 471238
rect 203614 471200 203670 471209
rect 203800 471174 203852 471180
rect 203614 471135 203670 471144
rect 203628 166666 203656 471135
rect 203706 466032 203762 466041
rect 203706 465967 203762 465976
rect 203616 166660 203668 166666
rect 203616 166602 203668 166608
rect 203524 166524 203576 166530
rect 203524 166466 203576 166472
rect 203720 166462 203748 465967
rect 203812 272610 203840 471174
rect 203892 466200 203944 466206
rect 203892 466142 203944 466148
rect 203904 282878 203932 466142
rect 203996 378078 204024 484366
rect 203984 378072 204036 378078
rect 203984 378014 204036 378020
rect 204364 376718 204392 488022
rect 204444 484152 204496 484158
rect 204444 484094 204496 484100
rect 204456 411602 204484 484094
rect 204732 470594 204760 488022
rect 204812 486532 204864 486538
rect 204812 486474 204864 486480
rect 204548 470566 204760 470594
rect 204548 417790 204576 470566
rect 204628 466608 204680 466614
rect 204628 466550 204680 466556
rect 204536 417784 204588 417790
rect 204536 417726 204588 417732
rect 204444 411596 204496 411602
rect 204444 411538 204496 411544
rect 204352 376712 204404 376718
rect 204352 376654 204404 376660
rect 204640 359582 204668 466550
rect 204720 464772 204772 464778
rect 204720 464714 204772 464720
rect 204732 380458 204760 464714
rect 204720 380452 204772 380458
rect 204720 380394 204772 380400
rect 204628 359576 204680 359582
rect 204628 359518 204680 359524
rect 203892 282872 203944 282878
rect 203892 282814 203944 282820
rect 203800 272604 203852 272610
rect 203800 272546 203852 272552
rect 204824 271590 204852 486474
rect 204904 485784 204956 485790
rect 204904 485726 204956 485732
rect 204916 484838 204944 485726
rect 204904 484832 204956 484838
rect 204904 484774 204956 484780
rect 205192 484158 205220 488022
rect 205640 485308 205692 485314
rect 205640 485250 205692 485256
rect 205652 484809 205680 485250
rect 205638 484800 205694 484809
rect 205638 484735 205694 484744
rect 205732 484220 205784 484226
rect 205732 484162 205784 484168
rect 205180 484152 205232 484158
rect 205180 484094 205232 484100
rect 205640 484152 205692 484158
rect 205640 484094 205692 484100
rect 204996 478236 205048 478242
rect 204996 478178 205048 478184
rect 204904 466064 204956 466070
rect 204904 466006 204956 466012
rect 204812 271584 204864 271590
rect 204812 271526 204864 271532
rect 204916 178022 204944 466006
rect 205008 271522 205036 478178
rect 205088 471912 205140 471918
rect 205088 471854 205140 471860
rect 205100 272746 205128 471854
rect 205364 465724 205416 465730
rect 205364 465666 205416 465672
rect 205376 386414 205404 465666
rect 205456 414724 205508 414730
rect 205456 414666 205508 414672
rect 205284 386386 205404 386414
rect 205178 380760 205234 380769
rect 205178 380695 205234 380704
rect 205088 272740 205140 272746
rect 205088 272682 205140 272688
rect 204996 271516 205048 271522
rect 204996 271458 205048 271464
rect 204904 178016 204956 178022
rect 204904 177958 204956 177964
rect 203708 166456 203760 166462
rect 203708 166398 203760 166404
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204916 67658 204944 145522
rect 204904 67652 204956 67658
rect 204904 67594 204956 67600
rect 202788 58880 202840 58886
rect 202788 58822 202840 58828
rect 204916 57934 204944 67594
rect 205192 59090 205220 380695
rect 205284 379273 205312 386386
rect 205270 379264 205326 379273
rect 205270 379199 205326 379208
rect 205362 379128 205418 379137
rect 205468 379098 205496 414666
rect 205652 413302 205680 484094
rect 205744 414866 205772 484162
rect 205836 478174 205864 488022
rect 206112 484158 206140 488022
rect 206480 484226 206508 488022
rect 207112 487076 207164 487082
rect 207112 487018 207164 487024
rect 206836 485172 206888 485178
rect 206836 485114 206888 485120
rect 206468 484220 206520 484226
rect 206468 484162 206520 484168
rect 206100 484152 206152 484158
rect 206100 484094 206152 484100
rect 206376 483812 206428 483818
rect 206376 483754 206428 483760
rect 205824 478168 205876 478174
rect 205824 478110 205876 478116
rect 205824 474156 205876 474162
rect 205824 474098 205876 474104
rect 205732 414860 205784 414866
rect 205732 414802 205784 414808
rect 205640 413296 205692 413302
rect 205640 413238 205692 413244
rect 205640 411596 205692 411602
rect 205640 411538 205692 411544
rect 205652 410582 205680 411538
rect 205640 410576 205692 410582
rect 205640 410518 205692 410524
rect 205548 381540 205600 381546
rect 205548 381482 205600 381488
rect 205362 379063 205418 379072
rect 205456 379092 205508 379098
rect 205376 378536 205404 379063
rect 205456 379034 205508 379040
rect 205284 378508 205404 378536
rect 205284 269754 205312 378508
rect 205362 378448 205418 378457
rect 205362 378383 205418 378392
rect 205272 269748 205324 269754
rect 205272 269690 205324 269696
rect 205180 59084 205232 59090
rect 205180 59026 205232 59032
rect 205376 58750 205404 378383
rect 205364 58744 205416 58750
rect 205364 58686 205416 58692
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 183192 57792 183244 57798
rect 183190 57760 183192 57769
rect 197360 57792 197412 57798
rect 183244 57760 183246 57769
rect 197360 57734 197412 57740
rect 183190 57695 183246 57704
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 162858 57624 162914 57633
rect 162858 57559 162914 57568
rect 165618 57624 165674 57633
rect 165618 57559 165674 57568
rect 153290 56264 153346 56273
rect 153290 56199 153346 56208
rect 160112 54913 160140 57559
rect 162872 55049 162900 57559
rect 165632 55185 165660 57559
rect 205560 57390 205588 381482
rect 205836 380526 205864 474098
rect 205916 471368 205968 471374
rect 205916 471310 205968 471316
rect 205928 380662 205956 471310
rect 206284 466472 206336 466478
rect 206284 466414 206336 466420
rect 206296 389842 206324 466414
rect 206284 389836 206336 389842
rect 206284 389778 206336 389784
rect 205916 380656 205968 380662
rect 205916 380598 205968 380604
rect 205824 380520 205876 380526
rect 205824 380462 205876 380468
rect 205640 378888 205692 378894
rect 205640 378830 205692 378836
rect 206190 378856 206246 378865
rect 205652 378554 205680 378830
rect 206190 378791 206246 378800
rect 205640 378548 205692 378554
rect 205640 378490 205692 378496
rect 206204 270473 206232 378791
rect 206296 360262 206324 389778
rect 206284 360256 206336 360262
rect 206284 360198 206336 360204
rect 206388 271182 206416 483754
rect 206468 470008 206520 470014
rect 206468 469950 206520 469956
rect 206480 271726 206508 469950
rect 206560 467356 206612 467362
rect 206560 467298 206612 467304
rect 206468 271720 206520 271726
rect 206468 271662 206520 271668
rect 206376 271176 206428 271182
rect 206376 271118 206428 271124
rect 206572 271046 206600 467298
rect 206652 465520 206704 465526
rect 206652 465462 206704 465468
rect 206664 376650 206692 465462
rect 206744 410712 206796 410718
rect 206744 410654 206796 410660
rect 206652 376644 206704 376650
rect 206652 376586 206704 376592
rect 206756 374746 206784 410654
rect 206848 379030 206876 485114
rect 207020 484152 207072 484158
rect 207020 484094 207072 484100
rect 206926 415304 206982 415313
rect 206926 415239 206982 415248
rect 206836 379024 206888 379030
rect 206836 378966 206888 378972
rect 206836 378888 206888 378894
rect 206836 378830 206888 378836
rect 206744 374740 206796 374746
rect 206744 374682 206796 374688
rect 206560 271040 206612 271046
rect 206560 270982 206612 270988
rect 206190 270464 206246 270473
rect 206190 270399 206246 270408
rect 206742 270464 206798 270473
rect 206742 270399 206798 270408
rect 206756 147626 206784 270399
rect 206848 268394 206876 378830
rect 206836 268388 206888 268394
rect 206836 268330 206888 268336
rect 206744 147620 206796 147626
rect 206744 147562 206796 147568
rect 206940 58818 206968 415239
rect 207032 379930 207060 484094
rect 207124 466478 207152 487018
rect 207308 485774 207336 488022
rect 207400 488022 207690 488050
rect 207768 488022 208150 488050
rect 208412 488022 208610 488050
rect 208688 488022 209070 488050
rect 209148 488022 209438 488050
rect 207400 487082 207428 488022
rect 207388 487076 207440 487082
rect 207388 487018 207440 487024
rect 207308 485746 207428 485774
rect 207400 483970 207428 485746
rect 207768 484158 207796 488022
rect 207756 484152 207808 484158
rect 207756 484094 207808 484100
rect 207216 483942 207428 483970
rect 207216 474094 207244 483942
rect 207756 482724 207808 482730
rect 207756 482666 207808 482672
rect 207296 482316 207348 482322
rect 207296 482258 207348 482264
rect 207204 474088 207256 474094
rect 207204 474030 207256 474036
rect 207112 466472 207164 466478
rect 207112 466414 207164 466420
rect 207112 465860 207164 465866
rect 207112 465802 207164 465808
rect 207124 380118 207152 465802
rect 207204 400920 207256 400926
rect 207204 400862 207256 400868
rect 207112 380112 207164 380118
rect 207112 380054 207164 380060
rect 207032 379902 207152 379930
rect 207124 379574 207152 379902
rect 207112 379568 207164 379574
rect 207112 379510 207164 379516
rect 207018 379400 207074 379409
rect 207018 379335 207074 379344
rect 207032 378593 207060 379335
rect 207018 378584 207074 378593
rect 207018 378519 207074 378528
rect 207124 376446 207152 379510
rect 207112 376440 207164 376446
rect 207112 376382 207164 376388
rect 207216 369850 207244 400862
rect 207308 377330 207336 482258
rect 207664 476876 207716 476882
rect 207664 476818 207716 476824
rect 207296 377324 207348 377330
rect 207296 377266 207348 377272
rect 207020 369844 207072 369850
rect 207020 369786 207072 369792
rect 207204 369844 207256 369850
rect 207204 369786 207256 369792
rect 207032 369170 207060 369786
rect 207020 369164 207072 369170
rect 207020 369106 207072 369112
rect 207676 165306 207704 476818
rect 207768 175234 207796 482666
rect 207848 475516 207900 475522
rect 207848 475458 207900 475464
rect 207860 271250 207888 475458
rect 208032 468308 208084 468314
rect 208032 468250 208084 468256
rect 207940 466336 207992 466342
rect 207940 466278 207992 466284
rect 207952 273018 207980 466278
rect 208044 376106 208072 468250
rect 208124 466472 208176 466478
rect 208124 466414 208176 466420
rect 208136 417450 208164 466414
rect 208308 465792 208360 465798
rect 208308 465734 208360 465740
rect 208216 417784 208268 417790
rect 208216 417726 208268 417732
rect 208124 417444 208176 417450
rect 208124 417386 208176 417392
rect 208228 409154 208256 417726
rect 208216 409148 208268 409154
rect 208216 409090 208268 409096
rect 208214 378584 208270 378593
rect 208214 378519 208270 378528
rect 208122 378312 208178 378321
rect 208122 378247 208178 378256
rect 208032 376100 208084 376106
rect 208032 376042 208084 376048
rect 207940 273012 207992 273018
rect 207940 272954 207992 272960
rect 207848 271244 207900 271250
rect 207848 271186 207900 271192
rect 208136 269793 208164 378247
rect 208122 269784 208178 269793
rect 208122 269719 208178 269728
rect 208228 268530 208256 378519
rect 208320 378185 208348 465734
rect 208412 380934 208440 488022
rect 208492 485444 208544 485450
rect 208492 485386 208544 485392
rect 208504 485353 208532 485386
rect 208490 485344 208546 485353
rect 208490 485279 208546 485288
rect 208492 484152 208544 484158
rect 208492 484094 208544 484100
rect 208400 380928 208452 380934
rect 208400 380870 208452 380876
rect 208398 380760 208454 380769
rect 208398 380695 208454 380704
rect 208412 380361 208440 380695
rect 208398 380352 208454 380361
rect 208398 380287 208454 380296
rect 208504 379506 208532 484094
rect 208688 470594 208716 488022
rect 209148 484158 209176 488022
rect 209688 485376 209740 485382
rect 209688 485318 209740 485324
rect 209136 484152 209188 484158
rect 209136 484094 209188 484100
rect 209412 482860 209464 482866
rect 209412 482802 209464 482808
rect 209044 481024 209096 481030
rect 209044 480966 209096 480972
rect 208596 470566 208716 470594
rect 208492 379500 208544 379506
rect 208492 379442 208544 379448
rect 208492 379364 208544 379370
rect 208492 379306 208544 379312
rect 208398 379128 208454 379137
rect 208398 379063 208454 379072
rect 208412 378729 208440 379063
rect 208398 378720 208454 378729
rect 208398 378655 208454 378664
rect 208504 378418 208532 379306
rect 208492 378412 208544 378418
rect 208492 378354 208544 378360
rect 208596 378282 208624 470566
rect 208952 464840 209004 464846
rect 208952 464782 209004 464788
rect 208676 380928 208728 380934
rect 208676 380870 208728 380876
rect 208584 378276 208636 378282
rect 208584 378218 208636 378224
rect 208306 378176 208362 378185
rect 208306 378111 208362 378120
rect 208306 378040 208362 378049
rect 208306 377975 208362 377984
rect 208216 268524 208268 268530
rect 208216 268466 208268 268472
rect 207756 175228 207808 175234
rect 207756 175170 207808 175176
rect 207664 165300 207716 165306
rect 207664 165242 207716 165248
rect 206928 58812 206980 58818
rect 206928 58754 206980 58760
rect 208320 57866 208348 377975
rect 208688 375358 208716 380870
rect 208858 379536 208914 379545
rect 208858 379471 208914 379480
rect 208400 375352 208452 375358
rect 208400 375294 208452 375300
rect 208676 375352 208728 375358
rect 208676 375294 208728 375300
rect 208412 374882 208440 375294
rect 208400 374876 208452 374882
rect 208400 374818 208452 374824
rect 208308 57860 208360 57866
rect 208308 57802 208360 57808
rect 208872 57526 208900 379471
rect 208964 375970 208992 464782
rect 208952 375964 209004 375970
rect 208952 375906 209004 375912
rect 209056 70378 209084 480966
rect 209228 474360 209280 474366
rect 209228 474302 209280 474308
rect 209136 468988 209188 468994
rect 209136 468930 209188 468936
rect 209148 166394 209176 468930
rect 209240 271318 209268 474302
rect 209320 464636 209372 464642
rect 209320 464578 209372 464584
rect 209332 273086 209360 464578
rect 209424 391950 209452 482802
rect 209412 391944 209464 391950
rect 209412 391886 209464 391892
rect 209410 381576 209466 381585
rect 209410 381511 209466 381520
rect 209320 273080 209372 273086
rect 209320 273022 209372 273028
rect 209228 271312 209280 271318
rect 209228 271254 209280 271260
rect 209424 270473 209452 381511
rect 209700 380769 209728 485318
rect 209884 485246 209912 488036
rect 209976 488022 210358 488050
rect 210528 488022 210818 488050
rect 211202 488022 211384 488050
rect 211662 488022 211936 488050
rect 209780 485240 209832 485246
rect 209780 485182 209832 485188
rect 209872 485240 209924 485246
rect 209872 485182 209924 485188
rect 209792 485042 209820 485182
rect 209780 485036 209832 485042
rect 209780 484978 209832 484984
rect 209780 484152 209832 484158
rect 209780 484094 209832 484100
rect 209686 380760 209742 380769
rect 209686 380695 209742 380704
rect 209596 379364 209648 379370
rect 209596 379306 209648 379312
rect 209502 379128 209558 379137
rect 209502 379063 209558 379072
rect 209410 270464 209466 270473
rect 209410 270399 209466 270408
rect 209516 269929 209544 379063
rect 209502 269920 209558 269929
rect 209502 269855 209558 269864
rect 209504 269748 209556 269754
rect 209504 269690 209556 269696
rect 209136 166388 209188 166394
rect 209136 166330 209188 166336
rect 209516 144906 209544 269690
rect 209608 268462 209636 379306
rect 209792 378350 209820 484094
rect 209976 470594 210004 488022
rect 210528 484158 210556 488022
rect 211068 485512 211120 485518
rect 211068 485454 211120 485460
rect 210516 484152 210568 484158
rect 210516 484094 210568 484100
rect 210516 479596 210568 479602
rect 210516 479538 210568 479544
rect 209884 470566 210004 470594
rect 209884 379302 209912 470566
rect 210424 469872 210476 469878
rect 210424 469814 210476 469820
rect 209872 379296 209924 379302
rect 209872 379238 209924 379244
rect 210332 379092 210384 379098
rect 210332 379034 210384 379040
rect 210238 378720 210294 378729
rect 210238 378655 210294 378664
rect 209780 378344 209832 378350
rect 209780 378286 209832 378292
rect 209596 268456 209648 268462
rect 209596 268398 209648 268404
rect 209504 144900 209556 144906
rect 209504 144842 209556 144848
rect 209044 70372 209096 70378
rect 209044 70314 209096 70320
rect 210252 57934 210280 378655
rect 210344 378418 210372 379034
rect 210332 378412 210384 378418
rect 210332 378354 210384 378360
rect 210344 269074 210372 378354
rect 210332 269068 210384 269074
rect 210332 269010 210384 269016
rect 210240 57928 210292 57934
rect 210240 57870 210292 57876
rect 208860 57520 208912 57526
rect 208860 57462 208912 57468
rect 205548 57384 205600 57390
rect 205548 57326 205600 57332
rect 210436 57254 210464 469814
rect 210528 164966 210556 479538
rect 210700 472796 210752 472802
rect 210700 472738 210752 472744
rect 210608 468920 210660 468926
rect 210608 468862 210660 468868
rect 210620 166598 210648 468862
rect 210712 271017 210740 472738
rect 210792 471640 210844 471646
rect 210792 471582 210844 471588
rect 210804 272814 210832 471582
rect 210884 469124 210936 469130
rect 210884 469066 210936 469072
rect 210792 272808 210844 272814
rect 210792 272750 210844 272756
rect 210896 271386 210924 469066
rect 210976 466132 211028 466138
rect 210976 466074 211028 466080
rect 210988 273290 211016 466074
rect 211080 378842 211108 485454
rect 211160 485444 211212 485450
rect 211160 485386 211212 485392
rect 211172 485353 211200 485386
rect 211158 485344 211214 485353
rect 211158 485279 211214 485288
rect 211160 484832 211212 484838
rect 211158 484800 211160 484809
rect 211212 484800 211214 484809
rect 211158 484735 211214 484744
rect 211356 379234 211384 488022
rect 211620 484968 211672 484974
rect 211620 484910 211672 484916
rect 211528 468376 211580 468382
rect 211528 468318 211580 468324
rect 211344 379228 211396 379234
rect 211344 379170 211396 379176
rect 211080 378814 211200 378842
rect 211068 378752 211120 378758
rect 211068 378694 211120 378700
rect 211080 378350 211108 378694
rect 211068 378344 211120 378350
rect 211068 378286 211120 378292
rect 211172 378196 211200 378814
rect 211080 378168 211200 378196
rect 211080 374814 211108 378168
rect 211540 376242 211568 468318
rect 211632 377330 211660 484910
rect 211908 484430 211936 488022
rect 212092 485790 212120 488036
rect 212582 488022 212672 488050
rect 212080 485784 212132 485790
rect 212080 485726 212132 485732
rect 212540 485648 212592 485654
rect 212540 485590 212592 485596
rect 212552 485489 212580 485590
rect 212538 485480 212594 485489
rect 212538 485415 212594 485424
rect 212540 484492 212592 484498
rect 212540 484434 212592 484440
rect 211896 484424 211948 484430
rect 211896 484366 211948 484372
rect 211804 482656 211856 482662
rect 211804 482598 211856 482604
rect 211712 378344 211764 378350
rect 211712 378286 211764 378292
rect 211620 377324 211672 377330
rect 211620 377266 211672 377272
rect 211528 376236 211580 376242
rect 211528 376178 211580 376184
rect 211068 374808 211120 374814
rect 211068 374750 211120 374756
rect 210976 273284 211028 273290
rect 210976 273226 211028 273232
rect 210884 271380 210936 271386
rect 210884 271322 210936 271328
rect 210698 271008 210754 271017
rect 210698 270943 210754 270952
rect 211724 270502 211752 378286
rect 211712 270496 211764 270502
rect 211712 270438 211764 270444
rect 210974 269784 211030 269793
rect 210974 269719 211030 269728
rect 210884 269068 210936 269074
rect 210884 269010 210936 269016
rect 210896 268870 210924 269010
rect 210884 268864 210936 268870
rect 210884 268806 210936 268812
rect 210896 166802 210924 268806
rect 210884 166796 210936 166802
rect 210884 166738 210936 166744
rect 210608 166592 210660 166598
rect 210608 166534 210660 166540
rect 210516 164960 210568 164966
rect 210516 164902 210568 164908
rect 210988 147422 211016 269719
rect 211816 165034 211844 482598
rect 211896 475448 211948 475454
rect 211896 475390 211948 475396
rect 211908 165442 211936 475390
rect 212080 474020 212132 474026
rect 212080 473962 212132 473968
rect 211986 471336 212042 471345
rect 211986 471271 212042 471280
rect 211896 165436 211948 165442
rect 211896 165378 211948 165384
rect 211804 165028 211856 165034
rect 211804 164970 211856 164976
rect 212000 164218 212028 471271
rect 212092 271697 212120 473962
rect 212172 472660 212224 472666
rect 212172 472602 212224 472608
rect 212184 271794 212212 472602
rect 212264 467424 212316 467430
rect 212264 467366 212316 467372
rect 212276 272950 212304 467366
rect 212552 379778 212580 484434
rect 212644 484242 212672 488022
rect 212736 488022 213026 488050
rect 212736 484498 212764 488022
rect 212724 484492 212776 484498
rect 212724 484434 212776 484440
rect 213380 484430 213408 488036
rect 213472 488022 213854 488050
rect 214024 488022 214314 488050
rect 214790 488022 214880 488050
rect 212908 484424 212960 484430
rect 212908 484366 212960 484372
rect 213368 484424 213420 484430
rect 213368 484366 213420 484372
rect 212644 484214 212764 484242
rect 212632 484152 212684 484158
rect 212632 484094 212684 484100
rect 212540 379772 212592 379778
rect 212540 379714 212592 379720
rect 212448 379500 212500 379506
rect 212448 379442 212500 379448
rect 212356 379024 212408 379030
rect 212356 378966 212408 378972
rect 212264 272944 212316 272950
rect 212264 272886 212316 272892
rect 212172 271788 212224 271794
rect 212172 271730 212224 271736
rect 212078 271688 212134 271697
rect 212078 271623 212134 271632
rect 212368 271538 212396 378966
rect 212460 378350 212488 379442
rect 212448 378344 212500 378350
rect 212448 378286 212500 378292
rect 212446 378040 212502 378049
rect 212446 377975 212502 377984
rect 212276 271510 212396 271538
rect 212276 269686 212304 271510
rect 212356 270496 212408 270502
rect 212356 270438 212408 270444
rect 212368 270298 212396 270438
rect 212356 270292 212408 270298
rect 212356 270234 212408 270240
rect 212264 269680 212316 269686
rect 212264 269622 212316 269628
rect 212172 268456 212224 268462
rect 212172 268398 212224 268404
rect 211988 164212 212040 164218
rect 211988 164154 212040 164160
rect 212184 148442 212212 268398
rect 212172 148436 212224 148442
rect 212172 148378 212224 148384
rect 212276 147558 212304 269622
rect 212264 147552 212316 147558
rect 212264 147494 212316 147500
rect 210976 147416 211028 147422
rect 210976 147358 211028 147364
rect 212368 144702 212396 270234
rect 212356 144696 212408 144702
rect 212356 144638 212408 144644
rect 212460 58954 212488 377975
rect 212552 377806 212580 379714
rect 212644 379710 212672 484094
rect 212632 379704 212684 379710
rect 212632 379646 212684 379652
rect 212540 377800 212592 377806
rect 212540 377742 212592 377748
rect 212644 377738 212672 379646
rect 212736 379642 212764 484214
rect 212920 470594 212948 484366
rect 213472 484158 213500 488022
rect 213460 484152 213512 484158
rect 213460 484094 213512 484100
rect 213920 484152 213972 484158
rect 213920 484094 213972 484100
rect 213184 475584 213236 475590
rect 213184 475526 213236 475532
rect 212828 470566 212948 470594
rect 212724 379636 212776 379642
rect 212724 379578 212776 379584
rect 212632 377732 212684 377738
rect 212632 377674 212684 377680
rect 212736 376514 212764 379578
rect 212828 379438 212856 470566
rect 212908 467220 212960 467226
rect 212908 467162 212960 467168
rect 212920 381546 212948 467162
rect 213092 466404 213144 466410
rect 213092 466346 213144 466352
rect 212908 381540 212960 381546
rect 212908 381482 212960 381488
rect 212816 379432 212868 379438
rect 212816 379374 212868 379380
rect 213000 378276 213052 378282
rect 213000 378218 213052 378224
rect 213012 377194 213040 378218
rect 213000 377188 213052 377194
rect 213000 377130 213052 377136
rect 212724 376508 212776 376514
rect 212724 376450 212776 376456
rect 213104 376446 213132 466346
rect 213092 376440 213144 376446
rect 213092 376382 213144 376388
rect 213196 271862 213224 475526
rect 213460 471980 213512 471986
rect 213460 471922 213512 471928
rect 213368 378480 213420 378486
rect 213368 378422 213420 378428
rect 213276 377800 213328 377806
rect 213276 377742 213328 377748
rect 213184 271856 213236 271862
rect 213184 271798 213236 271804
rect 213182 271552 213238 271561
rect 213182 271487 213238 271496
rect 213092 270496 213144 270502
rect 213092 270438 213144 270444
rect 213104 144770 213132 270438
rect 213196 164082 213224 271487
rect 213288 269074 213316 377742
rect 213276 269068 213328 269074
rect 213276 269010 213328 269016
rect 213380 267714 213408 378422
rect 213472 376310 213500 471922
rect 213826 380488 213882 380497
rect 213826 380423 213882 380432
rect 213644 380384 213696 380390
rect 213644 380326 213696 380332
rect 213552 380112 213604 380118
rect 213552 380054 213604 380060
rect 213564 377482 213592 380054
rect 213656 378282 213684 380326
rect 213840 380118 213868 380423
rect 213828 380112 213880 380118
rect 213828 380054 213880 380060
rect 213828 379976 213880 379982
rect 213828 379918 213880 379924
rect 213840 379574 213868 379918
rect 213828 379568 213880 379574
rect 213748 379516 213828 379522
rect 213748 379510 213880 379516
rect 213748 379494 213868 379510
rect 213644 378276 213696 378282
rect 213644 378218 213696 378224
rect 213564 377454 213684 377482
rect 213552 377188 213604 377194
rect 213552 377130 213604 377136
rect 213460 376304 213512 376310
rect 213460 376246 213512 376252
rect 213564 270502 213592 377130
rect 213656 271561 213684 377454
rect 213642 271552 213698 271561
rect 213642 271487 213698 271496
rect 213552 270496 213604 270502
rect 213552 270438 213604 270444
rect 213564 270094 213592 270438
rect 213552 270088 213604 270094
rect 213552 270030 213604 270036
rect 213550 269920 213606 269929
rect 213550 269855 213606 269864
rect 213460 268388 213512 268394
rect 213460 268330 213512 268336
rect 213368 267708 213420 267714
rect 213368 267650 213420 267656
rect 213184 164076 213236 164082
rect 213184 164018 213236 164024
rect 213380 151814 213408 267650
rect 213288 151786 213408 151814
rect 213288 149054 213316 151786
rect 213276 149048 213328 149054
rect 213276 148990 213328 148996
rect 213184 147620 213236 147626
rect 213184 147562 213236 147568
rect 213092 144764 213144 144770
rect 213092 144706 213144 144712
rect 212448 58948 212500 58954
rect 212448 58890 212500 58896
rect 210424 57248 210476 57254
rect 210424 57190 210476 57196
rect 213196 55758 213224 147562
rect 213288 147490 213316 148990
rect 213472 148986 213500 268330
rect 213460 148980 213512 148986
rect 213460 148922 213512 148928
rect 213368 147688 213420 147694
rect 213368 147630 213420 147636
rect 213276 147484 213328 147490
rect 213276 147426 213328 147432
rect 213274 145752 213330 145761
rect 213274 145687 213330 145696
rect 213288 144906 213316 145687
rect 213276 144900 213328 144906
rect 213276 144842 213328 144848
rect 213184 55752 213236 55758
rect 213184 55694 213236 55700
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 162858 55040 162914 55049
rect 162858 54975 162914 54984
rect 160098 54904 160154 54913
rect 160098 54839 160154 54848
rect 122840 54528 122892 54534
rect 122840 54470 122892 54476
rect 213288 54330 213316 144842
rect 213380 56370 213408 147630
rect 213368 56364 213420 56370
rect 213368 56306 213420 56312
rect 213472 54398 213500 148922
rect 213564 148782 213592 269855
rect 213748 268666 213776 379494
rect 213828 379432 213880 379438
rect 213828 379374 213880 379380
rect 213840 378554 213868 379374
rect 213828 378548 213880 378554
rect 213828 378490 213880 378496
rect 213826 378040 213882 378049
rect 213826 377975 213882 377984
rect 213736 268660 213788 268666
rect 213736 268602 213788 268608
rect 213644 268524 213696 268530
rect 213644 268466 213696 268472
rect 213552 148776 213604 148782
rect 213552 148718 213604 148724
rect 213564 55894 213592 148718
rect 213656 144838 213684 268466
rect 213736 148572 213788 148578
rect 213736 148514 213788 148520
rect 213748 147626 213776 148514
rect 213736 147620 213788 147626
rect 213736 147562 213788 147568
rect 213736 147484 213788 147490
rect 213736 147426 213788 147432
rect 213644 144832 213696 144838
rect 213644 144774 213696 144780
rect 213552 55888 213604 55894
rect 213552 55830 213604 55836
rect 213748 55690 213776 147426
rect 213840 59022 213868 377975
rect 213932 375290 213960 484094
rect 214024 376378 214052 488022
rect 214748 485036 214800 485042
rect 214748 484978 214800 484984
rect 214564 483744 214616 483750
rect 214564 483686 214616 483692
rect 214380 468444 214432 468450
rect 214380 468386 214432 468392
rect 214288 464704 214340 464710
rect 214288 464646 214340 464652
rect 214196 378616 214248 378622
rect 214196 378558 214248 378564
rect 214012 376372 214064 376378
rect 214012 376314 214064 376320
rect 214024 376281 214052 376314
rect 214010 376272 214066 376281
rect 214010 376207 214066 376216
rect 213920 375284 213972 375290
rect 213920 375226 213972 375232
rect 214208 273358 214236 378558
rect 214300 376514 214328 464646
rect 214288 376508 214340 376514
rect 214288 376450 214340 376456
rect 214392 376174 214420 468386
rect 214470 376544 214526 376553
rect 214470 376479 214526 376488
rect 214380 376168 214432 376174
rect 214380 376110 214432 376116
rect 214484 375902 214512 376479
rect 214472 375896 214524 375902
rect 214472 375838 214524 375844
rect 214196 273352 214248 273358
rect 214196 273294 214248 273300
rect 214380 269544 214432 269550
rect 214380 269486 214432 269492
rect 214288 162852 214340 162858
rect 214288 162794 214340 162800
rect 214300 59226 214328 162794
rect 214392 144906 214420 269486
rect 214484 252550 214512 375838
rect 214472 252544 214524 252550
rect 214472 252486 214524 252492
rect 214484 162858 214512 252486
rect 214576 165510 214604 483686
rect 214760 480254 214788 484978
rect 214852 484537 214880 488022
rect 214944 488022 215234 488050
rect 215312 488022 215602 488050
rect 215680 488022 216062 488050
rect 216538 488022 216628 488050
rect 214838 484528 214894 484537
rect 214838 484463 214894 484472
rect 214944 484158 214972 488022
rect 214932 484152 214984 484158
rect 214932 484094 214984 484100
rect 214760 480226 214972 480254
rect 214656 471572 214708 471578
rect 214656 471514 214708 471520
rect 214668 166734 214696 471514
rect 214748 468852 214800 468858
rect 214748 468794 214800 468800
rect 214656 166728 214708 166734
rect 214656 166670 214708 166676
rect 214760 165578 214788 468794
rect 214840 465928 214892 465934
rect 214840 465870 214892 465876
rect 214852 270978 214880 465870
rect 214944 377738 214972 480226
rect 215312 384282 215340 488022
rect 215680 470594 215708 488022
rect 216600 484430 216628 488022
rect 216220 484424 216272 484430
rect 216220 484366 216272 484372
rect 216588 484424 216640 484430
rect 216588 484366 216640 484372
rect 215944 483676 215996 483682
rect 215944 483618 215996 483624
rect 215404 470566 215708 470594
rect 215404 389174 215432 470566
rect 215404 389146 215524 389174
rect 215312 384254 215432 384282
rect 215300 379840 215352 379846
rect 215300 379782 215352 379788
rect 215206 378040 215262 378049
rect 215206 377975 215262 377984
rect 214932 377732 214984 377738
rect 214932 377674 214984 377680
rect 215114 376680 215170 376689
rect 215114 376615 215170 376624
rect 215024 376032 215076 376038
rect 215024 375974 215076 375980
rect 214932 273352 214984 273358
rect 214932 273294 214984 273300
rect 214840 270972 214892 270978
rect 214840 270914 214892 270920
rect 214840 251864 214892 251870
rect 214840 251806 214892 251812
rect 214748 165572 214800 165578
rect 214748 165514 214800 165520
rect 214564 165504 214616 165510
rect 214564 165446 214616 165452
rect 214852 162858 214880 251806
rect 214472 162852 214524 162858
rect 214472 162794 214524 162800
rect 214840 162852 214892 162858
rect 214840 162794 214892 162800
rect 214852 161474 214880 162794
rect 214760 161446 214880 161474
rect 214656 148436 214708 148442
rect 214656 148378 214708 148384
rect 214564 147416 214616 147422
rect 214564 147358 214616 147364
rect 214470 145616 214526 145625
rect 214470 145551 214526 145560
rect 214380 144900 214432 144906
rect 214380 144842 214432 144848
rect 214484 144838 214512 145551
rect 214472 144832 214524 144838
rect 214472 144774 214524 144780
rect 214288 59220 214340 59226
rect 214288 59162 214340 59168
rect 213828 59016 213880 59022
rect 213828 58958 213880 58964
rect 213736 55684 213788 55690
rect 213736 55626 213788 55632
rect 214484 55185 214512 144774
rect 214470 55176 214526 55185
rect 214576 55146 214604 147358
rect 214668 56302 214696 148378
rect 214760 59158 214788 161446
rect 214944 148850 214972 273294
rect 215036 268938 215064 375974
rect 215024 268932 215076 268938
rect 215024 268874 215076 268880
rect 214932 148844 214984 148850
rect 214932 148786 214984 148792
rect 214944 147694 214972 148786
rect 215024 148504 215076 148510
rect 215024 148446 215076 148452
rect 214932 147688 214984 147694
rect 214932 147630 214984 147636
rect 215036 147422 215064 148446
rect 215024 147416 215076 147422
rect 215024 147358 215076 147364
rect 215024 146328 215076 146334
rect 215024 146270 215076 146276
rect 214932 145784 214984 145790
rect 214932 145726 214984 145732
rect 214748 59152 214800 59158
rect 214748 59094 214800 59100
rect 214656 56296 214708 56302
rect 214656 56238 214708 56244
rect 214470 55111 214526 55120
rect 214564 55140 214616 55146
rect 214564 55082 214616 55088
rect 214944 54602 214972 145726
rect 215036 56506 215064 146270
rect 215128 57730 215156 376615
rect 215116 57724 215168 57730
rect 215116 57666 215168 57672
rect 215220 57594 215248 377975
rect 215312 376038 215340 379782
rect 215300 376032 215352 376038
rect 215300 375974 215352 375980
rect 215404 375358 215432 384254
rect 215496 377913 215524 389146
rect 215852 380044 215904 380050
rect 215852 379986 215904 379992
rect 215482 377904 215538 377913
rect 215482 377839 215538 377848
rect 215760 377800 215812 377806
rect 215760 377742 215812 377748
rect 215392 375352 215444 375358
rect 215392 375294 215444 375300
rect 215772 269006 215800 377742
rect 215864 376718 215892 379986
rect 215852 376712 215904 376718
rect 215852 376654 215904 376660
rect 215864 271833 215892 376654
rect 215850 271824 215906 271833
rect 215850 271759 215906 271768
rect 215852 269476 215904 269482
rect 215852 269418 215904 269424
rect 215760 269000 215812 269006
rect 215760 268942 215812 268948
rect 215760 148368 215812 148374
rect 215760 148310 215812 148316
rect 215772 147558 215800 148310
rect 215760 147552 215812 147558
rect 215760 147494 215812 147500
rect 215864 146130 215892 269418
rect 215956 165102 215984 483618
rect 216128 474292 216180 474298
rect 216128 474234 216180 474240
rect 216034 465760 216090 465769
rect 216034 465695 216090 465704
rect 216048 165238 216076 465695
rect 216140 271590 216168 474234
rect 216232 379846 216260 484366
rect 216772 484152 216824 484158
rect 216772 484094 216824 484100
rect 216404 471776 216456 471782
rect 216404 471718 216456 471724
rect 216220 379840 216272 379846
rect 216220 379782 216272 379788
rect 216310 379264 216366 379273
rect 216310 379199 216366 379208
rect 216218 271824 216274 271833
rect 216218 271759 216274 271768
rect 216128 271584 216180 271590
rect 216128 271526 216180 271532
rect 216232 271289 216260 271759
rect 216218 271280 216274 271289
rect 216218 271215 216274 271224
rect 216128 269068 216180 269074
rect 216128 269010 216180 269016
rect 216140 268734 216168 269010
rect 216128 268728 216180 268734
rect 216128 268670 216180 268676
rect 216036 165232 216088 165238
rect 216036 165174 216088 165180
rect 215944 165096 215996 165102
rect 215944 165038 215996 165044
rect 216140 161634 216168 268670
rect 216232 164014 216260 271215
rect 216324 267646 216352 379199
rect 216416 375902 216444 471718
rect 216496 469192 216548 469198
rect 216496 469134 216548 469140
rect 216508 376378 216536 469134
rect 216678 417888 216734 417897
rect 216678 417823 216734 417832
rect 216692 417450 216720 417823
rect 216680 417444 216732 417450
rect 216680 417386 216732 417392
rect 216784 414730 216812 484094
rect 216772 414724 216824 414730
rect 216772 414666 216824 414672
rect 216862 413808 216918 413817
rect 216862 413743 216918 413752
rect 216876 413302 216904 413743
rect 216864 413296 216916 413302
rect 216864 413238 216916 413244
rect 216678 410952 216734 410961
rect 216678 410887 216734 410896
rect 216692 410582 216720 410887
rect 216680 410576 216732 410582
rect 216680 410518 216732 410524
rect 216692 409306 216720 410518
rect 216692 409278 216812 409306
rect 216678 409184 216734 409193
rect 216678 409119 216680 409128
rect 216732 409119 216734 409128
rect 216680 409090 216732 409096
rect 216680 391944 216732 391950
rect 216680 391886 216732 391892
rect 216692 390969 216720 391886
rect 216678 390960 216734 390969
rect 216678 390895 216734 390904
rect 216680 389836 216732 389842
rect 216680 389778 216732 389784
rect 216692 389337 216720 389778
rect 216678 389328 216734 389337
rect 216678 389263 216734 389272
rect 216678 380896 216734 380905
rect 216678 380831 216734 380840
rect 216692 380497 216720 380831
rect 216678 380488 216734 380497
rect 216678 380423 216734 380432
rect 216784 377262 216812 409278
rect 216876 380798 216904 413238
rect 216968 410718 216996 488036
rect 217428 485518 217456 488036
rect 217520 488022 217810 488050
rect 218164 488022 218270 488050
rect 218348 488022 218730 488050
rect 217416 485512 217468 485518
rect 217416 485454 217468 485460
rect 217416 485104 217468 485110
rect 217416 485046 217468 485052
rect 217324 478168 217376 478174
rect 217324 478110 217376 478116
rect 217232 474088 217284 474094
rect 217232 474030 217284 474036
rect 217244 416945 217272 474030
rect 217230 416936 217286 416945
rect 217230 416871 217286 416880
rect 217140 414860 217192 414866
rect 217140 414802 217192 414808
rect 217152 414769 217180 414802
rect 217138 414760 217194 414769
rect 217138 414695 217194 414704
rect 216956 410712 217008 410718
rect 216956 410654 217008 410660
rect 216954 409184 217010 409193
rect 216954 409119 217010 409128
rect 216968 380905 216996 409119
rect 216954 380896 217010 380905
rect 216954 380831 217010 380840
rect 216864 380792 216916 380798
rect 216864 380734 216916 380740
rect 216968 380633 216996 380831
rect 217152 380633 217180 414695
rect 217244 380866 217272 416871
rect 217336 412049 217364 478110
rect 217322 412040 217378 412049
rect 217322 411975 217378 411984
rect 217336 411369 217364 411975
rect 217322 411360 217378 411369
rect 217322 411295 217378 411304
rect 217322 380896 217378 380905
rect 217232 380860 217284 380866
rect 217322 380831 217378 380840
rect 217232 380802 217284 380808
rect 216954 380624 217010 380633
rect 216954 380559 217010 380568
rect 217138 380624 217194 380633
rect 217138 380559 217194 380568
rect 217244 379514 217272 380802
rect 217060 379486 217272 379514
rect 216772 377256 216824 377262
rect 216772 377198 216824 377204
rect 216956 377256 217008 377262
rect 216956 377198 217008 377204
rect 216496 376372 216548 376378
rect 216496 376314 216548 376320
rect 216404 375896 216456 375902
rect 216404 375838 216456 375844
rect 216586 375456 216642 375465
rect 216586 375391 216642 375400
rect 216496 375284 216548 375290
rect 216496 375226 216548 375232
rect 216404 375012 216456 375018
rect 216404 374954 216456 374960
rect 216416 269074 216444 374954
rect 216508 374950 216536 375226
rect 216496 374944 216548 374950
rect 216496 374886 216548 374892
rect 216404 269068 216456 269074
rect 216404 269010 216456 269016
rect 216508 268802 216536 374886
rect 216496 268796 216548 268802
rect 216496 268738 216548 268744
rect 216496 268660 216548 268666
rect 216496 268602 216548 268608
rect 216508 268326 216536 268602
rect 216496 268320 216548 268326
rect 216496 268262 216548 268268
rect 216312 267640 216364 267646
rect 216312 267582 216364 267588
rect 216220 164008 216272 164014
rect 216220 163950 216272 163956
rect 216128 161628 216180 161634
rect 216128 161570 216180 161576
rect 216140 161474 216168 161570
rect 216140 161446 216260 161474
rect 215944 147552 215996 147558
rect 215944 147494 215996 147500
rect 215852 146124 215904 146130
rect 215852 146066 215904 146072
rect 215850 146024 215906 146033
rect 215850 145959 215906 145968
rect 215864 59430 215892 145959
rect 215852 59424 215904 59430
rect 215852 59366 215904 59372
rect 215208 57588 215260 57594
rect 215208 57530 215260 57536
rect 215024 56500 215076 56506
rect 215024 56442 215076 56448
rect 215956 55078 215984 147494
rect 216128 145920 216180 145926
rect 216128 145862 216180 145868
rect 216036 145648 216088 145654
rect 216036 145590 216088 145596
rect 216048 144770 216076 145590
rect 216036 144764 216088 144770
rect 216036 144706 216088 144712
rect 216048 55826 216076 144706
rect 216036 55820 216088 55826
rect 216036 55762 216088 55768
rect 215944 55072 215996 55078
rect 215944 55014 215996 55020
rect 216140 54670 216168 145862
rect 216232 59566 216260 161446
rect 216324 148918 216352 267582
rect 216508 258074 216536 268262
rect 216416 258046 216536 258074
rect 216312 148912 216364 148918
rect 216312 148854 216364 148860
rect 216220 59560 216272 59566
rect 216220 59502 216272 59508
rect 216128 54664 216180 54670
rect 216128 54606 216180 54612
rect 214932 54596 214984 54602
rect 214932 54538 214984 54544
rect 216324 54466 216352 148854
rect 216416 145858 216444 258046
rect 216496 146056 216548 146062
rect 216496 145998 216548 146004
rect 216404 145852 216456 145858
rect 216404 145794 216456 145800
rect 216416 55214 216444 145794
rect 216404 55208 216456 55214
rect 216404 55150 216456 55156
rect 216508 54738 216536 145998
rect 216600 57662 216628 375391
rect 216862 310040 216918 310049
rect 216862 309975 216918 309984
rect 216680 284300 216732 284306
rect 216680 284242 216732 284248
rect 216692 284073 216720 284242
rect 216678 284064 216734 284073
rect 216678 283999 216734 284008
rect 216772 282872 216824 282878
rect 216772 282814 216824 282820
rect 216678 282296 216734 282305
rect 216678 282231 216734 282240
rect 216692 282198 216720 282231
rect 216680 282192 216732 282198
rect 216784 282169 216812 282814
rect 216680 282134 216732 282140
rect 216770 282160 216826 282169
rect 216770 282095 216826 282104
rect 216772 270156 216824 270162
rect 216772 270098 216824 270104
rect 216680 269612 216732 269618
rect 216680 269554 216732 269560
rect 216692 176746 216720 269554
rect 216784 178106 216812 270098
rect 216876 203017 216904 309975
rect 216968 303929 216996 377198
rect 217060 310049 217088 379486
rect 217232 375352 217284 375358
rect 217232 375294 217284 375300
rect 217244 374882 217272 375294
rect 217232 374876 217284 374882
rect 217232 374818 217284 374824
rect 217140 358284 217192 358290
rect 217140 358226 217192 358232
rect 217046 310040 217102 310049
rect 217046 309975 217102 309984
rect 216954 303920 217010 303929
rect 216954 303855 217010 303864
rect 216954 302152 217010 302161
rect 216954 302087 217010 302096
rect 216862 203008 216918 203017
rect 216862 202943 216918 202952
rect 216862 198792 216918 198801
rect 216862 198727 216918 198736
rect 216876 178226 216904 198727
rect 216968 195265 216996 302087
rect 217152 269822 217180 358226
rect 217140 269816 217192 269822
rect 217140 269758 217192 269764
rect 217244 269278 217272 374818
rect 217336 302161 217364 380831
rect 217428 377806 217456 485046
rect 217520 484158 217548 488022
rect 217508 484152 217560 484158
rect 217508 484094 217560 484100
rect 217692 471844 217744 471850
rect 217692 471786 217744 471792
rect 217508 471708 217560 471714
rect 217508 471650 217560 471656
rect 217416 377800 217468 377806
rect 217416 377742 217468 377748
rect 217520 375834 217548 471650
rect 217600 466268 217652 466274
rect 217600 466210 217652 466216
rect 217612 380934 217640 466210
rect 217704 410106 217732 471786
rect 218060 467288 218112 467294
rect 218060 467230 218112 467236
rect 218072 466546 218100 467230
rect 218060 466540 218112 466546
rect 218060 466482 218112 466488
rect 217874 417888 217930 417897
rect 217874 417823 217930 417832
rect 217782 411360 217838 411369
rect 217782 411295 217838 411304
rect 217692 410100 217744 410106
rect 217692 410042 217744 410048
rect 217692 389156 217744 389162
rect 217692 389098 217744 389104
rect 217704 389065 217732 389098
rect 217690 389056 217746 389065
rect 217690 388991 217746 389000
rect 217600 380928 217652 380934
rect 217600 380870 217652 380876
rect 217692 380792 217744 380798
rect 217692 380734 217744 380740
rect 217598 380624 217654 380633
rect 217598 380559 217654 380568
rect 217612 380089 217640 380559
rect 217598 380080 217654 380089
rect 217598 380015 217654 380024
rect 217508 375828 217560 375834
rect 217508 375770 217560 375776
rect 217612 307873 217640 380015
rect 217598 307864 217654 307873
rect 217598 307799 217654 307808
rect 217506 303920 217562 303929
rect 217506 303855 217562 303864
rect 217322 302152 217378 302161
rect 217322 302087 217378 302096
rect 217232 269272 217284 269278
rect 217232 269214 217284 269220
rect 217140 268932 217192 268938
rect 217140 268874 217192 268880
rect 217152 268666 217180 268874
rect 217140 268660 217192 268666
rect 217140 268602 217192 268608
rect 216954 195256 217010 195265
rect 216954 195191 217010 195200
rect 216864 178220 216916 178226
rect 216864 178162 216916 178168
rect 216784 178078 216996 178106
rect 216772 178016 216824 178022
rect 216772 177958 216824 177964
rect 216864 178016 216916 178022
rect 216864 177958 216916 177964
rect 216784 177041 216812 177958
rect 216770 177032 216826 177041
rect 216770 176967 216826 176976
rect 216692 176718 216812 176746
rect 216680 176656 216732 176662
rect 216680 176598 216732 176604
rect 216692 175409 216720 176598
rect 216678 175400 216734 175409
rect 216678 175335 216734 175344
rect 216784 175250 216812 176718
rect 216692 175222 216812 175250
rect 216692 163538 216720 175222
rect 216772 175160 216824 175166
rect 216772 175102 216824 175108
rect 216680 163532 216732 163538
rect 216680 163474 216732 163480
rect 216784 145314 216812 175102
rect 216772 145308 216824 145314
rect 216772 145250 216824 145256
rect 216876 92857 216904 177958
rect 216968 175166 216996 178078
rect 217048 175228 217100 175234
rect 217048 175170 217100 175176
rect 216956 175160 217008 175166
rect 217060 175137 217088 175170
rect 216956 175102 217008 175108
rect 217046 175128 217102 175137
rect 217046 175063 217102 175072
rect 217152 161498 217180 268602
rect 217414 203960 217470 203969
rect 217414 203895 217470 203904
rect 217140 161492 217192 161498
rect 216968 161446 217140 161474
rect 216862 92848 216918 92857
rect 216862 92783 216918 92792
rect 216680 70372 216732 70378
rect 216680 70314 216732 70320
rect 216692 70009 216720 70314
rect 216678 70000 216734 70009
rect 216678 69935 216734 69944
rect 216678 68368 216734 68377
rect 216678 68303 216734 68312
rect 216692 67658 216720 68303
rect 216680 67652 216732 67658
rect 216680 67594 216732 67600
rect 216968 59634 216996 161446
rect 217140 161434 217192 161440
rect 217322 146296 217378 146305
rect 217322 146231 217378 146240
rect 217336 145926 217364 146231
rect 217324 145920 217376 145926
rect 217324 145862 217376 145868
rect 217048 145580 217100 145586
rect 217048 145522 217100 145528
rect 217060 144906 217088 145522
rect 217232 145308 217284 145314
rect 217232 145250 217284 145256
rect 217048 144900 217100 144906
rect 217048 144842 217100 144848
rect 217060 142154 217088 144842
rect 217060 142126 217180 142154
rect 216956 59628 217008 59634
rect 216956 59570 217008 59576
rect 216588 57656 216640 57662
rect 216588 57598 216640 57604
rect 217152 55962 217180 142126
rect 217140 55956 217192 55962
rect 217140 55898 217192 55904
rect 217244 54806 217272 145250
rect 217428 96937 217456 203895
rect 217520 197033 217548 303855
rect 217612 200841 217640 307799
rect 217704 306785 217732 380734
rect 217796 380497 217824 411295
rect 217782 380488 217838 380497
rect 217782 380423 217838 380432
rect 217690 306776 217746 306785
rect 217690 306711 217746 306720
rect 217598 200832 217654 200841
rect 217598 200767 217654 200776
rect 217506 197024 217562 197033
rect 217506 196959 217562 196968
rect 217414 96928 217470 96937
rect 217414 96863 217470 96872
rect 217520 90001 217548 196959
rect 217612 93809 217640 200767
rect 217704 199889 217732 306711
rect 217796 305017 217824 380423
rect 217888 311001 217916 417823
rect 218164 378593 218192 488022
rect 218244 466540 218296 466546
rect 218244 466482 218296 466488
rect 218256 381070 218284 466482
rect 218244 381064 218296 381070
rect 218244 381006 218296 381012
rect 218348 379302 218376 488022
rect 219176 485178 219204 488036
rect 219574 488022 219664 488050
rect 219164 485172 219216 485178
rect 219164 485114 219216 485120
rect 219164 484424 219216 484430
rect 219164 484366 219216 484372
rect 218796 476808 218848 476814
rect 218796 476750 218848 476756
rect 218704 467152 218756 467158
rect 218704 467094 218756 467100
rect 218336 379296 218388 379302
rect 218336 379238 218388 379244
rect 218150 378584 218206 378593
rect 218150 378519 218206 378528
rect 217966 377904 218022 377913
rect 217966 377839 218022 377848
rect 217874 310992 217930 311001
rect 217874 310927 217930 310936
rect 217782 305008 217838 305017
rect 217782 304943 217838 304952
rect 217690 199880 217746 199889
rect 217690 199815 217746 199824
rect 217704 198801 217732 199815
rect 217690 198792 217746 198801
rect 217690 198727 217746 198736
rect 217796 198121 217824 304943
rect 217888 203969 217916 310927
rect 217980 269618 218008 377839
rect 218520 375692 218572 375698
rect 218520 375634 218572 375640
rect 218426 273456 218482 273465
rect 218426 273391 218482 273400
rect 217968 269612 218020 269618
rect 217968 269554 218020 269560
rect 217966 252512 218022 252521
rect 217966 252447 217968 252456
rect 218020 252447 218022 252456
rect 217968 252418 218020 252424
rect 217874 203960 217930 203969
rect 217874 203895 217930 203904
rect 217874 203008 217930 203017
rect 217874 202943 217930 202952
rect 217782 198112 217838 198121
rect 217782 198047 217838 198056
rect 217690 195256 217746 195265
rect 217690 195191 217746 195200
rect 217598 93800 217654 93809
rect 217598 93735 217654 93744
rect 217506 89992 217562 90001
rect 217506 89927 217562 89936
rect 217704 88233 217732 195191
rect 217796 91089 217824 198047
rect 217888 95985 217916 202943
rect 217966 162752 218022 162761
rect 217966 162687 217968 162696
rect 218020 162687 218022 162696
rect 217968 162658 218020 162664
rect 218242 146296 218298 146305
rect 218242 146231 218298 146240
rect 218060 145716 218112 145722
rect 218060 145658 218112 145664
rect 218072 144702 218100 145658
rect 218060 144696 218112 144702
rect 218060 144638 218112 144644
rect 217874 95976 217930 95985
rect 217874 95911 217930 95920
rect 217782 91080 217838 91089
rect 217782 91015 217838 91024
rect 217690 88224 217746 88233
rect 217690 88159 217746 88168
rect 217966 68368 218022 68377
rect 217966 68303 218022 68312
rect 217980 59362 218008 68303
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218256 56166 218284 146231
rect 218440 57458 218468 273391
rect 218532 269414 218560 375634
rect 218612 358692 218664 358698
rect 218612 358634 218664 358640
rect 218624 270366 218652 358634
rect 218612 270360 218664 270366
rect 218612 270302 218664 270308
rect 218612 269816 218664 269822
rect 218612 269758 218664 269764
rect 218520 269408 218572 269414
rect 218520 269350 218572 269356
rect 218520 269000 218572 269006
rect 218520 268942 218572 268948
rect 218532 268598 218560 268942
rect 218520 268592 218572 268598
rect 218520 268534 218572 268540
rect 218532 162654 218560 268534
rect 218520 162648 218572 162654
rect 218520 162590 218572 162596
rect 218624 162178 218652 269758
rect 218612 162172 218664 162178
rect 218612 162114 218664 162120
rect 218520 145512 218572 145518
rect 218520 145454 218572 145460
rect 218532 59702 218560 145454
rect 218612 145444 218664 145450
rect 218612 145386 218664 145392
rect 218624 61266 218652 145386
rect 218612 61260 218664 61266
rect 218612 61202 218664 61208
rect 218716 61146 218744 467094
rect 218808 165374 218836 476750
rect 218888 474224 218940 474230
rect 218888 474166 218940 474172
rect 218796 165368 218848 165374
rect 218796 165310 218848 165316
rect 218900 164898 218928 474166
rect 218980 469940 219032 469946
rect 218980 469882 219032 469888
rect 218992 165170 219020 469882
rect 219072 465996 219124 466002
rect 219072 465938 219124 465944
rect 219084 271454 219112 465938
rect 219176 380866 219204 484366
rect 219532 484220 219584 484226
rect 219532 484162 219584 484168
rect 219440 484152 219492 484158
rect 219440 484094 219492 484100
rect 219256 410100 219308 410106
rect 219256 410042 219308 410048
rect 219164 380860 219216 380866
rect 219164 380802 219216 380808
rect 219268 376038 219296 410042
rect 219348 380860 219400 380866
rect 219348 380802 219400 380808
rect 219360 379506 219388 380802
rect 219348 379500 219400 379506
rect 219348 379442 219400 379448
rect 219256 376032 219308 376038
rect 219256 375974 219308 375980
rect 219360 375698 219388 379442
rect 219452 379438 219480 484094
rect 219544 381002 219572 484162
rect 219532 380996 219584 381002
rect 219532 380938 219584 380944
rect 219440 379432 219492 379438
rect 219440 379374 219492 379380
rect 219452 378894 219480 379374
rect 219636 379370 219664 488022
rect 219728 488022 220018 488050
rect 220096 488022 220478 488050
rect 220832 488022 220938 488050
rect 221016 488022 221398 488050
rect 219728 484158 219756 488022
rect 219900 485240 219952 485246
rect 219900 485182 219952 485188
rect 219716 484152 219768 484158
rect 219716 484094 219768 484100
rect 219912 380866 219940 485182
rect 219992 484424 220044 484430
rect 219992 484366 220044 484372
rect 219900 380860 219952 380866
rect 219900 380802 219952 380808
rect 219808 379908 219860 379914
rect 219808 379850 219860 379856
rect 219820 379642 219848 379850
rect 219808 379636 219860 379642
rect 219808 379578 219860 379584
rect 219900 379636 219952 379642
rect 219900 379578 219952 379584
rect 219624 379364 219676 379370
rect 219624 379306 219676 379312
rect 219532 379228 219584 379234
rect 219532 379170 219584 379176
rect 219440 378888 219492 378894
rect 219440 378830 219492 378836
rect 219348 375692 219400 375698
rect 219348 375634 219400 375640
rect 219440 374808 219492 374814
rect 219440 374750 219492 374756
rect 219348 374740 219400 374746
rect 219348 374682 219400 374688
rect 219256 358760 219308 358766
rect 219256 358702 219308 358708
rect 219164 357876 219216 357882
rect 219164 357818 219216 357824
rect 219072 271448 219124 271454
rect 219072 271390 219124 271396
rect 219176 270230 219204 357818
rect 219164 270224 219216 270230
rect 219164 270166 219216 270172
rect 219072 269068 219124 269074
rect 219072 269010 219124 269016
rect 219084 268258 219112 269010
rect 219072 268252 219124 268258
rect 219072 268194 219124 268200
rect 218980 165164 219032 165170
rect 218980 165106 219032 165112
rect 218888 164892 218940 164898
rect 218888 164834 218940 164840
rect 218980 163532 219032 163538
rect 218980 163474 219032 163480
rect 218888 162648 218940 162654
rect 218888 162590 218940 162596
rect 218796 144696 218848 144702
rect 218796 144638 218848 144644
rect 218624 61118 218744 61146
rect 218520 59696 218572 59702
rect 218520 59638 218572 59644
rect 218428 57452 218480 57458
rect 218428 57394 218480 57400
rect 218624 57322 218652 61118
rect 218702 60616 218758 60625
rect 218702 60551 218758 60560
rect 218716 57798 218744 60551
rect 218704 57792 218756 57798
rect 218704 57734 218756 57740
rect 218612 57316 218664 57322
rect 218612 57258 218664 57264
rect 218244 56160 218296 56166
rect 218244 56102 218296 56108
rect 217232 54800 217284 54806
rect 217232 54742 217284 54748
rect 216496 54732 216548 54738
rect 216496 54674 216548 54680
rect 218808 54534 218836 144638
rect 218900 59294 218928 162590
rect 218992 59498 219020 163474
rect 219084 145790 219112 268194
rect 219176 145994 219204 270166
rect 219268 270162 219296 358702
rect 219360 273426 219388 374682
rect 219452 358290 219480 374750
rect 219440 358284 219492 358290
rect 219440 358226 219492 358232
rect 219348 273420 219400 273426
rect 219348 273362 219400 273368
rect 219348 270360 219400 270366
rect 219348 270302 219400 270308
rect 219256 270156 219308 270162
rect 219256 270098 219308 270104
rect 219360 146130 219388 270302
rect 219544 269550 219572 379170
rect 219636 378622 219664 379306
rect 219716 378752 219768 378758
rect 219716 378694 219768 378700
rect 219624 378616 219676 378622
rect 219624 378558 219676 378564
rect 219624 378208 219676 378214
rect 219624 378150 219676 378156
rect 219636 270065 219664 378150
rect 219622 270056 219678 270065
rect 219622 269991 219678 270000
rect 219532 269544 219584 269550
rect 219532 269486 219584 269492
rect 219728 269482 219756 378694
rect 219716 269476 219768 269482
rect 219716 269418 219768 269424
rect 219624 269408 219676 269414
rect 219624 269350 219676 269356
rect 219440 269272 219492 269278
rect 219440 269214 219492 269220
rect 219348 146124 219400 146130
rect 219348 146066 219400 146072
rect 219164 145988 219216 145994
rect 219164 145930 219216 145936
rect 219072 145784 219124 145790
rect 219072 145726 219124 145732
rect 219072 61260 219124 61266
rect 219072 61202 219124 61208
rect 218980 59492 219032 59498
rect 218980 59434 219032 59440
rect 218888 59288 218940 59294
rect 218888 59230 218940 59236
rect 219084 56438 219112 61202
rect 219072 56432 219124 56438
rect 219072 56374 219124 56380
rect 219176 56030 219204 145930
rect 219360 142154 219388 146066
rect 219452 146033 219480 269214
rect 219636 164150 219664 269350
rect 219820 269006 219848 379578
rect 219912 377913 219940 379578
rect 219898 377904 219954 377913
rect 219898 377839 219954 377848
rect 219900 273420 219952 273426
rect 219900 273362 219952 273368
rect 219808 269000 219860 269006
rect 219808 268942 219860 268948
rect 219624 164144 219676 164150
rect 219624 164086 219676 164092
rect 219532 162172 219584 162178
rect 219532 162114 219584 162120
rect 219438 146024 219494 146033
rect 219438 145959 219494 145968
rect 219268 142126 219388 142154
rect 219268 74534 219296 142126
rect 219268 74506 219388 74534
rect 219254 60616 219310 60625
rect 219254 60551 219310 60560
rect 219268 58682 219296 60551
rect 219256 58676 219308 58682
rect 219256 58618 219308 58624
rect 219360 56098 219388 74506
rect 219348 56092 219400 56098
rect 219348 56034 219400 56040
rect 219164 56024 219216 56030
rect 219164 55966 219216 55972
rect 219544 55010 219572 162114
rect 219532 55004 219584 55010
rect 219532 54946 219584 54952
rect 219636 54942 219664 164086
rect 219820 145382 219848 268942
rect 219912 146305 219940 273362
rect 219898 146296 219954 146305
rect 219898 146231 219954 146240
rect 219898 146160 219954 146169
rect 219898 146095 219954 146104
rect 219808 145376 219860 145382
rect 219808 145318 219860 145324
rect 219624 54936 219676 54942
rect 219624 54878 219676 54884
rect 219820 54874 219848 145318
rect 219912 56234 219940 146095
rect 220004 56574 220032 484366
rect 220096 484226 220124 488022
rect 220084 484220 220136 484226
rect 220084 484162 220136 484168
rect 220832 480282 220860 488022
rect 221016 484242 221044 488022
rect 221752 485382 221780 488036
rect 222242 488022 222608 488050
rect 221740 485376 221792 485382
rect 221740 485318 221792 485324
rect 220924 484214 221044 484242
rect 220820 480276 220872 480282
rect 220820 480218 220872 480224
rect 220924 465730 220952 484214
rect 222580 482322 222608 488022
rect 222672 484430 222700 488036
rect 223162 488022 223528 488050
rect 223622 488022 223712 488050
rect 223990 488022 224080 488050
rect 223500 485110 223528 488022
rect 223488 485104 223540 485110
rect 223488 485046 223540 485052
rect 222660 484424 222712 484430
rect 222660 484366 222712 484372
rect 223580 484152 223632 484158
rect 223580 484094 223632 484100
rect 222568 482316 222620 482322
rect 222568 482258 222620 482264
rect 221004 480276 221056 480282
rect 221004 480218 221056 480224
rect 221016 465798 221044 480218
rect 223592 474065 223620 484094
rect 223684 479641 223712 488022
rect 224052 485246 224080 488022
rect 224144 488022 224434 488050
rect 224040 485240 224092 485246
rect 224040 485182 224092 485188
rect 224144 484158 224172 488022
rect 224880 484537 224908 488036
rect 225370 488022 225644 488050
rect 225738 488022 226104 488050
rect 225616 485382 225644 488022
rect 226076 485518 226104 488022
rect 226064 485512 226116 485518
rect 226064 485454 226116 485460
rect 225604 485376 225656 485382
rect 225604 485318 225656 485324
rect 226168 485081 226196 488036
rect 226154 485072 226210 485081
rect 226154 485007 226210 485016
rect 224866 484528 224922 484537
rect 224866 484463 224922 484472
rect 224132 484152 224184 484158
rect 224132 484094 224184 484100
rect 226340 484152 226392 484158
rect 226340 484094 226392 484100
rect 223670 479632 223726 479641
rect 223670 479567 223726 479576
rect 223578 474056 223634 474065
rect 223578 473991 223634 474000
rect 226352 472705 226380 484094
rect 226432 484016 226484 484022
rect 226432 483958 226484 483964
rect 226444 472734 226472 483958
rect 226628 475454 226656 488036
rect 226720 488022 227102 488050
rect 227272 488022 227562 488050
rect 227732 488022 227930 488050
rect 228406 488022 228496 488050
rect 226720 484158 226748 488022
rect 226708 484152 226760 484158
rect 226708 484094 226760 484100
rect 227272 484022 227300 488022
rect 227260 484016 227312 484022
rect 227260 483958 227312 483964
rect 226616 475448 226668 475454
rect 226616 475390 226668 475396
rect 226432 472728 226484 472734
rect 226338 472696 226394 472705
rect 226432 472670 226484 472676
rect 227732 472666 227760 488022
rect 228468 483857 228496 488022
rect 228560 488022 228850 488050
rect 229204 488022 229310 488050
rect 229480 488022 229770 488050
rect 229848 488022 230138 488050
rect 230614 488022 230888 488050
rect 231074 488022 231440 488050
rect 231534 488022 231808 488050
rect 231902 488022 232176 488050
rect 228454 483848 228510 483857
rect 228454 483783 228510 483792
rect 228560 478281 228588 488022
rect 229100 484152 229152 484158
rect 229100 484094 229152 484100
rect 228546 478272 228602 478281
rect 228546 478207 228602 478216
rect 226338 472631 226394 472640
rect 227720 472660 227772 472666
rect 227720 472602 227772 472608
rect 229112 472569 229140 484094
rect 229204 474026 229232 488022
rect 229480 484158 229508 488022
rect 229468 484152 229520 484158
rect 229468 484094 229520 484100
rect 229848 474094 229876 488022
rect 230860 485450 230888 488022
rect 230848 485444 230900 485450
rect 230848 485386 230900 485392
rect 231412 483721 231440 488022
rect 231780 485178 231808 488022
rect 231768 485172 231820 485178
rect 231768 485114 231820 485120
rect 231398 483712 231454 483721
rect 231398 483647 231454 483656
rect 232148 480865 232176 488022
rect 232332 485081 232360 488036
rect 232424 488022 232806 488050
rect 232318 485072 232374 485081
rect 232318 485007 232374 485016
rect 232134 480856 232190 480865
rect 232134 480791 232190 480800
rect 232424 475561 232452 488022
rect 233252 485489 233280 488036
rect 233344 488022 233726 488050
rect 234110 488022 234384 488050
rect 233238 485480 233294 485489
rect 233238 485415 233294 485424
rect 233344 478174 233372 488022
rect 234356 485217 234384 488022
rect 234540 485722 234568 488036
rect 234632 488022 235014 488050
rect 235490 488022 235856 488050
rect 234528 485716 234580 485722
rect 234528 485658 234580 485664
rect 234342 485208 234398 485217
rect 234342 485143 234398 485152
rect 233332 478168 233384 478174
rect 233332 478110 233384 478116
rect 234632 476785 234660 488022
rect 235828 485625 235856 488022
rect 235814 485616 235870 485625
rect 235814 485551 235870 485560
rect 235920 485353 235948 488036
rect 236318 488022 236592 488050
rect 235906 485344 235962 485353
rect 235906 485279 235962 485288
rect 236564 482361 236592 488022
rect 236748 483750 236776 488036
rect 236840 488022 237222 488050
rect 237392 488022 237682 488050
rect 237760 488022 238142 488050
rect 238220 488022 238510 488050
rect 238772 488022 238970 488050
rect 239446 488022 239720 488050
rect 239906 488022 240088 488050
rect 236736 483744 236788 483750
rect 236736 483686 236788 483692
rect 236550 482352 236606 482361
rect 236550 482287 236606 482296
rect 236840 476882 236868 488022
rect 237392 476950 237420 488022
rect 237760 484106 237788 488022
rect 237484 484078 237788 484106
rect 237484 478242 237512 484078
rect 238220 479534 238248 488022
rect 238208 479528 238260 479534
rect 238208 479470 238260 479476
rect 237472 478236 237524 478242
rect 237472 478178 237524 478184
rect 237380 476944 237432 476950
rect 237380 476886 237432 476892
rect 236828 476876 236880 476882
rect 236828 476818 236880 476824
rect 234618 476776 234674 476785
rect 234618 476711 234674 476720
rect 232410 475552 232466 475561
rect 232410 475487 232466 475496
rect 238772 475386 238800 488022
rect 239692 485654 239720 488022
rect 239680 485648 239732 485654
rect 239680 485590 239732 485596
rect 240060 485314 240088 488022
rect 240152 488022 240258 488050
rect 240336 488022 240718 488050
rect 240888 488022 241178 488050
rect 240048 485308 240100 485314
rect 240048 485250 240100 485256
rect 238760 475380 238812 475386
rect 238760 475322 238812 475328
rect 229836 474088 229888 474094
rect 229836 474030 229888 474036
rect 229192 474020 229244 474026
rect 229192 473962 229244 473968
rect 229098 472560 229154 472569
rect 229098 472495 229154 472504
rect 240152 471374 240180 488022
rect 240232 484152 240284 484158
rect 240232 484094 240284 484100
rect 240140 471368 240192 471374
rect 240140 471310 240192 471316
rect 240244 471306 240272 484094
rect 240336 478145 240364 488022
rect 240888 484158 240916 488022
rect 240876 484152 240928 484158
rect 240876 484094 240928 484100
rect 241520 484152 241572 484158
rect 241520 484094 241572 484100
rect 240322 478136 240378 478145
rect 240322 478071 240378 478080
rect 240232 471300 240284 471306
rect 240232 471242 240284 471248
rect 241532 465798 241560 484094
rect 241624 474230 241652 488036
rect 241716 488022 242098 488050
rect 242176 488022 242466 488050
rect 241716 478310 241744 488022
rect 242176 484158 242204 488022
rect 242928 487778 242956 488036
rect 243188 488022 243386 488050
rect 243464 488022 243846 488050
rect 244322 488022 244596 488050
rect 242928 487750 243124 487778
rect 242164 484152 242216 484158
rect 242164 484094 242216 484100
rect 243096 481098 243124 487750
rect 243084 481092 243136 481098
rect 243084 481034 243136 481040
rect 243188 480978 243216 488022
rect 242912 480950 243216 480978
rect 241704 478304 241756 478310
rect 241704 478246 241756 478252
rect 241612 474224 241664 474230
rect 241612 474166 241664 474172
rect 221004 465792 221056 465798
rect 221004 465734 221056 465740
rect 241520 465792 241572 465798
rect 241520 465734 241572 465740
rect 242912 465730 242940 480950
rect 243464 479670 243492 488022
rect 244568 485722 244596 488022
rect 244556 485716 244608 485722
rect 244556 485658 244608 485664
rect 244660 482458 244688 488036
rect 244752 488022 245134 488050
rect 245304 488022 245594 488050
rect 245672 488022 246054 488050
rect 246132 488022 246422 488050
rect 246898 488022 246988 488050
rect 244648 482452 244700 482458
rect 244648 482394 244700 482400
rect 243452 479664 243504 479670
rect 243452 479606 243504 479612
rect 244752 476114 244780 488022
rect 244292 476086 244780 476114
rect 244292 474162 244320 476086
rect 245304 475522 245332 488022
rect 245292 475516 245344 475522
rect 245292 475458 245344 475464
rect 244280 474156 244332 474162
rect 244280 474098 244332 474104
rect 245672 466070 245700 488022
rect 246132 479602 246160 488022
rect 246960 483682 246988 488022
rect 247052 488022 247342 488050
rect 247818 488022 248092 488050
rect 248278 488022 248368 488050
rect 246948 483676 247000 483682
rect 246948 483618 247000 483624
rect 246120 479596 246172 479602
rect 246120 479538 246172 479544
rect 247052 476814 247080 488022
rect 248064 481030 248092 488022
rect 248340 482390 248368 488022
rect 248524 488022 248630 488050
rect 248800 488022 249090 488050
rect 249168 488022 249550 488050
rect 249904 488022 250010 488050
rect 250088 488022 250470 488050
rect 250548 488022 250838 488050
rect 251314 488022 251404 488050
rect 248328 482384 248380 482390
rect 248328 482326 248380 482332
rect 248052 481024 248104 481030
rect 248052 480966 248104 480972
rect 248420 480888 248472 480894
rect 248420 480830 248472 480836
rect 247040 476808 247092 476814
rect 247040 476750 247092 476756
rect 245660 466064 245712 466070
rect 245660 466006 245712 466012
rect 248432 465769 248460 480830
rect 248524 465934 248552 488022
rect 248800 480894 248828 488022
rect 248788 480888 248840 480894
rect 248788 480830 248840 480836
rect 249168 470594 249196 488022
rect 249800 480888 249852 480894
rect 249800 480830 249852 480836
rect 248616 470566 249196 470594
rect 248512 465928 248564 465934
rect 248512 465870 248564 465876
rect 248616 465866 248644 470566
rect 249812 466138 249840 480830
rect 249800 466132 249852 466138
rect 249800 466074 249852 466080
rect 249904 466002 249932 488022
rect 250088 470594 250116 488022
rect 250548 480894 250576 488022
rect 251376 481166 251404 488022
rect 251468 488022 251758 488050
rect 251928 488022 252218 488050
rect 252602 488022 252692 488050
rect 251364 481160 251416 481166
rect 251364 481102 251416 481108
rect 250536 480888 250588 480894
rect 250536 480830 250588 480836
rect 251180 480888 251232 480894
rect 251180 480830 251232 480836
rect 249996 470566 250116 470594
rect 249996 468654 250024 470566
rect 249984 468648 250036 468654
rect 249984 468590 250036 468596
rect 251192 467294 251220 480830
rect 251468 478122 251496 488022
rect 251548 481160 251600 481166
rect 251548 481102 251600 481108
rect 251284 478094 251496 478122
rect 251284 467362 251312 478094
rect 251560 473354 251588 481102
rect 251928 480894 251956 488022
rect 251916 480888 251968 480894
rect 251916 480830 251968 480836
rect 252560 480888 252612 480894
rect 252560 480830 252612 480836
rect 251376 473326 251588 473354
rect 251376 468586 251404 473326
rect 251364 468580 251416 468586
rect 251364 468522 251416 468528
rect 252572 468518 252600 480830
rect 252664 472977 252692 488022
rect 252756 488022 253046 488050
rect 253216 488022 253506 488050
rect 252756 478378 252784 488022
rect 253216 480894 253244 488022
rect 253204 480888 253256 480894
rect 253204 480830 253256 480836
rect 252744 478372 252796 478378
rect 252744 478314 252796 478320
rect 252650 472968 252706 472977
rect 252650 472903 252706 472912
rect 252560 468512 252612 468518
rect 252560 468454 252612 468460
rect 251272 467356 251324 467362
rect 251272 467298 251324 467304
rect 251180 467288 251232 467294
rect 251180 467230 251232 467236
rect 253952 467226 253980 488036
rect 254044 488022 254426 488050
rect 254504 488022 254794 488050
rect 254872 488022 255254 488050
rect 255332 488022 255714 488050
rect 256190 488022 256280 488050
rect 254044 475590 254072 488022
rect 254504 479738 254532 488022
rect 254492 479732 254544 479738
rect 254492 479674 254544 479680
rect 254872 478514 254900 488022
rect 254860 478508 254912 478514
rect 254860 478450 254912 478456
rect 254032 475584 254084 475590
rect 254032 475526 254084 475532
rect 255332 468790 255360 488022
rect 256252 482497 256280 488022
rect 256344 488022 256634 488050
rect 256712 488022 257002 488050
rect 257478 488022 257568 488050
rect 256238 482488 256294 482497
rect 256238 482423 256294 482432
rect 256344 479942 256372 488022
rect 256332 479936 256384 479942
rect 256332 479878 256384 479884
rect 255320 468784 255372 468790
rect 255320 468726 255372 468732
rect 256712 467498 256740 488022
rect 257540 482526 257568 488022
rect 257632 488022 257922 488050
rect 258184 488022 258382 488050
rect 258552 488022 258842 488050
rect 258920 488022 259210 488050
rect 259564 488022 259670 488050
rect 257528 482520 257580 482526
rect 257528 482462 257580 482468
rect 257632 474434 257660 488022
rect 258080 480888 258132 480894
rect 258080 480830 258132 480836
rect 257620 474428 257672 474434
rect 257620 474370 257672 474376
rect 256700 467492 256752 467498
rect 256700 467434 256752 467440
rect 253940 467220 253992 467226
rect 253940 467162 253992 467168
rect 258092 466274 258120 480830
rect 258184 467430 258212 488022
rect 258552 480894 258580 488022
rect 258540 480888 258592 480894
rect 258540 480830 258592 480836
rect 258920 475658 258948 488022
rect 259564 479806 259592 488022
rect 260116 483818 260144 488036
rect 260208 488022 260590 488050
rect 260974 488022 261248 488050
rect 260104 483812 260156 483818
rect 260104 483754 260156 483760
rect 259552 479800 259604 479806
rect 259552 479742 259604 479748
rect 260208 476114 260236 488022
rect 261220 481234 261248 488022
rect 261404 482594 261432 488036
rect 261496 488022 261878 488050
rect 262354 488022 262444 488050
rect 261392 482588 261444 482594
rect 261392 482530 261444 482536
rect 261208 481228 261260 481234
rect 261208 481170 261260 481176
rect 259472 476086 260236 476114
rect 258908 475652 258960 475658
rect 258908 475594 258960 475600
rect 259472 474298 259500 476086
rect 259460 474292 259512 474298
rect 259460 474234 259512 474240
rect 261496 470594 261524 488022
rect 262416 485790 262444 488022
rect 262508 488022 262798 488050
rect 262876 488022 263166 488050
rect 262404 485784 262456 485790
rect 262404 485726 262456 485732
rect 262508 481114 262536 488022
rect 262588 485784 262640 485790
rect 262588 485726 262640 485732
rect 260852 470566 261524 470594
rect 262232 481086 262536 481114
rect 258172 467424 258224 467430
rect 258172 467366 258224 467372
rect 258080 466268 258132 466274
rect 258080 466210 258132 466216
rect 260852 466206 260880 470566
rect 262232 467158 262260 481086
rect 262312 480888 262364 480894
rect 262312 480830 262364 480836
rect 262324 472870 262352 480830
rect 262600 474366 262628 485726
rect 262876 480894 262904 488022
rect 262864 480888 262916 480894
rect 262864 480830 262916 480836
rect 262588 474360 262640 474366
rect 262588 474302 262640 474308
rect 262312 472864 262364 472870
rect 262312 472806 262364 472812
rect 263612 472802 263640 488036
rect 263796 488022 264086 488050
rect 264256 488022 264546 488050
rect 265022 488022 265112 488050
rect 263692 484152 263744 484158
rect 263692 484094 263744 484100
rect 263704 477086 263732 484094
rect 263692 477080 263744 477086
rect 263692 477022 263744 477028
rect 263796 477018 263824 488022
rect 264256 484158 264284 488022
rect 264244 484152 264296 484158
rect 264244 484094 264296 484100
rect 264980 484152 265032 484158
rect 264980 484094 265032 484100
rect 263784 477012 263836 477018
rect 263784 476954 263836 476960
rect 263600 472796 263652 472802
rect 263600 472738 263652 472744
rect 264992 468858 265020 484094
rect 265084 477154 265112 488022
rect 265176 488022 265374 488050
rect 265544 488022 265834 488050
rect 265912 488022 266294 488050
rect 266372 488022 266754 488050
rect 266832 488022 267122 488050
rect 267200 488022 267582 488050
rect 267752 488022 268042 488050
rect 268120 488022 268502 488050
rect 268978 488022 269068 488050
rect 265176 477358 265204 488022
rect 265544 484158 265572 488022
rect 265532 484152 265584 484158
rect 265532 484094 265584 484100
rect 265912 479874 265940 488022
rect 265900 479868 265952 479874
rect 265900 479810 265952 479816
rect 265164 477352 265216 477358
rect 265164 477294 265216 477300
rect 265072 477148 265124 477154
rect 265072 477090 265124 477096
rect 266372 468994 266400 488022
rect 266832 484106 266860 488022
rect 266464 484078 266860 484106
rect 266464 469062 266492 484078
rect 267200 470594 267228 488022
rect 266556 470566 267228 470594
rect 266556 469130 266584 470566
rect 266544 469124 266596 469130
rect 266544 469066 266596 469072
rect 266452 469056 266504 469062
rect 266452 468998 266504 469004
rect 266360 468988 266412 468994
rect 266360 468930 266412 468936
rect 264980 468852 265032 468858
rect 264980 468794 265032 468800
rect 267752 468722 267780 488022
rect 268120 477290 268148 488022
rect 269040 481302 269068 488022
rect 269120 484152 269172 484158
rect 269120 484094 269172 484100
rect 269028 481296 269080 481302
rect 269028 481238 269080 481244
rect 268108 477284 268160 477290
rect 268108 477226 268160 477232
rect 269132 475726 269160 484094
rect 269316 481166 269344 488036
rect 269408 488022 269790 488050
rect 269960 488022 270250 488050
rect 270604 488022 270710 488050
rect 270880 488022 271170 488050
rect 271554 488022 271828 488050
rect 269304 481160 269356 481166
rect 269304 481102 269356 481108
rect 269408 478446 269436 488022
rect 269960 484158 269988 488022
rect 269948 484152 270000 484158
rect 269948 484094 270000 484100
rect 270500 484152 270552 484158
rect 270500 484094 270552 484100
rect 269396 478440 269448 478446
rect 269396 478382 269448 478388
rect 269120 475720 269172 475726
rect 270512 475697 270540 484094
rect 270604 478582 270632 488022
rect 270880 484158 270908 488022
rect 270868 484152 270920 484158
rect 270868 484094 270920 484100
rect 271800 482798 271828 488022
rect 271892 488022 271998 488050
rect 272076 488022 272458 488050
rect 272536 488022 272918 488050
rect 271788 482792 271840 482798
rect 271788 482734 271840 482740
rect 270592 478576 270644 478582
rect 270592 478518 270644 478524
rect 269120 475662 269172 475668
rect 270498 475688 270554 475697
rect 270498 475623 270554 475632
rect 267740 468716 267792 468722
rect 267740 468658 267792 468664
rect 262220 467152 262272 467158
rect 262220 467094 262272 467100
rect 260840 466200 260892 466206
rect 260840 466142 260892 466148
rect 249892 465996 249944 466002
rect 249892 465938 249944 465944
rect 248604 465860 248656 465866
rect 248604 465802 248656 465808
rect 248418 465760 248474 465769
rect 220912 465724 220964 465730
rect 220912 465666 220964 465672
rect 242900 465724 242952 465730
rect 248418 465695 248474 465704
rect 242900 465666 242952 465672
rect 271892 464370 271920 488022
rect 271972 484152 272024 484158
rect 271972 484094 272024 484100
rect 271984 466342 272012 484094
rect 272076 468926 272104 488022
rect 272536 484158 272564 488022
rect 272524 484152 272576 484158
rect 272524 484094 272576 484100
rect 273272 469198 273300 488036
rect 273456 488022 273746 488050
rect 273824 488022 274206 488050
rect 273352 484152 273404 484158
rect 273352 484094 273404 484100
rect 273364 472938 273392 484094
rect 273456 474638 273484 488022
rect 273824 484158 273852 488022
rect 274668 487830 274696 488036
rect 274744 488022 275126 488050
rect 275510 488022 275600 488050
rect 274656 487824 274708 487830
rect 274656 487766 274708 487772
rect 273812 484152 273864 484158
rect 274744 484106 274772 488022
rect 274824 487824 274876 487830
rect 274824 487766 274876 487772
rect 273812 484094 273864 484100
rect 274652 484078 274772 484106
rect 273444 474632 273496 474638
rect 273444 474574 273496 474580
rect 273352 472932 273404 472938
rect 273352 472874 273404 472880
rect 273260 469192 273312 469198
rect 273260 469134 273312 469140
rect 272064 468920 272116 468926
rect 272064 468862 272116 468868
rect 274652 467566 274680 484078
rect 274836 482866 274864 487766
rect 275572 483886 275600 488022
rect 275664 488022 275954 488050
rect 276430 488022 276704 488050
rect 275560 483880 275612 483886
rect 275560 483822 275612 483828
rect 274824 482860 274876 482866
rect 274824 482802 274876 482808
rect 275664 477222 275692 488022
rect 276676 482730 276704 488022
rect 276664 482724 276716 482730
rect 276664 482666 276716 482672
rect 276860 482662 276888 488036
rect 276952 488022 277334 488050
rect 277412 488022 277702 488050
rect 277780 488022 278162 488050
rect 278240 488022 278622 488050
rect 278792 488022 279082 488050
rect 279558 488022 279832 488050
rect 279926 488022 280108 488050
rect 276848 482656 276900 482662
rect 276848 482598 276900 482604
rect 275652 477216 275704 477222
rect 275652 477158 275704 477164
rect 276952 471510 276980 488022
rect 276940 471504 276992 471510
rect 276940 471446 276992 471452
rect 274640 467560 274692 467566
rect 274640 467502 274692 467508
rect 271972 466336 272024 466342
rect 271972 466278 272024 466284
rect 277412 465905 277440 488022
rect 277780 484140 277808 488022
rect 277504 484112 277808 484140
rect 277504 467634 277532 484112
rect 278240 474502 278268 488022
rect 278792 480010 278820 488022
rect 279804 483954 279832 488022
rect 280080 484022 280108 488022
rect 280172 488022 280370 488050
rect 280448 488022 280830 488050
rect 281306 488022 281488 488050
rect 280068 484016 280120 484022
rect 280068 483958 280120 483964
rect 279792 483948 279844 483954
rect 279792 483890 279844 483896
rect 278780 480004 278832 480010
rect 278780 479946 278832 479952
rect 278228 474496 278280 474502
rect 278228 474438 278280 474444
rect 280172 468450 280200 488022
rect 280448 474570 280476 488022
rect 281460 481370 281488 488022
rect 281644 484294 281672 488036
rect 281736 488022 282118 488050
rect 282196 488022 282578 488050
rect 281632 484288 281684 484294
rect 281632 484230 281684 484236
rect 281736 484140 281764 488022
rect 281552 484112 281764 484140
rect 281448 481364 281500 481370
rect 281448 481306 281500 481312
rect 280436 474564 280488 474570
rect 280436 474506 280488 474512
rect 281552 469946 281580 484112
rect 282196 470594 282224 488022
rect 282920 480888 282972 480894
rect 282920 480830 282972 480836
rect 281644 470566 282224 470594
rect 281540 469940 281592 469946
rect 281540 469882 281592 469888
rect 281644 469878 281672 470566
rect 282932 470490 282960 480830
rect 282920 470484 282972 470490
rect 282920 470426 282972 470432
rect 283024 470354 283052 488036
rect 283116 488022 283498 488050
rect 283576 488022 283866 488050
rect 284342 488022 284432 488050
rect 283116 470422 283144 488022
rect 283576 480894 283604 488022
rect 283564 480888 283616 480894
rect 283564 480830 283616 480836
rect 284300 480888 284352 480894
rect 284300 480830 284352 480836
rect 283104 470416 283156 470422
rect 283104 470358 283156 470364
rect 283012 470348 283064 470354
rect 283012 470290 283064 470296
rect 284312 470082 284340 480830
rect 284300 470076 284352 470082
rect 284300 470018 284352 470024
rect 284404 470014 284432 488022
rect 284496 488022 284786 488050
rect 285262 488022 285536 488050
rect 285722 488022 285812 488050
rect 284496 480894 284524 488022
rect 285508 481438 285536 488022
rect 285784 485790 285812 488022
rect 285876 488022 286074 488050
rect 286152 488022 286534 488050
rect 286704 488022 286994 488050
rect 287348 488022 287454 488050
rect 287532 488022 287822 488050
rect 287992 488022 288282 488050
rect 288452 488022 288742 488050
rect 288820 488022 289202 488050
rect 289280 488022 289662 488050
rect 290046 488022 290136 488050
rect 285772 485784 285824 485790
rect 285772 485726 285824 485732
rect 285496 481432 285548 481438
rect 285496 481374 285548 481380
rect 285876 481114 285904 488022
rect 285956 485784 286008 485790
rect 285956 485726 286008 485732
rect 285692 481086 285904 481114
rect 284484 480888 284536 480894
rect 284484 480830 284536 480836
rect 285692 470286 285720 481086
rect 285968 480842 285996 485726
rect 285784 480814 285996 480842
rect 285680 470280 285732 470286
rect 285680 470222 285732 470228
rect 285784 470150 285812 480814
rect 286152 479777 286180 488022
rect 286138 479768 286194 479777
rect 286138 479703 286194 479712
rect 286704 476114 286732 488022
rect 287060 480888 287112 480894
rect 287060 480830 287112 480836
rect 285876 476086 286732 476114
rect 285876 471442 285904 476086
rect 285864 471436 285916 471442
rect 285864 471378 285916 471384
rect 287072 470218 287100 480830
rect 287348 477426 287376 488022
rect 287336 477420 287388 477426
rect 287336 477362 287388 477368
rect 287532 476114 287560 488022
rect 287992 480894 288020 488022
rect 287980 480888 288032 480894
rect 287980 480830 288032 480836
rect 287164 476086 287560 476114
rect 287164 471918 287192 476086
rect 287152 471912 287204 471918
rect 287152 471854 287204 471860
rect 287060 470212 287112 470218
rect 287060 470154 287112 470160
rect 285772 470144 285824 470150
rect 285772 470086 285824 470092
rect 284392 470008 284444 470014
rect 284392 469950 284444 469956
rect 281632 469872 281684 469878
rect 281632 469814 281684 469820
rect 280160 468444 280212 468450
rect 280160 468386 280212 468392
rect 288452 467702 288480 488022
rect 288820 476114 288848 488022
rect 289280 477494 289308 488022
rect 290108 482934 290136 488022
rect 290200 488022 290490 488050
rect 290568 488022 290950 488050
rect 291304 488022 291410 488050
rect 291488 488022 291870 488050
rect 291948 488022 292238 488050
rect 292592 488022 292698 488050
rect 292776 488022 293158 488050
rect 293328 488022 293618 488050
rect 290096 482928 290148 482934
rect 290096 482870 290148 482876
rect 289820 480888 289872 480894
rect 289820 480830 289872 480836
rect 289268 477488 289320 477494
rect 289268 477430 289320 477436
rect 288544 476086 288848 476114
rect 288544 471578 288572 476086
rect 289832 473074 289860 480830
rect 290200 473958 290228 488022
rect 290568 480894 290596 488022
rect 291304 481506 291332 488022
rect 291488 485774 291516 488022
rect 291396 485746 291516 485774
rect 291292 481500 291344 481506
rect 291292 481442 291344 481448
rect 290556 480888 290608 480894
rect 290556 480830 290608 480836
rect 291396 478122 291424 485746
rect 291476 481500 291528 481506
rect 291476 481442 291528 481448
rect 291212 478094 291424 478122
rect 290188 473952 290240 473958
rect 290188 473894 290240 473900
rect 289820 473068 289872 473074
rect 289820 473010 289872 473016
rect 288532 471572 288584 471578
rect 288532 471514 288584 471520
rect 288440 467696 288492 467702
rect 288440 467638 288492 467644
rect 277492 467628 277544 467634
rect 277492 467570 277544 467576
rect 277398 465896 277454 465905
rect 277398 465831 277454 465840
rect 291212 464438 291240 478094
rect 291488 473354 291516 481442
rect 291948 474706 291976 488022
rect 292592 475794 292620 488022
rect 292776 476746 292804 488022
rect 293328 480146 293356 488022
rect 293972 484158 294000 488036
rect 294064 488022 294446 488050
rect 294616 488022 294906 488050
rect 295382 488022 295564 488050
rect 293960 484152 294012 484158
rect 293960 484094 294012 484100
rect 293960 480888 294012 480894
rect 293960 480830 294012 480836
rect 293316 480140 293368 480146
rect 293316 480082 293368 480088
rect 292764 476740 292816 476746
rect 292764 476682 292816 476688
rect 292580 475788 292632 475794
rect 292580 475730 292632 475736
rect 291936 474700 291988 474706
rect 291936 474642 291988 474648
rect 291304 473326 291516 473354
rect 291304 467770 291332 473326
rect 293972 467838 294000 480830
rect 294064 473006 294092 488022
rect 294616 480894 294644 488022
rect 295536 481506 295564 488022
rect 295628 488022 295826 488050
rect 295904 488022 296194 488050
rect 296272 488022 296654 488050
rect 296824 488022 297114 488050
rect 297192 488022 297574 488050
rect 297744 488022 298034 488050
rect 298204 488022 298402 488050
rect 298480 488022 298862 488050
rect 299032 488022 299322 488050
rect 299492 488022 299782 488050
rect 295524 481500 295576 481506
rect 295524 481442 295576 481448
rect 294604 480888 294656 480894
rect 294604 480830 294656 480836
rect 295340 480888 295392 480894
rect 295340 480830 295392 480836
rect 294052 473000 294104 473006
rect 294052 472942 294104 472948
rect 293960 467832 294012 467838
rect 293960 467774 294012 467780
rect 291292 467764 291344 467770
rect 291292 467706 291344 467712
rect 295352 464506 295380 480830
rect 295628 478122 295656 488022
rect 295708 481500 295760 481506
rect 295708 481442 295760 481448
rect 295444 478094 295656 478122
rect 295444 466410 295472 478094
rect 295720 473354 295748 481442
rect 295904 480894 295932 488022
rect 295892 480888 295944 480894
rect 295892 480830 295944 480836
rect 295536 473326 295748 473354
rect 295536 471209 295564 473326
rect 296272 471986 296300 488022
rect 296720 480888 296772 480894
rect 296720 480830 296772 480836
rect 296260 471980 296312 471986
rect 296260 471922 296312 471928
rect 295522 471200 295578 471209
rect 295522 471135 295578 471144
rect 296732 468489 296760 480830
rect 296824 471345 296852 488022
rect 297192 480894 297220 488022
rect 297180 480888 297232 480894
rect 297180 480830 297232 480836
rect 297744 471646 297772 488022
rect 298204 485774 298232 488022
rect 298480 485774 298508 488022
rect 298112 485746 298232 485774
rect 298388 485746 298508 485774
rect 298112 483014 298140 485746
rect 298388 483014 298416 485746
rect 298020 482986 298140 483014
rect 298204 482986 298416 483014
rect 298020 478106 298048 482986
rect 298204 478122 298232 482986
rect 298008 478100 298060 478106
rect 298008 478042 298060 478048
rect 298112 478094 298232 478122
rect 298284 478100 298336 478106
rect 298112 471782 298140 478094
rect 298284 478042 298336 478048
rect 298192 477624 298244 477630
rect 298192 477566 298244 477572
rect 298204 471850 298232 477566
rect 298192 471844 298244 471850
rect 298192 471786 298244 471792
rect 298100 471776 298152 471782
rect 298100 471718 298152 471724
rect 298296 471714 298324 478042
rect 299032 477630 299060 488022
rect 299492 480078 299520 488022
rect 318076 482225 318104 623766
rect 318168 567934 318196 642330
rect 322296 642252 322348 642258
rect 322296 642194 322348 642200
rect 320916 642048 320968 642054
rect 320916 641990 320968 641996
rect 319444 641232 319496 641238
rect 319444 641174 319496 641180
rect 319456 575006 319484 641174
rect 319536 640552 319588 640558
rect 319536 640494 319588 640500
rect 319444 575000 319496 575006
rect 319444 574942 319496 574948
rect 319548 574666 319576 640494
rect 319628 640416 319680 640422
rect 319628 640358 319680 640364
rect 319640 575278 319668 640358
rect 320822 639296 320878 639305
rect 320822 639231 320878 639240
rect 319628 575272 319680 575278
rect 319628 575214 319680 575220
rect 319536 574660 319588 574666
rect 319536 574602 319588 574608
rect 318156 567928 318208 567934
rect 318156 567870 318208 567876
rect 320836 554266 320864 639231
rect 320928 558278 320956 641990
rect 322204 640484 322256 640490
rect 322204 640426 322256 640432
rect 321008 638240 321060 638246
rect 321008 638182 321060 638188
rect 321020 576745 321048 638182
rect 321558 634536 321614 634545
rect 321558 634471 321614 634480
rect 321572 633486 321600 634471
rect 321560 633480 321612 633486
rect 321560 633422 321612 633428
rect 321558 629776 321614 629785
rect 321558 629711 321614 629720
rect 321572 629338 321600 629711
rect 321560 629332 321612 629338
rect 321560 629274 321612 629280
rect 321558 625016 321614 625025
rect 321558 624951 321614 624960
rect 321572 623830 321600 624951
rect 321560 623824 321612 623830
rect 321560 623766 321612 623772
rect 321558 620256 321614 620265
rect 321558 620191 321614 620200
rect 321572 619682 321600 620191
rect 321560 619676 321612 619682
rect 321560 619618 321612 619624
rect 321558 615496 321614 615505
rect 321558 615431 321614 615440
rect 321572 614174 321600 615431
rect 321560 614168 321612 614174
rect 321560 614110 321612 614116
rect 321558 610736 321614 610745
rect 321558 610671 321614 610680
rect 321572 610026 321600 610671
rect 321560 610020 321612 610026
rect 321560 609962 321612 609968
rect 321558 605976 321614 605985
rect 321558 605911 321614 605920
rect 321572 605878 321600 605911
rect 321560 605872 321612 605878
rect 321560 605814 321612 605820
rect 321558 596456 321614 596465
rect 321558 596391 321614 596400
rect 321572 596222 321600 596391
rect 321560 596216 321612 596222
rect 321560 596158 321612 596164
rect 321558 591696 321614 591705
rect 321558 591631 321614 591640
rect 321572 590714 321600 591631
rect 321560 590708 321612 590714
rect 321560 590650 321612 590656
rect 321558 586936 321614 586945
rect 321558 586871 321614 586880
rect 321572 586566 321600 586871
rect 321560 586560 321612 586566
rect 321560 586502 321612 586508
rect 321558 581496 321614 581505
rect 321558 581431 321614 581440
rect 321572 581058 321600 581431
rect 321560 581052 321612 581058
rect 321560 580994 321612 581000
rect 321006 576736 321062 576745
rect 321006 576671 321062 576680
rect 321558 571976 321614 571985
rect 321558 571911 321614 571920
rect 321572 570654 321600 571911
rect 321560 570648 321612 570654
rect 321560 570590 321612 570596
rect 321560 567248 321612 567254
rect 321558 567216 321560 567225
rect 321612 567216 321614 567225
rect 321558 567151 321614 567160
rect 321558 562456 321614 562465
rect 321558 562391 321614 562400
rect 321572 561746 321600 562391
rect 321560 561740 321612 561746
rect 321560 561682 321612 561688
rect 321560 558884 321612 558890
rect 321560 558826 321612 558832
rect 320916 558272 320968 558278
rect 320916 558214 320968 558220
rect 321572 557705 321600 558826
rect 321558 557696 321614 557705
rect 321558 557631 321614 557640
rect 320824 554260 320876 554266
rect 320824 554202 320876 554208
rect 321558 552936 321614 552945
rect 321558 552871 321614 552880
rect 319536 552560 319588 552566
rect 319536 552502 319588 552508
rect 319444 550656 319496 550662
rect 319444 550598 319496 550604
rect 319456 524414 319484 550598
rect 319548 528562 319576 552502
rect 321008 552492 321060 552498
rect 321008 552434 321060 552440
rect 320916 552152 320968 552158
rect 320916 552094 320968 552100
rect 320824 552084 320876 552090
rect 320824 552026 320876 552032
rect 319536 528556 319588 528562
rect 319536 528498 319588 528504
rect 319444 524408 319496 524414
rect 319444 524350 319496 524356
rect 320836 524278 320864 552026
rect 320824 524272 320876 524278
rect 320824 524214 320876 524220
rect 320928 524210 320956 552094
rect 321020 524346 321048 552434
rect 321100 552288 321152 552294
rect 321100 552230 321152 552236
rect 321112 525570 321140 552230
rect 321572 552226 321600 552871
rect 321560 552220 321612 552226
rect 321560 552162 321612 552168
rect 321192 551472 321244 551478
rect 321192 551414 321244 551420
rect 321204 526969 321232 551414
rect 321284 550044 321336 550050
rect 321284 549986 321336 549992
rect 321296 528086 321324 549986
rect 322216 549953 322244 640426
rect 322308 556986 322336 642194
rect 322388 641844 322440 641850
rect 322388 641786 322440 641792
rect 322400 563854 322428 641786
rect 322492 572014 322520 642670
rect 322584 573578 322612 643078
rect 346584 642728 346636 642734
rect 346584 642670 346636 642676
rect 323676 642660 323728 642666
rect 323676 642602 323728 642608
rect 323584 640960 323636 640966
rect 323584 640902 323636 640908
rect 322664 640892 322716 640898
rect 322664 640834 322716 640840
rect 322676 603770 322704 640834
rect 322664 603764 322716 603770
rect 322664 603706 322716 603712
rect 322572 573572 322624 573578
rect 322572 573514 322624 573520
rect 322480 572008 322532 572014
rect 322480 571950 322532 571956
rect 322388 563848 322440 563854
rect 322388 563790 322440 563796
rect 322296 556980 322348 556986
rect 322296 556922 322348 556928
rect 322480 552628 322532 552634
rect 322480 552570 322532 552576
rect 322296 552356 322348 552362
rect 322296 552298 322348 552304
rect 322202 549944 322258 549953
rect 322202 549879 322258 549888
rect 321560 548616 321612 548622
rect 321560 548558 321612 548564
rect 321572 548185 321600 548558
rect 322112 548548 322164 548554
rect 322112 548490 322164 548496
rect 321558 548176 321614 548185
rect 321558 548111 321614 548120
rect 321560 543720 321612 543726
rect 321560 543662 321612 543668
rect 321572 543425 321600 543662
rect 321558 543416 321614 543425
rect 321558 543351 321614 543360
rect 321560 539572 321612 539578
rect 321560 539514 321612 539520
rect 321572 538665 321600 539514
rect 321558 538656 321614 538665
rect 321558 538591 321614 538600
rect 322124 533905 322152 548490
rect 322202 548040 322258 548049
rect 322202 547975 322258 547984
rect 322110 533896 322166 533905
rect 322110 533831 322166 533840
rect 321284 528080 321336 528086
rect 321284 528022 321336 528028
rect 321190 526960 321246 526969
rect 321190 526895 321246 526904
rect 322216 526833 322244 547975
rect 322202 526824 322258 526833
rect 322202 526759 322258 526768
rect 322308 525638 322336 552298
rect 322388 550792 322440 550798
rect 322388 550734 322440 550740
rect 322400 525706 322428 550734
rect 322492 528426 322520 552570
rect 322664 552424 322716 552430
rect 322664 552366 322716 552372
rect 322572 551064 322624 551070
rect 322572 551006 322624 551012
rect 322480 528420 322532 528426
rect 322480 528362 322532 528368
rect 322584 526794 322612 551006
rect 322676 528494 322704 552366
rect 322756 550112 322808 550118
rect 322756 550054 322808 550060
rect 322768 529514 322796 550054
rect 323596 549914 323624 640902
rect 323688 554198 323716 642602
rect 342260 642592 342312 642598
rect 342260 642534 342312 642540
rect 323768 642456 323820 642462
rect 323768 642398 323820 642404
rect 323780 555626 323808 642398
rect 324872 642320 324924 642326
rect 324872 642262 324924 642268
rect 323952 642116 324004 642122
rect 323952 642058 324004 642064
rect 323860 641776 323912 641782
rect 323860 641718 323912 641724
rect 323872 561066 323900 641718
rect 323964 561134 323992 642058
rect 324778 641744 324834 641753
rect 324778 641679 324834 641688
rect 324228 641096 324280 641102
rect 324228 641038 324280 641044
rect 324240 601225 324268 641038
rect 324226 601216 324282 601225
rect 324226 601151 324282 601160
rect 324044 573368 324096 573374
rect 324044 573310 324096 573316
rect 323952 561128 324004 561134
rect 323952 561070 324004 561076
rect 323860 561060 323912 561066
rect 323860 561002 323912 561008
rect 323768 555620 323820 555626
rect 323768 555562 323820 555568
rect 323676 554192 323728 554198
rect 323676 554134 323728 554140
rect 323676 550996 323728 551002
rect 323676 550938 323728 550944
rect 323584 549908 323636 549914
rect 323584 549850 323636 549856
rect 322848 548820 322900 548826
rect 322848 548762 322900 548768
rect 322756 529508 322808 529514
rect 322756 529450 322808 529456
rect 322664 528488 322716 528494
rect 322664 528430 322716 528436
rect 322860 528358 322888 548762
rect 323584 548072 323636 548078
rect 323584 548014 323636 548020
rect 322848 528352 322900 528358
rect 322848 528294 322900 528300
rect 323596 526998 323624 548014
rect 323584 526992 323636 526998
rect 323584 526934 323636 526940
rect 322572 526788 322624 526794
rect 322572 526730 322624 526736
rect 323688 526386 323716 550938
rect 323950 549808 324006 549817
rect 323950 549743 324006 549752
rect 323768 549364 323820 549370
rect 323768 549306 323820 549312
rect 323780 528290 323808 549306
rect 323860 548208 323912 548214
rect 323860 548150 323912 548156
rect 323768 528284 323820 528290
rect 323768 528226 323820 528232
rect 323872 527066 323900 548150
rect 323964 528193 323992 549743
rect 323950 528184 324006 528193
rect 323950 528119 324006 528128
rect 323860 527060 323912 527066
rect 323860 527002 323912 527008
rect 324056 526697 324084 573310
rect 324792 569362 324820 641679
rect 324780 569356 324832 569362
rect 324780 569298 324832 569304
rect 324884 566642 324912 642262
rect 337568 642184 337620 642190
rect 337568 642126 337620 642132
rect 337108 641912 337160 641918
rect 337108 641854 337160 641860
rect 328552 641776 328604 641782
rect 328552 641718 328604 641724
rect 328564 639962 328592 641718
rect 328564 639934 328900 639962
rect 337120 639742 337148 641854
rect 337580 639962 337608 642126
rect 342272 639962 342300 642534
rect 346596 639962 346624 642670
rect 401692 642660 401744 642666
rect 401692 642602 401744 642608
rect 374000 642524 374052 642530
rect 374000 642466 374052 642472
rect 369124 642456 369176 642462
rect 369124 642398 369176 642404
rect 364616 642388 364668 642394
rect 355520 642348 355732 642376
rect 347596 642184 347648 642190
rect 347596 642126 347648 642132
rect 337580 639934 337916 639962
rect 342272 639934 342424 639962
rect 346596 639934 346932 639962
rect 337108 639736 337160 639742
rect 337108 639678 337160 639684
rect 347608 639674 347636 642126
rect 351092 641912 351144 641918
rect 351092 641854 351144 641860
rect 351104 639962 351132 641854
rect 351104 639934 351440 639962
rect 347596 639668 347648 639674
rect 347596 639610 347648 639616
rect 355520 639606 355548 642348
rect 355704 642258 355732 642348
rect 364616 642330 364668 642336
rect 355600 642252 355652 642258
rect 355600 642194 355652 642200
rect 355692 642252 355744 642258
rect 355692 642194 355744 642200
rect 355612 639962 355640 642194
rect 360200 641164 360252 641170
rect 360200 641106 360252 641112
rect 360212 639962 360240 641106
rect 364628 639962 364656 642330
rect 365628 641776 365680 641782
rect 365628 641718 365680 641724
rect 365640 641034 365668 641718
rect 365628 641028 365680 641034
rect 365628 640970 365680 640976
rect 369136 639962 369164 642398
rect 374012 639962 374040 642466
rect 378140 642320 378192 642326
rect 378140 642262 378192 642268
rect 355612 639934 355948 639962
rect 360212 639934 360456 639962
rect 364628 639934 364964 639962
rect 369136 639934 369472 639962
rect 373980 639934 374040 639962
rect 378152 639962 378180 642262
rect 387800 642116 387852 642122
rect 387800 642058 387852 642064
rect 383660 641980 383712 641986
rect 383660 641922 383712 641928
rect 383672 639962 383700 641922
rect 378152 639934 378488 639962
rect 383640 639934 383700 639962
rect 387812 639962 387840 642058
rect 392308 642048 392360 642054
rect 392308 641990 392360 641996
rect 392320 639962 392348 641990
rect 396816 640688 396868 640694
rect 396816 640630 396868 640636
rect 396828 639962 396856 640630
rect 387812 639934 388148 639962
rect 392320 639934 392656 639962
rect 396828 639934 397164 639962
rect 401704 639826 401732 642602
rect 405936 639962 405964 646478
rect 428372 645176 428424 645182
rect 428372 645118 428424 645124
rect 414848 642252 414900 642258
rect 414848 642194 414900 642200
rect 410340 642184 410392 642190
rect 410340 642126 410392 642132
rect 410352 639962 410380 642126
rect 414860 639962 414888 642194
rect 419540 641776 419592 641782
rect 419540 641718 419592 641724
rect 423862 641744 423918 641753
rect 419552 639962 419580 641718
rect 423862 641679 423918 641688
rect 423876 639962 423904 641679
rect 428384 639962 428412 645118
rect 432880 641844 432932 641850
rect 432880 641786 432932 641792
rect 432892 639962 432920 641786
rect 405936 639934 406180 639962
rect 410352 639934 410688 639962
rect 414860 639934 415196 639962
rect 419552 639934 419704 639962
rect 423876 639934 424212 639962
rect 428384 639934 428720 639962
rect 432892 639934 433228 639962
rect 401672 639798 401732 639826
rect 355508 639600 355560 639606
rect 333058 639568 333114 639577
rect 333114 639526 333408 639554
rect 355508 639542 355560 639548
rect 333058 639503 333114 639512
rect 433340 639124 433392 639130
rect 433340 639066 433392 639072
rect 433352 626249 433380 639066
rect 433338 626240 433394 626249
rect 433338 626175 433394 626184
rect 433338 615904 433394 615913
rect 433338 615839 433394 615848
rect 324872 566636 324924 566642
rect 324872 566578 324924 566584
rect 324780 550928 324832 550934
rect 324780 550870 324832 550876
rect 324688 550860 324740 550866
rect 324688 550802 324740 550808
rect 324136 549500 324188 549506
rect 324136 549442 324188 549448
rect 324148 528018 324176 549442
rect 324596 548480 324648 548486
rect 324596 548422 324648 548428
rect 324504 548276 324556 548282
rect 324504 548218 324556 548224
rect 324136 528012 324188 528018
rect 324136 527954 324188 527960
rect 324516 526862 324544 548218
rect 324608 527134 324636 548422
rect 324700 533458 324728 550802
rect 324688 533452 324740 533458
rect 324688 533394 324740 533400
rect 324792 533338 324820 550870
rect 324872 550724 324924 550730
rect 324872 550666 324924 550672
rect 324700 533310 324820 533338
rect 324596 527128 324648 527134
rect 324596 527070 324648 527076
rect 324504 526856 324556 526862
rect 324504 526798 324556 526804
rect 324042 526688 324098 526697
rect 324042 526623 324098 526632
rect 324700 526454 324728 533310
rect 324780 533248 324832 533254
rect 324780 533190 324832 533196
rect 324792 526658 324820 533190
rect 324884 526930 324912 550666
rect 325036 529094 325096 529122
rect 329544 529094 329788 529122
rect 334052 529094 334112 529122
rect 325068 528554 325096 529094
rect 324976 528526 325096 528554
rect 324976 527202 325004 528526
rect 324964 527196 325016 527202
rect 324964 527138 325016 527144
rect 324872 526924 324924 526930
rect 324872 526866 324924 526872
rect 324780 526652 324832 526658
rect 324780 526594 324832 526600
rect 324688 526448 324740 526454
rect 324688 526390 324740 526396
rect 323676 526380 323728 526386
rect 323676 526322 323728 526328
rect 322388 525700 322440 525706
rect 322388 525642 322440 525648
rect 322296 525632 322348 525638
rect 322296 525574 322348 525580
rect 321100 525564 321152 525570
rect 321100 525506 321152 525512
rect 321008 524340 321060 524346
rect 321008 524282 321060 524288
rect 320916 524204 320968 524210
rect 320916 524146 320968 524152
rect 329760 524142 329788 529094
rect 334084 528554 334112 529094
rect 333992 528526 334112 528554
rect 338224 529094 338560 529122
rect 342732 529094 343068 529122
rect 347240 529094 347576 529122
rect 351932 529094 352084 529122
rect 356256 529094 356592 529122
rect 360764 529094 361100 529122
rect 365272 529094 365608 529122
rect 369872 529094 370116 529122
rect 374288 529094 374624 529122
rect 379532 529094 379776 529122
rect 383672 529094 384284 529122
rect 388456 529094 388792 529122
rect 393300 529094 393360 529122
rect 333992 526250 334020 528526
rect 338224 526998 338252 529094
rect 338212 526992 338264 526998
rect 338212 526934 338264 526940
rect 342732 526697 342760 529094
rect 347240 527066 347268 529094
rect 347228 527060 347280 527066
rect 347228 527002 347280 527008
rect 342718 526688 342774 526697
rect 342718 526623 342774 526632
rect 351932 526522 351960 529094
rect 356256 527882 356284 529094
rect 356244 527876 356296 527882
rect 356244 527818 356296 527824
rect 360764 526833 360792 529094
rect 360750 526824 360806 526833
rect 360750 526759 360806 526768
rect 365272 526590 365300 529094
rect 365260 526584 365312 526590
rect 365260 526526 365312 526532
rect 351920 526516 351972 526522
rect 351920 526458 351972 526464
rect 369872 526454 369900 529094
rect 374288 527950 374316 529094
rect 374276 527944 374328 527950
rect 374276 527886 374328 527892
rect 379532 526726 379560 529094
rect 379520 526720 379572 526726
rect 379520 526662 379572 526668
rect 369860 526448 369912 526454
rect 369860 526390 369912 526396
rect 333980 526244 334032 526250
rect 333980 526186 334032 526192
rect 329748 524136 329800 524142
rect 329748 524078 329800 524084
rect 383672 486470 383700 529094
rect 388456 526658 388484 529094
rect 388444 526652 388496 526658
rect 388444 526594 388496 526600
rect 393332 526318 393360 529094
rect 397472 529094 397808 529122
rect 401980 529094 402316 529122
rect 406488 529094 406824 529122
rect 411332 529094 411392 529122
rect 393320 526312 393372 526318
rect 393320 526254 393372 526260
rect 397472 523705 397500 529094
rect 401980 526794 402008 529094
rect 406488 526862 406516 529094
rect 411364 528554 411392 529094
rect 411272 528526 411392 528554
rect 415596 529094 415840 529122
rect 420012 529094 420348 529122
rect 424520 529094 424856 529122
rect 429212 529094 429364 529122
rect 411272 526930 411300 528526
rect 411260 526924 411312 526930
rect 411260 526866 411312 526872
rect 406476 526856 406528 526862
rect 406476 526798 406528 526804
rect 401968 526788 402020 526794
rect 401968 526730 402020 526736
rect 415596 526386 415624 529094
rect 420012 527134 420040 529094
rect 420000 527128 420052 527134
rect 424520 527105 424548 529094
rect 420000 527070 420052 527076
rect 424506 527096 424562 527105
rect 424506 527031 424562 527040
rect 429212 526969 429240 529094
rect 429198 526960 429254 526969
rect 429198 526895 429254 526904
rect 415584 526380 415636 526386
rect 415584 526322 415636 526328
rect 433352 525570 433380 615839
rect 433430 601624 433486 601633
rect 433430 601559 433486 601568
rect 433340 525564 433392 525570
rect 433340 525506 433392 525512
rect 433444 524210 433472 601559
rect 433522 567488 433578 567497
rect 433522 567423 433578 567432
rect 433536 524278 433564 567423
rect 434626 529816 434682 529825
rect 434626 529751 434682 529760
rect 434640 524346 434668 529751
rect 434628 524340 434680 524346
rect 434628 524282 434680 524288
rect 433524 524272 433576 524278
rect 433524 524214 433576 524220
rect 433432 524204 433484 524210
rect 433432 524146 433484 524152
rect 434732 524142 434760 700402
rect 434812 700392 434864 700398
rect 434812 700334 434864 700340
rect 434824 635225 434852 700334
rect 434904 647896 434956 647902
rect 434904 647838 434956 647844
rect 434810 635216 434866 635225
rect 434810 635151 434866 635160
rect 434810 592376 434866 592385
rect 434810 592311 434866 592320
rect 434720 524136 434772 524142
rect 434720 524078 434772 524084
rect 397458 523696 397514 523705
rect 397458 523631 397514 523640
rect 383660 486464 383712 486470
rect 383660 486406 383712 486412
rect 356796 485716 356848 485722
rect 356796 485658 356848 485664
rect 356704 485512 356756 485518
rect 356704 485454 356756 485460
rect 318062 482216 318118 482225
rect 318062 482151 318118 482160
rect 299480 480072 299532 480078
rect 299480 480014 299532 480020
rect 299020 477624 299072 477630
rect 299020 477566 299072 477572
rect 298284 471708 298336 471714
rect 298284 471650 298336 471656
rect 297732 471640 297784 471646
rect 297732 471582 297784 471588
rect 296810 471336 296866 471345
rect 296810 471271 296866 471280
rect 296718 468480 296774 468489
rect 296718 468415 296774 468424
rect 338488 466608 338540 466614
rect 338486 466576 338488 466585
rect 338540 466576 338542 466585
rect 338486 466511 338542 466520
rect 339774 466576 339830 466585
rect 339774 466511 339776 466520
rect 339828 466511 339830 466520
rect 350998 466576 351054 466585
rect 350998 466511 351054 466520
rect 339776 466482 339828 466488
rect 351012 466478 351040 466511
rect 351000 466472 351052 466478
rect 351000 466414 351052 466420
rect 295432 466404 295484 466410
rect 295432 466346 295484 466352
rect 295340 464500 295392 464506
rect 295340 464442 295392 464448
rect 291200 464432 291252 464438
rect 291200 464374 291252 464380
rect 271880 464364 271932 464370
rect 271880 464306 271932 464312
rect 220084 380996 220136 381002
rect 220084 380938 220136 380944
rect 220096 379506 220124 380938
rect 248236 380928 248288 380934
rect 248234 380896 248236 380905
rect 248288 380896 248290 380905
rect 220728 380860 220780 380866
rect 248234 380831 248290 380840
rect 220728 380802 220780 380808
rect 220084 379500 220136 379506
rect 220084 379442 220136 379448
rect 220096 378486 220124 379442
rect 220176 379228 220228 379234
rect 220176 379170 220228 379176
rect 220188 378690 220216 379170
rect 220740 378894 220768 380802
rect 235998 380624 236054 380633
rect 235998 380559 236054 380568
rect 237102 380624 237158 380633
rect 237102 380559 237158 380568
rect 243082 380624 243138 380633
rect 243082 380559 243138 380568
rect 245382 380624 245438 380633
rect 245382 380559 245438 380568
rect 247590 380624 247646 380633
rect 247590 380559 247646 380568
rect 254490 380624 254546 380633
rect 254490 380559 254546 380568
rect 255870 380624 255926 380633
rect 255870 380559 255926 380568
rect 256974 380624 257030 380633
rect 256974 380559 257030 380568
rect 258078 380624 258134 380633
rect 258078 380559 258134 380568
rect 259458 380624 259514 380633
rect 259458 380559 259514 380568
rect 265254 380624 265310 380633
rect 265254 380559 265310 380568
rect 265530 380624 265586 380633
rect 265530 380559 265586 380568
rect 270958 380624 271014 380633
rect 270958 380559 271014 380568
rect 222016 380384 222068 380390
rect 222016 380326 222068 380332
rect 221004 379092 221056 379098
rect 221004 379034 221056 379040
rect 220912 378956 220964 378962
rect 220912 378898 220964 378904
rect 220728 378888 220780 378894
rect 220728 378830 220780 378836
rect 220176 378684 220228 378690
rect 220176 378626 220228 378632
rect 220084 378480 220136 378486
rect 220084 378422 220136 378428
rect 220740 378214 220768 378830
rect 220820 378480 220872 378486
rect 220820 378422 220872 378428
rect 220728 378208 220780 378214
rect 220728 378150 220780 378156
rect 220832 358766 220860 378422
rect 220924 378214 220952 378898
rect 221016 378554 221044 379034
rect 222028 378826 222056 380326
rect 236012 380118 236040 380559
rect 236000 380112 236052 380118
rect 236000 380054 236052 380060
rect 237116 380050 237144 380559
rect 237104 380044 237156 380050
rect 237104 379986 237156 379992
rect 239128 380044 239180 380050
rect 239128 379986 239180 379992
rect 222016 378820 222068 378826
rect 222016 378762 222068 378768
rect 221004 378548 221056 378554
rect 221004 378490 221056 378496
rect 220912 378208 220964 378214
rect 220912 378150 220964 378156
rect 221016 375850 221044 378490
rect 221188 378208 221240 378214
rect 221188 378150 221240 378156
rect 220924 375822 221044 375850
rect 220820 358760 220872 358766
rect 220820 358702 220872 358708
rect 220924 357882 220952 375822
rect 221200 375442 221228 378150
rect 239140 376009 239168 379986
rect 243096 379982 243124 380559
rect 243084 379976 243136 379982
rect 243084 379918 243136 379924
rect 245396 378826 245424 380559
rect 246210 379400 246266 379409
rect 246210 379335 246266 379344
rect 245384 378820 245436 378826
rect 245384 378762 245436 378768
rect 246224 378350 246252 379335
rect 247604 378894 247632 380559
rect 254504 379914 254532 380559
rect 254492 379908 254544 379914
rect 254492 379850 254544 379856
rect 255884 379778 255912 380559
rect 256988 379846 257016 380559
rect 256976 379840 257028 379846
rect 256976 379782 257028 379788
rect 255872 379772 255924 379778
rect 255872 379714 255924 379720
rect 258092 379710 258120 380559
rect 259472 380050 259500 380559
rect 259460 380044 259512 380050
rect 259460 379986 259512 379992
rect 258080 379704 258132 379710
rect 258080 379646 258132 379652
rect 263876 379636 263928 379642
rect 263876 379578 263928 379584
rect 263888 379409 263916 379578
rect 265268 379574 265296 380559
rect 265256 379568 265308 379574
rect 265256 379510 265308 379516
rect 248602 379400 248658 379409
rect 248602 379335 248658 379344
rect 250074 379400 250130 379409
rect 250074 379335 250130 379344
rect 251178 379400 251234 379409
rect 251178 379335 251234 379344
rect 252282 379400 252338 379409
rect 252282 379335 252338 379344
rect 253386 379400 253442 379409
rect 253386 379335 253442 379344
rect 261666 379400 261722 379409
rect 261666 379335 261722 379344
rect 263874 379400 263930 379409
rect 263874 379335 263930 379344
rect 247592 378888 247644 378894
rect 247592 378830 247644 378836
rect 248616 378690 248644 379335
rect 248604 378684 248656 378690
rect 248604 378626 248656 378632
rect 250088 378622 250116 379335
rect 250076 378616 250128 378622
rect 250076 378558 250128 378564
rect 251192 378554 251220 379335
rect 251180 378548 251232 378554
rect 251180 378490 251232 378496
rect 252296 378486 252324 379335
rect 253110 379128 253166 379137
rect 253110 379063 253166 379072
rect 252284 378480 252336 378486
rect 253124 378457 253152 379063
rect 252284 378422 252336 378428
rect 253110 378448 253166 378457
rect 253110 378383 253166 378392
rect 246212 378344 246264 378350
rect 244278 378312 244334 378321
rect 246212 378286 246264 378292
rect 250626 378312 250682 378321
rect 244278 378247 244334 378256
rect 250626 378247 250682 378256
rect 239126 376000 239182 376009
rect 239126 375935 239182 375944
rect 221016 375414 221228 375442
rect 221016 358698 221044 375414
rect 244292 375018 244320 378247
rect 250640 376106 250668 378247
rect 253400 378214 253428 379335
rect 253570 378584 253626 378593
rect 253570 378519 253626 378528
rect 255962 378584 256018 378593
rect 255962 378519 256018 378528
rect 258354 378584 258410 378593
rect 258354 378519 258410 378528
rect 260930 378584 260986 378593
rect 260930 378519 260986 378528
rect 253388 378208 253440 378214
rect 253388 378150 253440 378156
rect 250628 376100 250680 376106
rect 250628 376042 250680 376048
rect 253584 375834 253612 378519
rect 255976 375902 256004 378519
rect 258368 375970 258396 378519
rect 260944 376038 260972 378519
rect 260932 376032 260984 376038
rect 260932 375974 260984 375980
rect 258356 375964 258408 375970
rect 258356 375906 258408 375912
rect 255964 375896 256016 375902
rect 255964 375838 256016 375844
rect 253572 375828 253624 375834
rect 253572 375770 253624 375776
rect 244280 375012 244332 375018
rect 244280 374954 244332 374960
rect 261680 374950 261708 379335
rect 263598 378584 263654 378593
rect 263598 378519 263654 378528
rect 262770 378312 262826 378321
rect 262770 378247 262826 378256
rect 261668 374944 261720 374950
rect 261668 374886 261720 374892
rect 262784 374882 262812 378247
rect 263612 376174 263640 378519
rect 265544 378457 265572 380559
rect 268658 379400 268714 379409
rect 268658 379335 268714 379344
rect 265898 378584 265954 378593
rect 265898 378519 265954 378528
rect 268106 378584 268162 378593
rect 268106 378519 268162 378528
rect 265530 378448 265586 378457
rect 265530 378383 265586 378392
rect 265912 376242 265940 378519
rect 266358 378312 266414 378321
rect 266358 378247 266414 378256
rect 267554 378312 267610 378321
rect 267554 378247 267610 378256
rect 265900 376236 265952 376242
rect 265900 376178 265952 376184
rect 263600 376168 263652 376174
rect 263600 376110 263652 376116
rect 262772 374876 262824 374882
rect 262772 374818 262824 374824
rect 266372 374746 266400 378247
rect 267568 374814 267596 378247
rect 268120 376310 268148 378519
rect 268672 378418 268700 379335
rect 268660 378412 268712 378418
rect 268660 378354 268712 378360
rect 270972 376378 271000 380559
rect 295340 380316 295392 380322
rect 295340 380258 295392 380264
rect 275652 379500 275704 379506
rect 275652 379442 275704 379448
rect 274364 379432 274416 379438
rect 271050 379400 271106 379409
rect 271050 379335 271106 379344
rect 272154 379400 272210 379409
rect 272154 379335 272210 379344
rect 273258 379400 273314 379409
rect 273258 379335 273260 379344
rect 271064 379302 271092 379335
rect 271052 379296 271104 379302
rect 271052 379238 271104 379244
rect 272168 379030 272196 379335
rect 273312 379335 273314 379344
rect 274362 379400 274364 379409
rect 275664 379409 275692 379442
rect 274416 379400 274418 379409
rect 274362 379335 274418 379344
rect 275650 379400 275706 379409
rect 275650 379335 275706 379344
rect 276110 379400 276166 379409
rect 276110 379335 276166 379344
rect 277030 379400 277086 379409
rect 277030 379335 277086 379344
rect 278226 379400 278282 379409
rect 278226 379335 278282 379344
rect 285954 379400 286010 379409
rect 285954 379335 286010 379344
rect 287610 379400 287666 379409
rect 287610 379335 287666 379344
rect 290922 379400 290978 379409
rect 290922 379335 290978 379344
rect 292670 379400 292726 379409
rect 295352 379370 295380 380258
rect 301504 380248 301556 380254
rect 301504 380190 301556 380196
rect 301516 379506 301544 380190
rect 310428 380180 310480 380186
rect 310428 380122 310480 380128
rect 301504 379500 301556 379506
rect 301504 379442 301556 379448
rect 310440 379438 310468 380122
rect 313372 379500 313424 379506
rect 313372 379442 313424 379448
rect 310428 379432 310480 379438
rect 295430 379400 295486 379409
rect 292670 379335 292726 379344
rect 295340 379364 295392 379370
rect 273260 379306 273312 379312
rect 272156 379024 272208 379030
rect 272156 378966 272208 378972
rect 273442 378584 273498 378593
rect 273442 378519 273498 378528
rect 273260 378344 273312 378350
rect 273260 378286 273312 378292
rect 271788 378208 271840 378214
rect 271788 378150 271840 378156
rect 271800 377398 271828 378150
rect 273272 377466 273300 378286
rect 273260 377460 273312 377466
rect 273260 377402 273312 377408
rect 271788 377392 271840 377398
rect 271788 377334 271840 377340
rect 273456 376446 273484 378519
rect 276020 378276 276072 378282
rect 276020 378218 276072 378224
rect 276032 378185 276060 378218
rect 276018 378176 276074 378185
rect 276018 378111 276074 378120
rect 276124 376514 276152 379335
rect 277044 378282 277072 379335
rect 277032 378276 277084 378282
rect 277032 378218 277084 378224
rect 278240 377534 278268 379335
rect 280250 379264 280306 379273
rect 280250 379199 280306 379208
rect 283378 379264 283434 379273
rect 283378 379199 283434 379208
rect 278228 377528 278280 377534
rect 278228 377470 278280 377476
rect 280264 377330 280292 379199
rect 280252 377324 280304 377330
rect 280252 377266 280304 377272
rect 283392 376650 283420 379199
rect 285968 377602 285996 379335
rect 287624 378146 287652 379335
rect 287612 378140 287664 378146
rect 287612 378082 287664 378088
rect 290936 377670 290964 379335
rect 292684 377874 292712 379335
rect 295430 379335 295486 379344
rect 298466 379400 298522 379409
rect 298466 379335 298522 379344
rect 300858 379400 300914 379409
rect 300858 379335 300914 379344
rect 303250 379400 303306 379409
rect 303250 379335 303306 379344
rect 305826 379400 305882 379409
rect 305826 379335 305882 379344
rect 307850 379400 307906 379409
rect 313384 379409 313412 379442
rect 315764 379432 315816 379438
rect 310428 379374 310480 379380
rect 310978 379400 311034 379409
rect 307850 379335 307906 379344
rect 310978 379335 310980 379344
rect 295340 379306 295392 379312
rect 295444 377942 295472 379335
rect 298480 378010 298508 379335
rect 300872 378350 300900 379335
rect 300860 378344 300912 378350
rect 300860 378286 300912 378292
rect 298468 378004 298520 378010
rect 298468 377946 298520 377952
rect 295432 377936 295484 377942
rect 295432 377878 295484 377884
rect 292672 377868 292724 377874
rect 292672 377810 292724 377816
rect 303264 377738 303292 379335
rect 305840 378214 305868 379335
rect 305828 378208 305880 378214
rect 305828 378150 305880 378156
rect 307864 377806 307892 379335
rect 311032 379335 311034 379344
rect 313370 379400 313426 379409
rect 313370 379335 313426 379344
rect 315762 379400 315764 379409
rect 315816 379400 315818 379409
rect 315762 379335 315818 379344
rect 317418 379400 317474 379409
rect 317418 379335 317474 379344
rect 310980 379306 311032 379312
rect 317432 378078 317460 379335
rect 325882 379264 325938 379273
rect 325882 379199 325938 379208
rect 320914 378584 320970 378593
rect 320914 378519 320970 378528
rect 317420 378072 317472 378078
rect 317420 378014 317472 378020
rect 307852 377800 307904 377806
rect 307852 377742 307904 377748
rect 303252 377732 303304 377738
rect 303252 377674 303304 377680
rect 290924 377664 290976 377670
rect 290924 377606 290976 377612
rect 285956 377596 286008 377602
rect 285956 377538 286008 377544
rect 283380 376644 283432 376650
rect 283380 376586 283432 376592
rect 320928 376582 320956 378519
rect 320916 376576 320968 376582
rect 320916 376518 320968 376524
rect 276112 376508 276164 376514
rect 276112 376450 276164 376456
rect 273444 376440 273496 376446
rect 273444 376382 273496 376388
rect 270960 376372 271012 376378
rect 270960 376314 271012 376320
rect 268108 376304 268160 376310
rect 268108 376246 268160 376252
rect 325896 375766 325924 379199
rect 343178 378448 343234 378457
rect 343178 378383 343234 378392
rect 343192 378350 343220 378383
rect 342260 378344 342312 378350
rect 342260 378286 342312 378292
rect 343180 378344 343232 378350
rect 343180 378286 343232 378292
rect 343546 378312 343602 378321
rect 325884 375760 325936 375766
rect 325884 375702 325936 375708
rect 267556 374808 267608 374814
rect 267556 374750 267608 374756
rect 266360 374740 266412 374746
rect 266360 374682 266412 374688
rect 342272 374678 342300 378286
rect 343546 378247 343602 378256
rect 356612 378276 356664 378282
rect 343560 378214 343588 378247
rect 356612 378218 356664 378224
rect 343548 378208 343600 378214
rect 343548 378150 343600 378156
rect 342260 374672 342312 374678
rect 342260 374614 342312 374620
rect 340052 359644 340104 359650
rect 340052 359586 340104 359592
rect 338488 359576 338540 359582
rect 338488 359518 338540 359524
rect 338500 358873 338528 359518
rect 340064 358873 340092 359586
rect 338486 358864 338542 358873
rect 338486 358799 338542 358808
rect 340050 358864 340106 358873
rect 343560 358834 343588 378150
rect 351736 359508 351788 359514
rect 351736 359450 351788 359456
rect 351748 358873 351776 359450
rect 351734 358864 351790 358873
rect 340050 358799 340106 358808
rect 342260 358828 342312 358834
rect 342260 358770 342312 358776
rect 343548 358828 343600 358834
rect 351734 358799 351790 358808
rect 343548 358770 343600 358776
rect 221004 358692 221056 358698
rect 221004 358634 221056 358640
rect 342272 358086 342300 358770
rect 342260 358080 342312 358086
rect 342260 358022 342312 358028
rect 220912 357876 220964 357882
rect 220912 357818 220964 357824
rect 266358 273592 266414 273601
rect 266358 273527 266414 273536
rect 283470 273592 283526 273601
rect 283470 273527 283526 273536
rect 266372 273426 266400 273527
rect 273258 273456 273314 273465
rect 266360 273420 266412 273426
rect 273258 273391 273314 273400
rect 266360 273362 266412 273368
rect 273272 273358 273300 273391
rect 273260 273352 273312 273358
rect 273260 273294 273312 273300
rect 283484 273290 283512 273527
rect 283472 273284 283524 273290
rect 283472 273226 283524 273232
rect 288164 273080 288216 273086
rect 288164 273022 288216 273028
rect 285956 273012 286008 273018
rect 285956 272954 286008 272960
rect 285968 272921 285996 272954
rect 288176 272921 288204 273022
rect 295892 272944 295944 272950
rect 285954 272912 286010 272921
rect 285954 272847 286010 272856
rect 288162 272912 288218 272921
rect 288162 272847 288218 272856
rect 290922 272912 290978 272921
rect 290922 272847 290924 272856
rect 290976 272847 290978 272856
rect 295890 272912 295892 272921
rect 295944 272912 295946 272921
rect 295890 272847 295946 272856
rect 303434 272912 303490 272921
rect 303434 272847 303490 272856
rect 290924 272818 290976 272824
rect 303448 272814 303476 272847
rect 303436 272808 303488 272814
rect 298466 272776 298522 272785
rect 298466 272711 298468 272720
rect 298520 272711 298522 272720
rect 300858 272776 300914 272785
rect 303436 272750 303488 272756
rect 300858 272711 300914 272720
rect 298468 272682 298520 272688
rect 300872 272678 300900 272711
rect 300860 272672 300912 272678
rect 300860 272614 300912 272620
rect 305826 272640 305882 272649
rect 305826 272575 305828 272584
rect 305880 272575 305882 272584
rect 320914 272640 320970 272649
rect 320914 272575 320970 272584
rect 305828 272546 305880 272552
rect 320928 272542 320956 272575
rect 320916 272536 320968 272542
rect 320916 272478 320968 272484
rect 265162 272232 265218 272241
rect 265162 272167 265218 272176
rect 263598 271824 263654 271833
rect 263598 271759 263654 271768
rect 264978 271824 265034 271833
rect 264978 271759 265034 271768
rect 263612 271522 263640 271759
rect 263600 271516 263652 271522
rect 263600 271458 263652 271464
rect 264992 271318 265020 271759
rect 264980 271312 265032 271318
rect 258262 271280 258318 271289
rect 258262 271215 258318 271224
rect 260838 271280 260894 271289
rect 264980 271254 265032 271260
rect 260838 271215 260840 271224
rect 258276 271182 258304 271215
rect 260892 271215 260894 271224
rect 260840 271186 260892 271192
rect 258264 271176 258316 271182
rect 247038 271144 247094 271153
rect 247038 271079 247094 271088
rect 252558 271144 252614 271153
rect 252558 271079 252560 271088
rect 247052 270978 247080 271079
rect 252612 271079 252614 271088
rect 255318 271144 255374 271153
rect 258264 271118 258316 271124
rect 255318 271079 255374 271088
rect 252560 271050 252612 271056
rect 255332 271046 255360 271079
rect 255320 271040 255372 271046
rect 255320 270982 255372 270988
rect 247040 270972 247092 270978
rect 247040 270914 247092 270920
rect 253938 270872 253994 270881
rect 253938 270807 253994 270816
rect 244370 270736 244426 270745
rect 244370 270671 244426 270680
rect 251270 270736 251326 270745
rect 251270 270671 251326 270680
rect 237378 270600 237434 270609
rect 237378 270535 237434 270544
rect 242898 270600 242954 270609
rect 242898 270535 242954 270544
rect 244278 270600 244334 270609
rect 244278 270535 244334 270544
rect 220544 270496 220596 270502
rect 220544 270438 220596 270444
rect 220360 270020 220412 270026
rect 220360 269962 220412 269968
rect 220372 269482 220400 269962
rect 220556 269550 220584 270438
rect 220728 270428 220780 270434
rect 220728 270370 220780 270376
rect 220740 270065 220768 270370
rect 220726 270056 220782 270065
rect 220726 269991 220782 270000
rect 220636 269952 220688 269958
rect 220636 269894 220688 269900
rect 220544 269544 220596 269550
rect 220544 269486 220596 269492
rect 220360 269476 220412 269482
rect 220360 269418 220412 269424
rect 220648 269278 220676 269894
rect 220728 269884 220780 269890
rect 220728 269826 220780 269832
rect 220740 269414 220768 269826
rect 237392 269754 237420 270535
rect 237380 269748 237432 269754
rect 237380 269690 237432 269696
rect 220728 269408 220780 269414
rect 220728 269350 220780 269356
rect 220636 269272 220688 269278
rect 220636 269214 220688 269220
rect 232504 268932 232556 268938
rect 232504 268874 232556 268880
rect 231124 268864 231176 268870
rect 231124 268806 231176 268812
rect 229100 268796 229152 268802
rect 229100 268738 229152 268744
rect 229112 251870 229140 268738
rect 231136 252550 231164 268806
rect 231124 252544 231176 252550
rect 231124 252486 231176 252492
rect 232516 252482 232544 268874
rect 242912 268326 242940 270535
rect 244292 270094 244320 270535
rect 244280 270088 244332 270094
rect 244280 270030 244332 270036
rect 242900 268320 242952 268326
rect 242900 268262 242952 268268
rect 244384 268258 244412 270671
rect 245658 270600 245714 270609
rect 245658 270535 245714 270544
rect 247038 270600 247094 270609
rect 247038 270535 247094 270544
rect 248510 270600 248566 270609
rect 248510 270535 248566 270544
rect 249798 270600 249854 270609
rect 249798 270535 249854 270544
rect 251178 270600 251234 270609
rect 251178 270535 251234 270544
rect 245672 270298 245700 270535
rect 247052 270434 247080 270535
rect 248524 270502 248552 270535
rect 248512 270496 248564 270502
rect 248512 270438 248564 270444
rect 247040 270428 247092 270434
rect 247040 270370 247092 270376
rect 245660 270292 245712 270298
rect 245660 270234 245712 270240
rect 249812 270026 249840 270535
rect 251192 270230 251220 270535
rect 251180 270224 251232 270230
rect 251180 270166 251232 270172
rect 251284 270162 251312 270671
rect 252558 270600 252614 270609
rect 252558 270535 252614 270544
rect 252572 270366 252600 270535
rect 252560 270360 252612 270366
rect 252560 270302 252612 270308
rect 251272 270156 251324 270162
rect 251272 270098 251324 270104
rect 249800 270020 249852 270026
rect 249800 269962 249852 269968
rect 253952 269006 253980 270807
rect 255318 270736 255374 270745
rect 255318 270671 255374 270680
rect 259550 270736 259606 270745
rect 259550 270671 259606 270680
rect 253940 269000 253992 269006
rect 253940 268942 253992 268948
rect 255332 268734 255360 270671
rect 256698 270600 256754 270609
rect 256698 270535 256754 270544
rect 258078 270600 258134 270609
rect 258078 270535 258134 270544
rect 259458 270600 259514 270609
rect 259458 270535 259514 270544
rect 255320 268728 255372 268734
rect 255320 268670 255372 268676
rect 256712 268666 256740 270535
rect 256700 268660 256752 268666
rect 256700 268602 256752 268608
rect 258092 268598 258120 270535
rect 259472 268938 259500 270535
rect 259460 268932 259512 268938
rect 259460 268874 259512 268880
rect 259564 268870 259592 270671
rect 260838 270600 260894 270609
rect 260838 270535 260894 270544
rect 262218 270600 262274 270609
rect 262218 270535 262274 270544
rect 263598 270600 263654 270609
rect 263598 270535 263654 270544
rect 259552 268864 259604 268870
rect 259552 268806 259604 268812
rect 260852 268802 260880 270535
rect 262232 269958 262260 270535
rect 262220 269952 262272 269958
rect 262220 269894 262272 269900
rect 263612 269618 263640 270535
rect 265176 269890 265204 272167
rect 313280 271856 313332 271862
rect 268014 271824 268070 271833
rect 268014 271759 268070 271768
rect 270498 271824 270554 271833
rect 270498 271759 270554 271768
rect 271878 271824 271934 271833
rect 271878 271759 271934 271768
rect 276018 271824 276074 271833
rect 276018 271759 276074 271768
rect 277950 271824 278006 271833
rect 277950 271759 278006 271768
rect 280066 271824 280122 271833
rect 280066 271759 280122 271768
rect 280250 271824 280306 271833
rect 280250 271759 280306 271768
rect 307758 271824 307814 271833
rect 307758 271759 307760 271768
rect 268028 271386 268056 271759
rect 270512 271658 270540 271759
rect 270500 271652 270552 271658
rect 270500 271594 270552 271600
rect 268016 271380 268068 271386
rect 268016 271322 268068 271328
rect 270498 271280 270554 271289
rect 270498 271215 270554 271224
rect 267922 270872 267978 270881
rect 267922 270807 267978 270816
rect 266358 270600 266414 270609
rect 266358 270535 266414 270544
rect 265164 269884 265216 269890
rect 265164 269826 265216 269832
rect 266372 269822 266400 270535
rect 266360 269816 266412 269822
rect 266360 269758 266412 269764
rect 263600 269612 263652 269618
rect 263600 269554 263652 269560
rect 267936 269074 267964 270807
rect 269118 270600 269174 270609
rect 269118 270535 269174 270544
rect 267924 269068 267976 269074
rect 267924 269010 267976 269016
rect 260840 268796 260892 268802
rect 260840 268738 260892 268744
rect 258080 268592 258132 268598
rect 258080 268534 258132 268540
rect 269132 268530 269160 270535
rect 269120 268524 269172 268530
rect 269120 268466 269172 268472
rect 270512 268462 270540 271215
rect 271892 269686 271920 271759
rect 276032 271590 276060 271759
rect 276020 271584 276072 271590
rect 276020 271526 276072 271532
rect 277214 271552 277270 271561
rect 277214 271487 277270 271496
rect 277228 271182 277256 271487
rect 277964 271454 277992 271759
rect 277952 271448 278004 271454
rect 277952 271390 278004 271396
rect 280080 271250 280108 271759
rect 280264 271726 280292 271759
rect 307812 271759 307814 271768
rect 313278 271824 313280 271833
rect 313332 271824 313334 271833
rect 313278 271759 313334 271768
rect 307760 271730 307812 271736
rect 280252 271720 280304 271726
rect 280252 271662 280304 271668
rect 343546 271552 343602 271561
rect 343546 271487 343602 271496
rect 343560 271454 343588 271487
rect 343548 271448 343600 271454
rect 343454 271416 343510 271425
rect 343548 271390 343600 271396
rect 343454 271351 343510 271360
rect 343468 271318 343496 271351
rect 343456 271312 343508 271318
rect 343456 271254 343508 271260
rect 280068 271244 280120 271250
rect 280068 271186 280120 271192
rect 356624 271182 356652 378218
rect 277216 271176 277268 271182
rect 277216 271118 277268 271124
rect 356612 271176 356664 271182
rect 356612 271118 356664 271124
rect 277398 270872 277454 270881
rect 277398 270807 277454 270816
rect 273166 270600 273222 270609
rect 273166 270535 273222 270544
rect 274638 270600 274694 270609
rect 274638 270535 274694 270544
rect 271880 269680 271932 269686
rect 271880 269622 271932 269628
rect 270500 268456 270552 268462
rect 270500 268398 270552 268404
rect 273180 268394 273208 270535
rect 273168 268388 273220 268394
rect 273168 268330 273220 268336
rect 244372 268252 244424 268258
rect 244372 268194 244424 268200
rect 274652 267714 274680 270535
rect 274640 267708 274692 267714
rect 274640 267650 274692 267656
rect 277412 267646 277440 270807
rect 277400 267640 277452 267646
rect 277400 267582 277452 267588
rect 339408 253904 339460 253910
rect 339408 253846 339460 253852
rect 339420 253609 339448 253846
rect 339406 253600 339462 253609
rect 339406 253535 339462 253544
rect 340788 253292 340840 253298
rect 340788 253234 340840 253240
rect 340800 253065 340828 253234
rect 351828 253224 351880 253230
rect 351826 253192 351828 253201
rect 351880 253192 351882 253201
rect 351826 253127 351882 253136
rect 340786 253056 340842 253065
rect 340786 252991 340842 253000
rect 232504 252476 232556 252482
rect 232504 252418 232556 252424
rect 229100 251864 229152 251870
rect 229100 251806 229152 251812
rect 220820 166796 220872 166802
rect 220820 166738 220872 166744
rect 220832 146169 220860 166738
rect 260932 166728 260984 166734
rect 260932 166670 260984 166676
rect 303526 166696 303582 166705
rect 260944 166433 260972 166670
rect 265900 166660 265952 166666
rect 303526 166631 303582 166640
rect 265900 166602 265952 166608
rect 265912 166433 265940 166602
rect 293408 166592 293460 166598
rect 285954 166560 286010 166569
rect 285954 166495 285956 166504
rect 286008 166495 286010 166504
rect 288254 166560 288310 166569
rect 288254 166495 288310 166504
rect 293406 166560 293408 166569
rect 293460 166560 293462 166569
rect 293406 166495 293462 166504
rect 295890 166560 295946 166569
rect 295890 166495 295946 166504
rect 285956 166466 286008 166472
rect 288268 166462 288296 166495
rect 288256 166456 288308 166462
rect 260930 166424 260986 166433
rect 260930 166359 260986 166368
rect 265898 166424 265954 166433
rect 288256 166398 288308 166404
rect 295904 166394 295932 166495
rect 265898 166359 265954 166368
rect 295892 166388 295944 166394
rect 295892 166330 295944 166336
rect 303540 166326 303568 166631
rect 303528 166320 303580 166326
rect 303528 166262 303580 166268
rect 235998 165608 236054 165617
rect 235998 165543 236054 165552
rect 238758 165608 238814 165617
rect 238758 165543 238814 165552
rect 242898 165608 242954 165617
rect 242898 165543 242954 165552
rect 247038 165608 247094 165617
rect 247038 165543 247094 165552
rect 247682 165608 247738 165617
rect 247682 165543 247738 165552
rect 249798 165608 249854 165617
rect 249798 165543 249854 165552
rect 252558 165608 252614 165617
rect 252558 165543 252614 165552
rect 258078 165608 258134 165617
rect 258078 165543 258134 165552
rect 260838 165608 260894 165617
rect 260838 165543 260894 165552
rect 264978 165608 265034 165617
rect 264978 165543 265034 165552
rect 267738 165608 267794 165617
rect 267738 165543 267794 165552
rect 271878 165608 271934 165617
rect 271878 165543 271934 165552
rect 273442 165608 273498 165617
rect 273442 165543 273498 165552
rect 275926 165608 275982 165617
rect 276202 165608 276258 165617
rect 275982 165566 276152 165594
rect 275926 165543 275982 165552
rect 236012 164082 236040 165543
rect 236090 164248 236146 164257
rect 236090 164183 236146 164192
rect 237378 164248 237434 164257
rect 237378 164183 237434 164192
rect 236000 164076 236052 164082
rect 236000 164018 236052 164024
rect 235264 161560 235316 161566
rect 235264 161502 235316 161508
rect 235276 146198 235304 161502
rect 235264 146192 235316 146198
rect 220818 146160 220874 146169
rect 235264 146134 235316 146140
rect 220818 146095 220874 146104
rect 236012 145450 236040 164018
rect 236104 164014 236132 164183
rect 236092 164008 236144 164014
rect 236092 163950 236144 163956
rect 236104 145518 236132 163950
rect 236644 161492 236696 161498
rect 236644 161434 236696 161440
rect 236656 146266 236684 161434
rect 236644 146260 236696 146266
rect 236644 146202 236696 146208
rect 237392 145761 237420 164183
rect 238772 148578 238800 165543
rect 240138 164248 240194 164257
rect 240138 164183 240194 164192
rect 241518 164248 241574 164257
rect 241518 164183 241574 164192
rect 238760 148572 238812 148578
rect 238760 148514 238812 148520
rect 240152 148510 240180 164183
rect 241532 148782 241560 164183
rect 241520 148776 241572 148782
rect 241520 148718 241572 148724
rect 240140 148504 240192 148510
rect 240140 148446 240192 148452
rect 242912 145858 242940 165543
rect 244370 164520 244426 164529
rect 244370 164455 244426 164464
rect 244278 164248 244334 164257
rect 244278 164183 244334 164192
rect 242900 145852 242952 145858
rect 242900 145794 242952 145800
rect 237378 145752 237434 145761
rect 237378 145687 237434 145696
rect 244292 145654 244320 164183
rect 244384 145790 244412 164455
rect 245658 164248 245714 164257
rect 245658 164183 245714 164192
rect 244372 145784 244424 145790
rect 244372 145726 244424 145732
rect 245672 145722 245700 164183
rect 247052 145926 247080 165543
rect 247696 164898 247724 165543
rect 249812 164966 249840 165543
rect 252572 165034 252600 165543
rect 258092 165102 258120 165543
rect 258080 165096 258132 165102
rect 258080 165038 258132 165044
rect 252560 165028 252612 165034
rect 252560 164970 252612 164976
rect 249800 164960 249852 164966
rect 249800 164902 249852 164908
rect 247684 164892 247736 164898
rect 247684 164834 247736 164840
rect 251270 164520 251326 164529
rect 251270 164455 251326 164464
rect 259550 164520 259606 164529
rect 259550 164455 259606 164464
rect 248418 164248 248474 164257
rect 248418 164183 248474 164192
rect 249798 164248 249854 164257
rect 249798 164183 249854 164192
rect 251178 164248 251234 164257
rect 251178 164183 251234 164192
rect 247040 145920 247092 145926
rect 247040 145862 247092 145868
rect 245660 145716 245712 145722
rect 245660 145658 245712 145664
rect 244280 145648 244332 145654
rect 244280 145590 244332 145596
rect 248432 145586 248460 164183
rect 249812 146062 249840 164183
rect 249800 146056 249852 146062
rect 249800 145998 249852 146004
rect 251192 145994 251220 164183
rect 251180 145988 251232 145994
rect 251180 145930 251232 145936
rect 248420 145580 248472 145586
rect 248420 145522 248472 145528
rect 236092 145512 236144 145518
rect 236092 145454 236144 145460
rect 236000 145444 236052 145450
rect 236000 145386 236052 145392
rect 251284 145314 251312 164455
rect 252558 164248 252614 164257
rect 252558 164183 252614 164192
rect 253938 164248 253994 164257
rect 253938 164183 253994 164192
rect 255318 164248 255374 164257
rect 255318 164183 255374 164192
rect 256698 164248 256754 164257
rect 256698 164183 256754 164192
rect 258078 164248 258134 164257
rect 258078 164183 258134 164192
rect 259458 164248 259514 164257
rect 259458 164183 259514 164192
rect 252572 146130 252600 164183
rect 252560 146124 252612 146130
rect 252560 146066 252612 146072
rect 253952 145382 253980 164183
rect 255332 146198 255360 164183
rect 256712 146266 256740 164183
rect 258092 162654 258120 164183
rect 259472 162722 259500 164183
rect 259564 162790 259592 164455
rect 260852 162858 260880 165543
rect 263506 164248 263562 164257
rect 263782 164248 263838 164257
rect 263562 164206 263640 164234
rect 263506 164183 263562 164192
rect 260840 162852 260892 162858
rect 260840 162794 260892 162800
rect 259552 162784 259604 162790
rect 259552 162726 259604 162732
rect 259460 162716 259512 162722
rect 259460 162658 259512 162664
rect 258080 162648 258132 162654
rect 258080 162590 258132 162596
rect 256700 146260 256752 146266
rect 256700 146202 256752 146208
rect 255320 146192 255372 146198
rect 255320 146134 255372 146140
rect 263612 146033 263640 164206
rect 263782 164183 263838 164192
rect 263796 163538 263824 164183
rect 264992 164150 265020 165543
rect 267752 165306 267780 165543
rect 267740 165300 267792 165306
rect 267740 165242 267792 165248
rect 266358 164656 266414 164665
rect 266358 164591 266414 164600
rect 264980 164144 265032 164150
rect 264980 164086 265032 164092
rect 263784 163532 263836 163538
rect 263784 163474 263836 163480
rect 266372 162178 266400 164591
rect 267646 164520 267702 164529
rect 267702 164478 267780 164506
rect 267646 164455 267702 164464
rect 266360 162172 266412 162178
rect 266360 162114 266412 162120
rect 267752 146305 267780 164478
rect 267830 164248 267886 164257
rect 267830 164183 267886 164192
rect 269118 164248 269174 164257
rect 269118 164183 269174 164192
rect 270498 164248 270554 164257
rect 270498 164183 270554 164192
rect 267738 146296 267794 146305
rect 267738 146231 267794 146240
rect 267844 146169 267872 164183
rect 267830 146160 267886 146169
rect 267830 146095 267886 146104
rect 263598 146024 263654 146033
rect 263598 145959 263654 145968
rect 269132 145625 269160 164183
rect 270512 148442 270540 164183
rect 270500 148436 270552 148442
rect 270500 148378 270552 148384
rect 271892 148374 271920 165543
rect 273456 165238 273484 165543
rect 273444 165232 273496 165238
rect 273444 165174 273496 165180
rect 274454 164520 274510 164529
rect 274454 164455 274510 164464
rect 274468 164098 274496 164455
rect 274546 164248 274602 164257
rect 276018 164248 276074 164257
rect 274602 164206 274772 164234
rect 274546 164183 274602 164192
rect 274468 164070 274680 164098
rect 274652 148850 274680 164070
rect 274744 148986 274772 164206
rect 276018 164183 276074 164192
rect 274732 148980 274784 148986
rect 274732 148922 274784 148928
rect 274640 148844 274692 148850
rect 274640 148786 274692 148792
rect 271880 148368 271932 148374
rect 271880 148310 271932 148316
rect 276032 146334 276060 164183
rect 276124 149054 276152 165566
rect 276202 165543 276258 165552
rect 277398 165608 277454 165617
rect 277398 165543 277454 165552
rect 280066 165608 280122 165617
rect 280066 165543 280122 165552
rect 280250 165608 280306 165617
rect 280250 165543 280306 165552
rect 283378 165608 283434 165617
rect 283378 165543 283434 165552
rect 300858 165608 300914 165617
rect 300858 165543 300860 165552
rect 276216 165170 276244 165543
rect 277412 165442 277440 165543
rect 277400 165436 277452 165442
rect 277400 165378 277452 165384
rect 276204 165164 276256 165170
rect 276204 165106 276256 165112
rect 277398 164248 277454 164257
rect 277398 164183 277454 164192
rect 276112 149048 276164 149054
rect 276112 148990 276164 148996
rect 277412 148918 277440 164183
rect 277400 148912 277452 148918
rect 277400 148854 277452 148860
rect 276020 146328 276072 146334
rect 276020 146270 276072 146276
rect 280080 145654 280108 165543
rect 280264 165510 280292 165543
rect 280252 165504 280304 165510
rect 280252 165446 280304 165452
rect 283392 165374 283420 165543
rect 300912 165543 300914 165552
rect 323306 165608 323362 165617
rect 323306 165543 323362 165552
rect 343454 165608 343510 165617
rect 343454 165543 343510 165552
rect 300860 165514 300912 165520
rect 283380 165368 283432 165374
rect 283380 165310 283432 165316
rect 323320 164218 323348 165543
rect 343468 165034 343496 165543
rect 343546 165472 343602 165481
rect 343546 165407 343602 165416
rect 343456 165028 343508 165034
rect 343456 164970 343508 164976
rect 343560 164898 343588 165407
rect 343548 164892 343600 164898
rect 343548 164834 343600 164840
rect 323308 164212 323360 164218
rect 323308 164154 323360 164160
rect 356624 146266 356652 271118
rect 356612 146260 356664 146266
rect 356612 146202 356664 146208
rect 338488 146192 338540 146198
rect 338488 146134 338540 146140
rect 280068 145648 280120 145654
rect 269118 145616 269174 145625
rect 280068 145590 280120 145596
rect 269118 145551 269174 145560
rect 253940 145376 253992 145382
rect 253940 145318 253992 145324
rect 251272 145308 251324 145314
rect 251272 145250 251324 145256
rect 338500 144945 338528 146134
rect 340236 146124 340288 146130
rect 340236 146066 340288 146072
rect 340248 144945 340276 146066
rect 356612 145648 356664 145654
rect 356612 145590 356664 145596
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 351642 144871 351698 144880
rect 237102 59800 237158 59809
rect 237102 59735 237158 59744
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 256974 59800 257030 59809
rect 256974 59735 257030 59744
rect 262862 59800 262918 59809
rect 262862 59735 262918 59744
rect 263874 59800 263930 59809
rect 263874 59735 263930 59744
rect 237116 59702 237144 59735
rect 237104 59696 237156 59702
rect 237104 59638 237156 59644
rect 255884 59566 255912 59735
rect 256988 59634 257016 59735
rect 258078 59664 258134 59673
rect 256976 59628 257028 59634
rect 258078 59599 258134 59608
rect 260654 59664 260710 59673
rect 260654 59599 260710 59608
rect 261758 59664 261814 59673
rect 261758 59599 261814 59608
rect 256976 59570 257028 59576
rect 255872 59560 255924 59566
rect 255872 59502 255924 59508
rect 258092 59294 258120 59599
rect 258080 59288 258132 59294
rect 258080 59230 258132 59236
rect 260668 59226 260696 59599
rect 260656 59220 260708 59226
rect 260656 59162 260708 59168
rect 261772 59158 261800 59599
rect 262876 59430 262904 59735
rect 263888 59498 263916 59735
rect 308494 59664 308550 59673
rect 308494 59599 308550 59608
rect 315854 59664 315910 59673
rect 315854 59599 315910 59608
rect 263876 59492 263928 59498
rect 263876 59434 263928 59440
rect 262864 59424 262916 59430
rect 262864 59366 262916 59372
rect 279238 59392 279294 59401
rect 279238 59327 279294 59336
rect 279252 59158 279280 59327
rect 290922 59256 290978 59265
rect 290922 59191 290978 59200
rect 300858 59256 300914 59265
rect 300858 59191 300914 59200
rect 261760 59152 261812 59158
rect 261760 59094 261812 59100
rect 279240 59152 279292 59158
rect 279240 59094 279292 59100
rect 290936 59090 290964 59191
rect 290924 59084 290976 59090
rect 290924 59026 290976 59032
rect 300872 59022 300900 59191
rect 300860 59016 300912 59022
rect 300860 58958 300912 58964
rect 308508 58886 308536 59599
rect 315868 58954 315896 59599
rect 320914 59256 320970 59265
rect 320914 59191 320970 59200
rect 325882 59256 325938 59265
rect 325882 59191 325938 59200
rect 315856 58948 315908 58954
rect 315856 58890 315908 58896
rect 308496 58880 308548 58886
rect 308496 58822 308548 58828
rect 320928 58818 320956 59191
rect 320916 58812 320968 58818
rect 320916 58754 320968 58760
rect 325896 58750 325924 59191
rect 356624 59158 356652 145590
rect 356612 59152 356664 59158
rect 356612 59094 356664 59100
rect 356716 58954 356744 485454
rect 356808 166734 356836 485658
rect 358268 485648 358320 485654
rect 358268 485590 358320 485596
rect 358176 485376 358228 485382
rect 358176 485318 358228 485324
rect 357072 481364 357124 481370
rect 357072 481306 357124 481312
rect 356888 479936 356940 479942
rect 356888 479878 356940 479884
rect 356900 273358 356928 479878
rect 356980 466608 357032 466614
rect 356980 466550 357032 466556
rect 356992 359582 357020 466550
rect 357084 380186 357112 481306
rect 357164 473952 357216 473958
rect 357164 473894 357216 473900
rect 357072 380180 357124 380186
rect 357072 380122 357124 380128
rect 357176 375970 357204 473894
rect 358084 470484 358136 470490
rect 358084 470426 358136 470432
rect 357992 467832 358044 467838
rect 357992 467774 358044 467780
rect 357532 466540 357584 466546
rect 357532 466482 357584 466488
rect 357256 466404 357308 466410
rect 357256 466346 357308 466352
rect 357164 375964 357216 375970
rect 357164 375906 357216 375912
rect 357268 374678 357296 466346
rect 357438 380216 357494 380225
rect 357438 380151 357494 380160
rect 357256 374672 357308 374678
rect 357256 374614 357308 374620
rect 356980 359576 357032 359582
rect 356980 359518 357032 359524
rect 356888 273352 356940 273358
rect 356888 273294 356940 273300
rect 356888 272128 356940 272134
rect 356888 272070 356940 272076
rect 356900 271454 356928 272070
rect 356888 271448 356940 271454
rect 356888 271390 356940 271396
rect 356796 166728 356848 166734
rect 356796 166670 356848 166676
rect 356900 165034 356928 271390
rect 356992 253978 357020 359518
rect 357452 271250 357480 380151
rect 357544 359650 357572 466482
rect 358004 380730 358032 467774
rect 358096 411942 358124 470426
rect 358084 411936 358136 411942
rect 358084 411878 358136 411884
rect 358084 389224 358136 389230
rect 358084 389166 358136 389172
rect 357992 380724 358044 380730
rect 357992 380666 358044 380672
rect 357532 359644 357584 359650
rect 357532 359586 357584 359592
rect 357440 271244 357492 271250
rect 357440 271186 357492 271192
rect 356980 253972 357032 253978
rect 356980 253914 357032 253920
rect 357452 171134 357480 271186
rect 357544 253298 357572 359586
rect 358096 359514 358124 389166
rect 358084 359508 358136 359514
rect 358084 359450 358136 359456
rect 358096 282198 358124 359450
rect 358084 282192 358136 282198
rect 358084 282134 358136 282140
rect 357808 253972 357860 253978
rect 357808 253914 357860 253920
rect 357532 253292 357584 253298
rect 357532 253234 357584 253240
rect 357716 253292 357768 253298
rect 357716 253234 357768 253240
rect 357452 171106 357572 171134
rect 357440 165640 357492 165646
rect 357440 165582 357492 165588
rect 356888 165028 356940 165034
rect 356888 164970 356940 164976
rect 356900 161474 356928 164970
rect 357452 164898 357480 165582
rect 357440 164892 357492 164898
rect 357440 164834 357492 164840
rect 356808 161446 356928 161474
rect 356704 58948 356756 58954
rect 356704 58890 356756 58896
rect 325884 58744 325936 58750
rect 325884 58686 325936 58692
rect 323308 57928 323360 57934
rect 235998 57896 236054 57905
rect 235998 57831 236054 57840
rect 237378 57896 237434 57905
rect 237378 57831 237434 57840
rect 239218 57896 239274 57905
rect 239218 57831 239274 57840
rect 240138 57896 240194 57905
rect 240138 57831 240194 57840
rect 241610 57896 241666 57905
rect 241610 57831 241666 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 245290 57896 245346 57905
rect 245290 57831 245346 57840
rect 245658 57896 245714 57905
rect 245658 57831 245714 57840
rect 247038 57896 247094 57905
rect 247038 57831 247094 57840
rect 248234 57896 248290 57905
rect 248234 57831 248290 57840
rect 248602 57896 248658 57905
rect 248602 57831 248658 57840
rect 249798 57896 249854 57905
rect 249798 57831 249854 57840
rect 251178 57896 251234 57905
rect 251178 57831 251234 57840
rect 251362 57896 251418 57905
rect 251362 57831 251418 57840
rect 253386 57896 253442 57905
rect 253386 57831 253442 57840
rect 253938 57896 253994 57905
rect 253938 57831 253994 57840
rect 258354 57896 258410 57905
rect 258354 57831 258410 57840
rect 264978 57896 265034 57905
rect 264978 57831 265034 57840
rect 266450 57896 266506 57905
rect 266450 57831 266506 57840
rect 268106 57896 268162 57905
rect 268106 57831 268162 57840
rect 268934 57896 268990 57905
rect 268934 57831 268990 57840
rect 271050 57896 271106 57905
rect 271050 57831 271106 57840
rect 271878 57896 271934 57905
rect 271878 57831 271934 57840
rect 273258 57896 273314 57905
rect 273258 57831 273314 57840
rect 275098 57896 275154 57905
rect 275098 57831 275154 57840
rect 276938 57896 276994 57905
rect 276938 57831 276994 57840
rect 278318 57896 278374 57905
rect 278318 57831 278374 57840
rect 295890 57896 295946 57905
rect 295890 57831 295946 57840
rect 298098 57896 298154 57905
rect 298098 57831 298154 57840
rect 303434 57896 303490 57905
rect 303434 57831 303490 57840
rect 305826 57896 305882 57905
rect 305826 57831 305882 57840
rect 310978 57896 311034 57905
rect 310978 57831 311034 57840
rect 313370 57896 313426 57905
rect 313370 57831 313372 57840
rect 219992 56568 220044 56574
rect 219992 56510 220044 56516
rect 236012 56438 236040 57831
rect 236000 56432 236052 56438
rect 236000 56374 236052 56380
rect 219900 56228 219952 56234
rect 219900 56170 219952 56176
rect 219808 54868 219860 54874
rect 219808 54810 219860 54816
rect 218796 54528 218848 54534
rect 218796 54470 218848 54476
rect 216312 54460 216364 54466
rect 216312 54402 216364 54408
rect 213460 54392 213512 54398
rect 213460 54334 213512 54340
rect 237392 54330 237420 57831
rect 239232 55758 239260 57831
rect 239220 55752 239272 55758
rect 239220 55694 239272 55700
rect 240152 55146 240180 57831
rect 241624 55894 241652 57831
rect 241612 55888 241664 55894
rect 241612 55830 241664 55836
rect 242912 55214 242940 57831
rect 242900 55208 242952 55214
rect 242900 55150 242952 55156
rect 240140 55140 240192 55146
rect 240140 55082 240192 55088
rect 244384 54602 244412 57831
rect 245304 55826 245332 57831
rect 245292 55820 245344 55826
rect 245292 55762 245344 55768
rect 244372 54596 244424 54602
rect 244372 54538 244424 54544
rect 245672 54534 245700 57831
rect 247052 54670 247080 57831
rect 248248 57254 248276 57831
rect 248236 57248 248288 57254
rect 248236 57190 248288 57196
rect 248616 55962 248644 57831
rect 248604 55956 248656 55962
rect 248604 55898 248656 55904
rect 249812 54738 249840 57831
rect 251192 56030 251220 57831
rect 251180 56024 251232 56030
rect 251180 55966 251232 55972
rect 251376 54806 251404 57831
rect 253400 56098 253428 57831
rect 253388 56092 253440 56098
rect 253388 56034 253440 56040
rect 253952 54874 253980 57831
rect 258368 57322 258396 57831
rect 258356 57316 258408 57322
rect 258356 57258 258408 57264
rect 264992 54942 265020 57831
rect 266358 57352 266414 57361
rect 266358 57287 266414 57296
rect 266372 56166 266400 57287
rect 266360 56160 266412 56166
rect 266360 56102 266412 56108
rect 266464 55010 266492 57831
rect 268120 56234 268148 57831
rect 268948 57633 268976 57831
rect 268934 57624 268990 57633
rect 268934 57559 268990 57568
rect 269118 57624 269174 57633
rect 269118 57559 269174 57568
rect 268108 56228 268160 56234
rect 268108 56170 268160 56176
rect 269132 55185 269160 57559
rect 271064 56302 271092 57831
rect 271052 56296 271104 56302
rect 271052 56238 271104 56244
rect 269118 55176 269174 55185
rect 269118 55111 269174 55120
rect 271892 55078 271920 57831
rect 273272 56370 273300 57831
rect 273350 57624 273406 57633
rect 273350 57559 273406 57568
rect 273260 56364 273312 56370
rect 273260 56306 273312 56312
rect 271880 55072 271932 55078
rect 271880 55014 271932 55020
rect 266452 55004 266504 55010
rect 266452 54946 266504 54952
rect 264980 54936 265032 54942
rect 264980 54878 265032 54884
rect 253940 54868 253992 54874
rect 253940 54810 253992 54816
rect 251364 54800 251416 54806
rect 251364 54742 251416 54748
rect 249800 54732 249852 54738
rect 249800 54674 249852 54680
rect 247040 54664 247092 54670
rect 247040 54606 247092 54612
rect 245660 54528 245712 54534
rect 245660 54470 245712 54476
rect 273364 54398 273392 57559
rect 275112 55690 275140 57831
rect 276952 56506 276980 57831
rect 277398 57624 277454 57633
rect 277398 57559 277454 57568
rect 276940 56500 276992 56506
rect 276940 56442 276992 56448
rect 275100 55684 275152 55690
rect 275100 55626 275152 55632
rect 277412 54466 277440 57559
rect 278332 57390 278360 57831
rect 295904 57526 295932 57831
rect 295892 57520 295944 57526
rect 295892 57462 295944 57468
rect 298112 57458 298140 57831
rect 303448 57594 303476 57831
rect 305840 57662 305868 57831
rect 310992 57730 311020 57831
rect 313424 57831 313426 57840
rect 318246 57896 318302 57905
rect 318246 57831 318302 57840
rect 323306 57896 323308 57905
rect 343180 57928 343232 57934
rect 323360 57896 323362 57905
rect 323306 57831 323362 57840
rect 343178 57896 343180 57905
rect 343232 57896 343234 57905
rect 343178 57831 343234 57840
rect 343454 57896 343510 57905
rect 356808 57866 356836 161446
rect 357544 145654 357572 171106
rect 357624 164892 357676 164898
rect 357624 164834 357676 164840
rect 357532 145648 357584 145654
rect 357532 145590 357584 145596
rect 357636 57934 357664 164834
rect 357728 146130 357756 253234
rect 357820 146198 357848 253914
rect 358096 253230 358124 282134
rect 358084 253224 358136 253230
rect 358084 253166 358136 253172
rect 358096 175982 358124 253166
rect 358084 175976 358136 175982
rect 358084 175918 358136 175924
rect 357808 146192 357860 146198
rect 357808 146134 357860 146140
rect 357716 146124 357768 146130
rect 357716 146066 357768 146072
rect 358096 145586 358124 175918
rect 358084 145580 358136 145586
rect 358084 145522 358136 145528
rect 358084 68196 358136 68202
rect 358084 68138 358136 68144
rect 358096 59362 358124 68138
rect 358188 59430 358216 485318
rect 358280 166870 358308 485590
rect 364984 485580 365036 485586
rect 364984 485522 365036 485528
rect 362224 485444 362276 485450
rect 362224 485386 362276 485392
rect 360844 485240 360896 485246
rect 360844 485182 360896 485188
rect 359464 484084 359516 484090
rect 359464 484026 359516 484032
rect 358360 481228 358412 481234
rect 358360 481170 358412 481176
rect 358372 271862 358400 481170
rect 358544 478576 358596 478582
rect 358544 478518 358596 478524
rect 358452 478508 358504 478514
rect 358452 478450 358504 478456
rect 358464 273086 358492 478450
rect 358556 377602 358584 478518
rect 358728 471912 358780 471918
rect 358728 471854 358780 471860
rect 358636 471504 358688 471510
rect 358636 471446 358688 471452
rect 358544 377596 358596 377602
rect 358544 377538 358596 377544
rect 358648 376514 358676 471446
rect 358740 378826 358768 471854
rect 358820 466472 358872 466478
rect 358820 466414 358872 466420
rect 358832 390522 358860 466414
rect 358912 465112 358964 465118
rect 358912 465054 358964 465060
rect 358924 460193 358952 465054
rect 358910 460184 358966 460193
rect 358910 460119 358966 460128
rect 358820 390516 358872 390522
rect 358820 390458 358872 390464
rect 358832 389230 358860 390458
rect 358820 389224 358872 389230
rect 358820 389166 358872 389172
rect 358728 378820 358780 378826
rect 358728 378762 358780 378768
rect 358636 376508 358688 376514
rect 358636 376450 358688 376456
rect 358820 358828 358872 358834
rect 358820 358770 358872 358776
rect 358452 273080 358504 273086
rect 358452 273022 358504 273028
rect 358832 272134 358860 358770
rect 358924 353161 358952 460119
rect 359002 400344 359058 400353
rect 359002 400279 359058 400288
rect 359016 369850 359044 400279
rect 359094 398168 359150 398177
rect 359094 398103 359150 398112
rect 359108 370530 359136 398103
rect 359186 395312 359242 395321
rect 359186 395247 359242 395256
rect 359200 371890 359228 395247
rect 359278 394088 359334 394097
rect 359278 394023 359334 394032
rect 359188 371884 359240 371890
rect 359188 371826 359240 371832
rect 359096 370524 359148 370530
rect 359096 370466 359148 370472
rect 359108 369918 359136 370466
rect 359096 369912 359148 369918
rect 359096 369854 359148 369860
rect 359004 369844 359056 369850
rect 359004 369786 359056 369792
rect 359016 366382 359044 369786
rect 359004 366376 359056 366382
rect 359004 366318 359056 366324
rect 359292 364334 359320 394023
rect 359476 391950 359504 484026
rect 359740 481432 359792 481438
rect 359740 481374 359792 481380
rect 359556 469124 359608 469130
rect 359556 469066 359608 469072
rect 359464 391944 359516 391950
rect 359464 391886 359516 391892
rect 359568 379506 359596 469066
rect 359648 469056 359700 469062
rect 359648 468998 359700 469004
rect 359660 389162 359688 468998
rect 359752 417450 359780 481374
rect 360752 473068 360804 473074
rect 360752 473010 360804 473016
rect 359924 470416 359976 470422
rect 359924 470358 359976 470364
rect 359832 470348 359884 470354
rect 359832 470290 359884 470296
rect 359740 417444 359792 417450
rect 359740 417386 359792 417392
rect 359844 409154 359872 470290
rect 359936 410582 359964 470358
rect 360660 464500 360712 464506
rect 360660 464442 360712 464448
rect 359924 410576 359976 410582
rect 359924 410518 359976 410524
rect 359832 409148 359884 409154
rect 359832 409090 359884 409096
rect 359738 396808 359794 396817
rect 359738 396743 359794 396752
rect 359648 389156 359700 389162
rect 359648 389098 359700 389104
rect 359556 379500 359608 379506
rect 359556 379442 359608 379448
rect 359752 371890 359780 396743
rect 360200 378344 360252 378350
rect 360200 378286 360252 378292
rect 359464 371884 359516 371890
rect 359464 371826 359516 371832
rect 359740 371884 359792 371890
rect 359740 371826 359792 371832
rect 359476 369170 359504 371826
rect 359648 369912 359700 369918
rect 359648 369854 359700 369860
rect 359464 369164 359516 369170
rect 359464 369106 359516 369112
rect 359200 364306 359320 364334
rect 359004 363656 359056 363662
rect 359004 363598 359056 363604
rect 359016 362982 359044 363598
rect 359004 362976 359056 362982
rect 359004 362918 359056 362924
rect 358910 353152 358966 353161
rect 358910 353087 358966 353096
rect 358820 272128 358872 272134
rect 358820 272070 358872 272076
rect 358360 271856 358412 271862
rect 358360 271798 358412 271804
rect 358924 246265 358952 353087
rect 359016 291009 359044 362918
rect 359200 362234 359228 364306
rect 359188 362228 359240 362234
rect 359188 362170 359240 362176
rect 359094 291816 359150 291825
rect 359094 291751 359150 291760
rect 359002 291000 359058 291009
rect 359002 290935 359058 290944
rect 359002 289776 359058 289785
rect 359002 289711 359058 289720
rect 359016 288833 359044 289711
rect 359002 288824 359058 288833
rect 359002 288759 359058 288768
rect 358910 246256 358966 246265
rect 358910 246191 358966 246200
rect 358818 186416 358874 186425
rect 358818 186351 358874 186360
rect 358268 166864 358320 166870
rect 358268 166806 358320 166812
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68338 358768 145522
rect 358832 79937 358860 186351
rect 358924 139369 358952 246191
rect 359016 182073 359044 288759
rect 359108 184929 359136 291751
rect 359200 287609 359228 362170
rect 359278 292768 359334 292777
rect 359278 292703 359334 292712
rect 359186 287600 359242 287609
rect 359186 287535 359242 287544
rect 359094 184920 359150 184929
rect 359094 184855 359150 184864
rect 359002 182064 359058 182073
rect 359002 181999 359058 182008
rect 358910 139360 358966 139369
rect 358910 139295 358966 139304
rect 358818 79928 358874 79937
rect 358818 79863 358874 79872
rect 359108 78305 359136 184855
rect 359200 180713 359228 287535
rect 359292 186425 359320 292703
rect 359370 291000 359426 291009
rect 359370 290935 359426 290944
rect 359278 186416 359334 186425
rect 359278 186351 359334 186360
rect 359384 183433 359412 290935
rect 359476 289785 359504 369106
rect 359556 366376 359608 366382
rect 359556 366318 359608 366324
rect 359568 292777 359596 366318
rect 359660 363730 359688 369854
rect 359648 363724 359700 363730
rect 359648 363666 359700 363672
rect 359554 292768 359610 292777
rect 359554 292703 359610 292712
rect 359660 291825 359688 363666
rect 359752 362982 359780 371826
rect 359740 362976 359792 362982
rect 359740 362918 359792 362924
rect 359646 291816 359702 291825
rect 359646 291751 359702 291760
rect 359462 289776 359518 289785
rect 359462 289711 359518 289720
rect 360212 271318 360240 378286
rect 360672 374814 360700 464442
rect 360764 377466 360792 473010
rect 360752 377460 360804 377466
rect 360752 377402 360804 377408
rect 360660 374808 360712 374814
rect 360660 374750 360712 374756
rect 360200 271312 360252 271318
rect 360200 271254 360252 271260
rect 359370 183424 359426 183433
rect 359370 183359 359426 183368
rect 359278 182064 359334 182073
rect 359278 181999 359334 182008
rect 359186 180704 359242 180713
rect 359186 180639 359242 180648
rect 359094 78296 359150 78305
rect 359094 78231 359150 78240
rect 359200 74089 359228 180639
rect 359292 75449 359320 181999
rect 359384 76945 359412 183359
rect 360212 165646 360240 271254
rect 360200 165640 360252 165646
rect 360200 165582 360252 165588
rect 359370 76936 359426 76945
rect 359370 76871 359426 76880
rect 359278 75440 359334 75449
rect 359278 75375 359334 75384
rect 359186 74080 359242 74089
rect 359186 74015 359242 74024
rect 358728 68332 358780 68338
rect 358728 68274 358780 68280
rect 358740 68202 358768 68274
rect 358728 68196 358780 68202
rect 358728 68138 358780 68144
rect 358176 59424 358228 59430
rect 358176 59366 358228 59372
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 360856 59022 360884 485182
rect 361396 481296 361448 481302
rect 361396 481238 361448 481244
rect 360936 479664 360988 479670
rect 360936 479606 360988 479612
rect 360948 165442 360976 479606
rect 361028 474224 361080 474230
rect 361028 474166 361080 474172
rect 360936 165436 360988 165442
rect 360936 165378 360988 165384
rect 361040 164218 361068 474166
rect 361304 468988 361356 468994
rect 361304 468930 361356 468936
rect 361212 468784 361264 468790
rect 361212 468726 361264 468732
rect 361120 467492 361172 467498
rect 361120 467434 361172 467440
rect 361132 271386 361160 467434
rect 361224 273154 361252 468726
rect 361316 284306 361344 468930
rect 361408 377534 361436 481238
rect 361488 474632 361540 474638
rect 361488 474574 361540 474580
rect 361500 380254 361528 474574
rect 362040 471980 362092 471986
rect 362040 471922 362092 471928
rect 362052 381546 362080 471922
rect 362132 467764 362184 467770
rect 362132 467706 362184 467712
rect 362040 381540 362092 381546
rect 362040 381482 362092 381488
rect 361488 380248 361540 380254
rect 361488 380190 361540 380196
rect 361486 378040 361542 378049
rect 361486 377975 361542 377984
rect 361396 377528 361448 377534
rect 361396 377470 361448 377476
rect 361304 284300 361356 284306
rect 361304 284242 361356 284248
rect 361212 273148 361264 273154
rect 361212 273090 361264 273096
rect 361120 271380 361172 271386
rect 361120 271322 361172 271328
rect 361028 164212 361080 164218
rect 361028 164154 361080 164160
rect 360844 59016 360896 59022
rect 360844 58958 360896 58964
rect 357624 57928 357676 57934
rect 357624 57870 357676 57876
rect 343454 57831 343456 57840
rect 313372 57802 313424 57808
rect 318260 57798 318288 57831
rect 343508 57831 343510 57840
rect 356796 57860 356848 57866
rect 343456 57802 343508 57808
rect 356796 57802 356848 57808
rect 361500 57798 361528 377975
rect 362144 377194 362172 467706
rect 362132 377188 362184 377194
rect 362132 377130 362184 377136
rect 362236 58818 362264 485386
rect 362776 484016 362828 484022
rect 362776 483958 362828 483964
rect 362316 483744 362368 483750
rect 362316 483686 362368 483692
rect 362328 70378 362356 483686
rect 362592 477352 362644 477358
rect 362592 477294 362644 477300
rect 362408 471368 362460 471374
rect 362408 471310 362460 471316
rect 362420 166938 362448 471310
rect 362500 466064 362552 466070
rect 362500 466006 362552 466012
rect 362408 166932 362460 166938
rect 362408 166874 362460 166880
rect 362512 165578 362540 466006
rect 362604 272678 362632 477294
rect 362684 474428 362736 474434
rect 362684 474370 362736 474376
rect 362592 272672 362644 272678
rect 362592 272614 362644 272620
rect 362696 271522 362724 474370
rect 362788 376718 362816 483958
rect 363880 478236 363932 478242
rect 363880 478178 363932 478184
rect 363604 475448 363656 475454
rect 363604 475390 363656 475396
rect 362868 472932 362920 472938
rect 362868 472874 362920 472880
rect 362880 377942 362908 472874
rect 363420 469192 363472 469198
rect 363420 469134 363472 469140
rect 363432 380322 363460 469134
rect 363512 468444 363564 468450
rect 363512 468386 363564 468392
rect 363420 380316 363472 380322
rect 363420 380258 363472 380264
rect 363524 378049 363552 468386
rect 363510 378040 363566 378049
rect 363510 377975 363566 377984
rect 362868 377936 362920 377942
rect 362868 377878 362920 377884
rect 362776 376712 362828 376718
rect 362776 376654 362828 376660
rect 362684 271516 362736 271522
rect 362684 271458 362736 271464
rect 362500 165572 362552 165578
rect 362500 165514 362552 165520
rect 362316 70372 362368 70378
rect 362316 70314 362368 70320
rect 362224 58812 362276 58818
rect 362224 58754 362276 58760
rect 318248 57792 318300 57798
rect 318248 57734 318300 57740
rect 361488 57792 361540 57798
rect 361488 57734 361540 57740
rect 310980 57724 311032 57730
rect 310980 57666 311032 57672
rect 305828 57656 305880 57662
rect 305828 57598 305880 57604
rect 303436 57588 303488 57594
rect 303436 57530 303488 57536
rect 363616 57458 363644 475390
rect 363788 474088 363840 474094
rect 363788 474030 363840 474036
rect 363696 474020 363748 474026
rect 363696 473962 363748 473968
rect 363708 57526 363736 473962
rect 363800 57594 363828 474030
rect 363892 164898 363920 478178
rect 363972 471300 364024 471306
rect 363972 471242 364024 471248
rect 363984 166802 364012 471242
rect 364248 470280 364300 470286
rect 364248 470222 364300 470228
rect 364064 468852 364116 468858
rect 364064 468794 364116 468800
rect 364076 272610 364104 468794
rect 364156 466268 364208 466274
rect 364156 466210 364208 466216
rect 364064 272604 364116 272610
rect 364064 272546 364116 272552
rect 364168 271590 364196 466210
rect 364260 378078 364288 470222
rect 364800 467696 364852 467702
rect 364800 467638 364852 467644
rect 364248 378072 364300 378078
rect 364248 378014 364300 378020
rect 364812 377330 364840 467638
rect 364892 464432 364944 464438
rect 364892 464374 364944 464380
rect 364800 377324 364852 377330
rect 364800 377266 364852 377272
rect 364904 374950 364932 464374
rect 364892 374944 364944 374950
rect 364892 374886 364944 374892
rect 364156 271584 364208 271590
rect 364156 271526 364208 271532
rect 363972 166796 364024 166802
rect 363972 166738 364024 166744
rect 363880 164892 363932 164898
rect 363880 164834 363932 164840
rect 364996 58750 365024 485522
rect 373264 485308 373316 485314
rect 373264 485250 373316 485256
rect 369124 485172 369176 485178
rect 369124 485114 369176 485120
rect 367008 482928 367060 482934
rect 367008 482870 367060 482876
rect 365536 482860 365588 482866
rect 365536 482802 365588 482808
rect 365352 479800 365404 479806
rect 365352 479742 365404 479748
rect 365076 476876 365128 476882
rect 365076 476818 365128 476824
rect 365088 175234 365116 476818
rect 365168 468648 365220 468654
rect 365168 468590 365220 468596
rect 365076 175228 365128 175234
rect 365076 175170 365128 175176
rect 365180 166462 365208 468590
rect 365260 467356 365312 467362
rect 365260 467298 365312 467304
rect 365272 178022 365300 467298
rect 365364 271726 365392 479742
rect 365444 477148 365496 477154
rect 365444 477090 365496 477096
rect 365456 272746 365484 477090
rect 365548 377670 365576 482802
rect 366916 482792 366968 482798
rect 366916 482734 366968 482740
rect 366640 482520 366692 482526
rect 366640 482462 366692 482468
rect 365628 480004 365680 480010
rect 365628 479946 365680 479952
rect 365536 377664 365588 377670
rect 365536 377606 365588 377612
rect 365640 376582 365668 479946
rect 366364 478168 366416 478174
rect 366364 478110 366416 478116
rect 366272 477284 366324 477290
rect 366272 477226 366324 477232
rect 366180 466336 366232 466342
rect 366180 466278 366232 466284
rect 366192 380390 366220 466278
rect 366180 380384 366232 380390
rect 366180 380326 366232 380332
rect 365628 376576 365680 376582
rect 365628 376518 365680 376524
rect 366284 376106 366312 477226
rect 366272 376100 366324 376106
rect 366272 376042 366324 376048
rect 365444 272740 365496 272746
rect 365444 272682 365496 272688
rect 365352 271720 365404 271726
rect 365352 271662 365404 271668
rect 365260 178016 365312 178022
rect 365260 177958 365312 177964
rect 365168 166456 365220 166462
rect 365168 166398 365220 166404
rect 364984 58744 365036 58750
rect 364984 58686 365036 58692
rect 366376 57866 366404 478110
rect 366456 476944 366508 476950
rect 366456 476886 366508 476892
rect 366468 164830 366496 476886
rect 366548 466132 366600 466138
rect 366548 466074 366600 466080
rect 366560 166326 366588 466074
rect 366652 271250 366680 482462
rect 366732 479868 366784 479874
rect 366732 479810 366784 479816
rect 366744 272542 366772 479810
rect 366824 467288 366876 467294
rect 366824 467230 366876 467236
rect 366836 282878 366864 467230
rect 366928 376310 366956 482734
rect 367020 380798 367048 482870
rect 368020 482588 368072 482594
rect 368020 482530 368072 482536
rect 367836 478304 367888 478310
rect 367836 478246 367888 478252
rect 367744 472728 367796 472734
rect 367744 472670 367796 472676
rect 367652 470212 367704 470218
rect 367652 470154 367704 470160
rect 367560 467560 367612 467566
rect 367560 467502 367612 467508
rect 367008 380792 367060 380798
rect 367008 380734 367060 380740
rect 367572 377874 367600 467502
rect 367560 377868 367612 377874
rect 367560 377810 367612 377816
rect 366916 376304 366968 376310
rect 366916 376246 366968 376252
rect 367664 375086 367692 470154
rect 367652 375080 367704 375086
rect 367652 375022 367704 375028
rect 366824 282872 366876 282878
rect 366824 282814 366876 282820
rect 366732 272536 366784 272542
rect 366732 272478 366784 272484
rect 366640 271244 366692 271250
rect 366640 271186 366692 271192
rect 366548 166320 366600 166326
rect 366548 166262 366600 166268
rect 366456 164824 366508 164830
rect 366456 164766 366508 164772
rect 366364 57860 366416 57866
rect 366364 57802 366416 57808
rect 363788 57588 363840 57594
rect 363788 57530 363840 57536
rect 363696 57520 363748 57526
rect 363696 57462 363748 57468
rect 298100 57452 298152 57458
rect 298100 57394 298152 57400
rect 363604 57452 363656 57458
rect 363604 57394 363656 57400
rect 367756 57390 367784 472670
rect 367848 165102 367876 478246
rect 367928 465996 367980 466002
rect 367928 465938 367980 465944
rect 367940 166530 367968 465938
rect 368032 271794 368060 482530
rect 368112 477080 368164 477086
rect 368112 477022 368164 477028
rect 368124 272814 368152 477022
rect 368388 474700 368440 474706
rect 368388 474642 368440 474648
rect 368296 474496 368348 474502
rect 368296 474438 368348 474444
rect 368204 467424 368256 467430
rect 368204 467366 368256 467372
rect 368112 272808 368164 272814
rect 368112 272750 368164 272756
rect 368020 271788 368072 271794
rect 368020 271730 368072 271736
rect 368216 271318 368244 467366
rect 368308 376446 368336 474438
rect 368400 379642 368428 474642
rect 369032 468920 369084 468926
rect 369032 468862 369084 468868
rect 369044 380458 369072 468862
rect 369032 380452 369084 380458
rect 369032 380394 369084 380400
rect 368388 379636 368440 379642
rect 368388 379578 368440 379584
rect 368388 376780 368440 376786
rect 368388 376722 368440 376728
rect 368296 376440 368348 376446
rect 368296 376382 368348 376388
rect 368204 271312 368256 271318
rect 368204 271254 368256 271260
rect 368400 252482 368428 376722
rect 368388 252476 368440 252482
rect 368388 252418 368440 252424
rect 367928 166524 367980 166530
rect 367928 166466 367980 166472
rect 367836 165096 367888 165102
rect 367836 165038 367888 165044
rect 369136 58886 369164 485114
rect 371884 485104 371936 485110
rect 371884 485046 371936 485052
rect 371700 484152 371752 484158
rect 371700 484094 371752 484100
rect 370412 483880 370464 483886
rect 370412 483822 370464 483828
rect 370320 480140 370372 480146
rect 370320 480082 370372 480088
rect 369492 479732 369544 479738
rect 369492 479674 369544 479680
rect 369216 479596 369268 479602
rect 369216 479538 369268 479544
rect 369228 165510 369256 479538
rect 369308 468580 369360 468586
rect 369308 468522 369360 468528
rect 369320 166394 369348 468522
rect 369400 465792 369452 465798
rect 369400 465734 369452 465740
rect 369308 166388 369360 166394
rect 369308 166330 369360 166336
rect 369216 165504 369268 165510
rect 369216 165446 369268 165452
rect 369412 164966 369440 465734
rect 369504 273562 369532 479674
rect 369676 474564 369728 474570
rect 369676 474506 369728 474512
rect 369584 467220 369636 467226
rect 369584 467162 369636 467168
rect 369492 273556 369544 273562
rect 369492 273498 369544 273504
rect 369596 271182 369624 467162
rect 369688 376650 369716 474506
rect 369768 473000 369820 473006
rect 369768 472942 369820 472948
rect 369676 376644 369728 376650
rect 369676 376586 369728 376592
rect 369780 375290 369808 472942
rect 370228 467628 370280 467634
rect 370228 467570 370280 467576
rect 369860 381540 369912 381546
rect 369860 381482 369912 381488
rect 369872 380934 369900 381482
rect 369860 380928 369912 380934
rect 369860 380870 369912 380876
rect 370240 376378 370268 467570
rect 370228 376372 370280 376378
rect 370228 376314 370280 376320
rect 369768 375284 369820 375290
rect 369768 375226 369820 375232
rect 370332 374882 370360 480082
rect 370424 377806 370452 483822
rect 370688 483812 370740 483818
rect 370688 483754 370740 483760
rect 370504 481092 370556 481098
rect 370504 481034 370556 481040
rect 370412 377800 370464 377806
rect 370412 377742 370464 377748
rect 370320 374876 370372 374882
rect 370320 374818 370372 374824
rect 369676 374672 369728 374678
rect 369676 374614 369728 374620
rect 369584 271176 369636 271182
rect 369584 271118 369636 271124
rect 369688 252006 369716 374614
rect 370412 273964 370464 273970
rect 370412 273906 370464 273912
rect 369768 273284 369820 273290
rect 369768 273226 369820 273232
rect 369676 252000 369728 252006
rect 369676 251942 369728 251948
rect 369400 164960 369452 164966
rect 369400 164902 369452 164908
rect 369780 145897 369808 273226
rect 370424 270026 370452 273906
rect 370412 270020 370464 270026
rect 370412 269962 370464 269968
rect 370516 165170 370544 481034
rect 370596 475516 370648 475522
rect 370596 475458 370648 475464
rect 370608 165374 370636 475458
rect 370700 271658 370728 483754
rect 370780 472864 370832 472870
rect 370780 472806 370832 472812
rect 370792 273018 370820 472806
rect 371148 471572 371200 471578
rect 371148 471514 371200 471520
rect 371056 380928 371108 380934
rect 371056 380870 371108 380876
rect 370962 379128 371018 379137
rect 370962 379063 371018 379072
rect 370870 378992 370926 379001
rect 370870 378927 370926 378936
rect 370884 273970 370912 378927
rect 370872 273964 370924 273970
rect 370872 273906 370924 273912
rect 370976 273850 371004 379063
rect 370884 273822 371004 273850
rect 370884 273254 370912 273822
rect 371068 273714 371096 380870
rect 371160 378962 371188 471514
rect 371608 464364 371660 464370
rect 371608 464306 371660 464312
rect 371620 380526 371648 464306
rect 371608 380520 371660 380526
rect 371608 380462 371660 380468
rect 371148 378956 371200 378962
rect 371148 378898 371200 378904
rect 371146 377904 371202 377913
rect 371146 377839 371202 377848
rect 370976 273686 371096 273714
rect 370976 273494 371004 273686
rect 371056 273624 371108 273630
rect 371056 273566 371108 273572
rect 370964 273488 371016 273494
rect 370964 273430 371016 273436
rect 370884 273226 371004 273254
rect 370780 273012 370832 273018
rect 370780 272954 370832 272960
rect 370688 271652 370740 271658
rect 370688 271594 370740 271600
rect 370976 270366 371004 273226
rect 370964 270360 371016 270366
rect 370964 270302 371016 270308
rect 370780 269136 370832 269142
rect 370780 269078 370832 269084
rect 370596 165368 370648 165374
rect 370596 165310 370648 165316
rect 370504 165164 370556 165170
rect 370504 165106 370556 165112
rect 370792 148510 370820 269078
rect 370780 148504 370832 148510
rect 370780 148446 370832 148452
rect 370976 148442 371004 270302
rect 370964 148436 371016 148442
rect 370964 148378 371016 148384
rect 369766 145888 369822 145897
rect 369766 145823 369822 145832
rect 371068 145761 371096 273566
rect 371054 145752 371110 145761
rect 371054 145687 371110 145696
rect 369124 58880 369176 58886
rect 369124 58822 369176 58828
rect 371160 57662 371188 377839
rect 371712 374678 371740 484094
rect 371790 380216 371846 380225
rect 371790 380151 371846 380160
rect 371700 374672 371752 374678
rect 371700 374614 371752 374620
rect 371698 273320 371754 273329
rect 371698 273255 371754 273264
rect 371712 145625 371740 273255
rect 371804 269958 371832 380151
rect 371792 269952 371844 269958
rect 371792 269894 371844 269900
rect 371698 145616 371754 145625
rect 371698 145551 371754 145560
rect 371896 59294 371924 485046
rect 372344 483948 372396 483954
rect 372344 483890 372396 483896
rect 372160 475652 372212 475658
rect 372160 475594 372212 475600
rect 371976 474156 372028 474162
rect 371976 474098 372028 474104
rect 371988 165306 372016 474098
rect 372068 465928 372120 465934
rect 372068 465870 372120 465876
rect 372080 166666 372108 465870
rect 372172 271454 372200 475594
rect 372252 472796 372304 472802
rect 372252 472738 372304 472744
rect 372264 272950 372292 472738
rect 372356 378146 372384 483890
rect 372436 471844 372488 471850
rect 372436 471786 372488 471792
rect 372448 379438 372476 471786
rect 372620 471776 372672 471782
rect 372620 471718 372672 471724
rect 372632 383654 372660 471718
rect 372632 383626 372844 383654
rect 372528 379636 372580 379642
rect 372528 379578 372580 379584
rect 372436 379432 372488 379438
rect 372436 379374 372488 379380
rect 372344 378140 372396 378146
rect 372344 378082 372396 378088
rect 372436 375352 372488 375358
rect 372436 375294 372488 375300
rect 372344 374808 372396 374814
rect 372344 374750 372396 374756
rect 372252 272944 372304 272950
rect 372252 272886 372304 272892
rect 372160 271448 372212 271454
rect 372160 271390 372212 271396
rect 372252 269816 372304 269822
rect 372252 269758 372304 269764
rect 372068 166660 372120 166666
rect 372068 166602 372120 166608
rect 371976 165300 372028 165306
rect 371976 165242 372028 165248
rect 372264 148578 372292 269758
rect 372356 251938 372384 374750
rect 372344 251932 372396 251938
rect 372344 251874 372396 251880
rect 372448 251190 372476 375294
rect 372540 270065 372568 379578
rect 372710 378856 372766 378865
rect 372620 378820 372672 378826
rect 372710 378791 372766 378800
rect 372620 378762 372672 378768
rect 372632 378418 372660 378762
rect 372724 378690 372752 378791
rect 372712 378684 372764 378690
rect 372712 378626 372764 378632
rect 372620 378412 372672 378418
rect 372620 378354 372672 378360
rect 372816 378298 372844 383626
rect 373172 378684 373224 378690
rect 373172 378626 373224 378632
rect 372632 378270 372844 378298
rect 372632 376786 372660 378270
rect 372620 376780 372672 376786
rect 372620 376722 372672 376728
rect 372632 376242 372660 376722
rect 372620 376236 372672 376242
rect 372620 376178 372672 376184
rect 372988 375420 373040 375426
rect 372988 375362 373040 375368
rect 372526 270056 372582 270065
rect 372526 269991 372582 270000
rect 373000 269249 373028 375362
rect 373080 273488 373132 273494
rect 373080 273430 373132 273436
rect 372986 269240 373042 269249
rect 372986 269175 373042 269184
rect 372528 252000 372580 252006
rect 372528 251942 372580 251948
rect 372436 251184 372488 251190
rect 372436 251126 372488 251132
rect 372252 148572 372304 148578
rect 372252 148514 372304 148520
rect 372540 148374 372568 251942
rect 373092 163538 373120 273430
rect 373184 270162 373212 378626
rect 373172 270156 373224 270162
rect 373172 270098 373224 270104
rect 373184 269142 373212 270098
rect 373172 269136 373224 269142
rect 373172 269078 373224 269084
rect 373276 167006 373304 485250
rect 378784 483676 378836 483682
rect 378784 483618 378836 483624
rect 374460 482724 374512 482730
rect 374460 482666 374512 482672
rect 373356 482452 373408 482458
rect 373356 482394 373408 482400
rect 373264 167000 373316 167006
rect 373264 166942 373316 166948
rect 373368 165238 373396 482394
rect 373908 478440 373960 478446
rect 373908 478382 373960 478388
rect 373816 477488 373868 477494
rect 373816 477430 373868 477436
rect 373724 477216 373776 477222
rect 373724 477158 373776 477164
rect 373540 474360 373592 474366
rect 373540 474302 373592 474308
rect 373448 465860 373500 465866
rect 373448 465802 373500 465808
rect 373460 166598 373488 465802
rect 373552 271017 373580 474302
rect 373632 474292 373684 474298
rect 373632 474234 373684 474240
rect 373644 273290 373672 474234
rect 373736 377738 373764 477158
rect 373828 379098 373856 477430
rect 373920 380594 373948 478382
rect 374368 475720 374420 475726
rect 374368 475662 374420 475668
rect 373908 380588 373960 380594
rect 373908 380530 373960 380536
rect 373816 379092 373868 379098
rect 373816 379034 373868 379040
rect 373908 378412 373960 378418
rect 373908 378354 373960 378360
rect 373724 377732 373776 377738
rect 373724 377674 373776 377680
rect 373816 358080 373868 358086
rect 373816 358022 373868 358028
rect 373828 273426 373856 358022
rect 373816 273420 373868 273426
rect 373816 273362 373868 273368
rect 373632 273284 373684 273290
rect 373632 273226 373684 273232
rect 373538 271008 373594 271017
rect 373538 270943 373594 270952
rect 373724 270020 373776 270026
rect 373724 269962 373776 269968
rect 373632 269952 373684 269958
rect 373632 269894 373684 269900
rect 373540 251932 373592 251938
rect 373540 251874 373592 251880
rect 373448 166592 373500 166598
rect 373448 166534 373500 166540
rect 373356 165232 373408 165238
rect 373356 165174 373408 165180
rect 373552 163606 373580 251874
rect 373540 163600 373592 163606
rect 373540 163542 373592 163548
rect 373080 163532 373132 163538
rect 373080 163474 373132 163480
rect 373264 148504 373316 148510
rect 373264 148446 373316 148452
rect 372528 148368 372580 148374
rect 372528 148310 372580 148316
rect 371884 59288 371936 59294
rect 371884 59230 371936 59236
rect 371148 57656 371200 57662
rect 371148 57598 371200 57604
rect 278320 57384 278372 57390
rect 278320 57326 278372 57332
rect 367744 57384 367796 57390
rect 367744 57326 367796 57332
rect 373276 55894 373304 148446
rect 373356 148436 373408 148442
rect 373356 148378 373408 148384
rect 373368 55962 373396 148378
rect 373644 144906 373672 269894
rect 373736 148850 373764 269962
rect 373828 148986 373856 273362
rect 373920 270094 373948 378354
rect 374380 376174 374408 475662
rect 374472 378010 374500 482666
rect 375840 482656 375892 482662
rect 375840 482598 375892 482604
rect 374736 479528 374788 479534
rect 374736 479470 374788 479476
rect 374644 472660 374696 472666
rect 374644 472602 374696 472608
rect 374552 379568 374604 379574
rect 374552 379510 374604 379516
rect 374460 378004 374512 378010
rect 374460 377946 374512 377952
rect 374564 377890 374592 379510
rect 374472 377862 374592 377890
rect 374472 377126 374500 377862
rect 374552 377256 374604 377262
rect 374552 377198 374604 377204
rect 374460 377120 374512 377126
rect 374460 377062 374512 377068
rect 374368 376168 374420 376174
rect 374368 376110 374420 376116
rect 374000 374876 374052 374882
rect 374000 374818 374052 374824
rect 374012 273222 374040 374818
rect 374000 273216 374052 273222
rect 374000 273158 374052 273164
rect 373908 270088 373960 270094
rect 373908 270030 373960 270036
rect 374460 270088 374512 270094
rect 374460 270030 374512 270036
rect 374472 269890 374500 270030
rect 374460 269884 374512 269890
rect 374460 269826 374512 269832
rect 374368 269068 374420 269074
rect 374368 269010 374420 269016
rect 374276 164144 374328 164150
rect 374276 164086 374328 164092
rect 373816 148980 373868 148986
rect 373816 148922 373868 148928
rect 373724 148844 373776 148850
rect 373724 148786 373776 148792
rect 373632 144900 373684 144906
rect 373632 144842 373684 144848
rect 373356 55956 373408 55962
rect 373356 55898 373408 55904
rect 373264 55888 373316 55894
rect 373264 55830 373316 55836
rect 277400 54460 277452 54466
rect 277400 54402 277452 54408
rect 273352 54392 273404 54398
rect 273352 54334 273404 54340
rect 373736 54330 373764 148786
rect 373828 55078 373856 148922
rect 373816 55072 373868 55078
rect 373816 55014 373868 55020
rect 374288 54398 374316 164086
rect 374380 162518 374408 269010
rect 374368 162512 374420 162518
rect 374368 162454 374420 162460
rect 374472 144838 374500 269826
rect 374564 268394 374592 377198
rect 374552 268388 374604 268394
rect 374552 268330 374604 268336
rect 374552 251184 374604 251190
rect 374552 251126 374604 251132
rect 374564 164082 374592 251126
rect 374552 164076 374604 164082
rect 374552 164018 374604 164024
rect 374460 144832 374512 144838
rect 374460 144774 374512 144780
rect 374564 56370 374592 164018
rect 374656 57322 374684 472602
rect 374748 164762 374776 479470
rect 374920 478372 374972 478378
rect 374920 478314 374972 478320
rect 374828 465724 374880 465730
rect 374828 465666 374880 465672
rect 374840 165034 374868 465666
rect 374932 270978 374960 478314
rect 375012 477012 375064 477018
rect 375012 476954 375064 476960
rect 375024 272882 375052 476954
rect 375748 476740 375800 476746
rect 375748 476682 375800 476688
rect 375196 471708 375248 471714
rect 375196 471650 375248 471656
rect 375104 471640 375156 471646
rect 375104 471582 375156 471588
rect 375116 379574 375144 471582
rect 375104 379568 375156 379574
rect 375104 379510 375156 379516
rect 375102 378720 375158 378729
rect 375102 378655 375158 378664
rect 375012 272876 375064 272882
rect 375012 272818 375064 272824
rect 374920 270972 374972 270978
rect 374920 270914 374972 270920
rect 375116 270094 375144 378655
rect 375208 378162 375236 471650
rect 375288 378752 375340 378758
rect 375286 378720 375288 378729
rect 375340 378720 375342 378729
rect 375286 378655 375342 378664
rect 375380 378344 375432 378350
rect 375380 378286 375432 378292
rect 375392 378162 375420 378286
rect 375208 378134 375420 378162
rect 375288 378072 375340 378078
rect 375288 378014 375340 378020
rect 375196 377392 375248 377398
rect 375196 377334 375248 377340
rect 375104 270088 375156 270094
rect 375104 270030 375156 270036
rect 374918 269920 374974 269929
rect 374918 269855 374974 269864
rect 374828 165028 374880 165034
rect 374828 164970 374880 164976
rect 374736 164756 374788 164762
rect 374736 164698 374788 164704
rect 374932 164150 374960 269855
rect 375116 269822 375144 270030
rect 375104 269816 375156 269822
rect 375104 269758 375156 269764
rect 375104 269680 375156 269686
rect 375104 269622 375156 269628
rect 375116 258074 375144 269622
rect 375024 258046 375144 258074
rect 374920 164144 374972 164150
rect 374920 164086 374972 164092
rect 375024 163946 375052 258046
rect 375208 252550 375236 377334
rect 375300 377262 375328 378014
rect 375288 377256 375340 377262
rect 375288 377198 375340 377204
rect 375288 377120 375340 377126
rect 375288 377062 375340 377068
rect 375300 267578 375328 377062
rect 375392 376922 375420 378134
rect 375380 376916 375432 376922
rect 375380 376858 375432 376864
rect 375760 375222 375788 476682
rect 375852 378078 375880 482598
rect 376024 482316 376076 482322
rect 376024 482258 376076 482264
rect 375840 378072 375892 378078
rect 375840 378014 375892 378020
rect 375932 377188 375984 377194
rect 375932 377130 375984 377136
rect 375748 375216 375800 375222
rect 375748 375158 375800 375164
rect 375760 373994 375788 375158
rect 375760 373966 375880 373994
rect 375746 270600 375802 270609
rect 375746 270535 375802 270544
rect 375288 267572 375340 267578
rect 375288 267514 375340 267520
rect 375196 252544 375248 252550
rect 375196 252486 375248 252492
rect 375196 251864 375248 251870
rect 375196 251806 375248 251812
rect 375208 251190 375236 251806
rect 375196 251184 375248 251190
rect 375196 251126 375248 251132
rect 375012 163940 375064 163946
rect 375012 163882 375064 163888
rect 375196 163600 375248 163606
rect 375196 163542 375248 163548
rect 375104 163532 375156 163538
rect 375104 163474 375156 163480
rect 374736 148572 374788 148578
rect 374736 148514 374788 148520
rect 374644 57316 374696 57322
rect 374644 57258 374696 57264
rect 374552 56364 374604 56370
rect 374552 56306 374604 56312
rect 374748 55146 374776 148514
rect 375012 145716 375064 145722
rect 375012 145658 375064 145664
rect 375024 144906 375052 145658
rect 374828 144900 374880 144906
rect 374828 144842 374880 144848
rect 375012 144900 375064 144906
rect 375012 144842 375064 144848
rect 374840 58614 374868 144842
rect 374828 58608 374880 58614
rect 374828 58550 374880 58556
rect 374736 55140 374788 55146
rect 374736 55082 374788 55088
rect 375116 55010 375144 163474
rect 375104 55004 375156 55010
rect 375104 54946 375156 54952
rect 375208 54942 375236 163542
rect 375300 162586 375328 267514
rect 375562 164112 375618 164121
rect 375562 164047 375618 164056
rect 375288 162580 375340 162586
rect 375288 162522 375340 162528
rect 375300 56438 375328 162522
rect 375288 56432 375340 56438
rect 375288 56374 375340 56380
rect 375196 54936 375248 54942
rect 375196 54878 375248 54884
rect 375576 54466 375604 164047
rect 375760 163878 375788 270535
rect 375852 269385 375880 373966
rect 375838 269376 375894 269385
rect 375838 269311 375894 269320
rect 375944 269074 375972 377130
rect 375932 269068 375984 269074
rect 375932 269010 375984 269016
rect 375932 252068 375984 252074
rect 375932 252010 375984 252016
rect 375944 171134 375972 252010
rect 375852 171106 375972 171134
rect 375852 165646 375880 171106
rect 375840 165640 375892 165646
rect 375840 165582 375892 165588
rect 375748 163872 375800 163878
rect 375748 163814 375800 163820
rect 375852 163690 375880 165582
rect 375668 163662 375880 163690
rect 375668 56506 375696 163662
rect 375748 162648 375800 162654
rect 375748 162590 375800 162596
rect 375760 59158 375788 162590
rect 375932 146260 375984 146266
rect 375932 146202 375984 146208
rect 375840 145852 375892 145858
rect 375840 145794 375892 145800
rect 375748 59152 375800 59158
rect 375748 59094 375800 59100
rect 375852 58478 375880 145794
rect 375840 58472 375892 58478
rect 375840 58414 375892 58420
rect 375656 56500 375708 56506
rect 375656 56442 375708 56448
rect 375944 56098 375972 146202
rect 376036 68105 376064 482258
rect 377496 481160 377548 481166
rect 377496 481102 377548 481108
rect 376116 481024 376168 481030
rect 376116 480966 376168 480972
rect 376128 164665 376156 480966
rect 376300 476808 376352 476814
rect 376300 476750 376352 476756
rect 376208 468512 376260 468518
rect 376208 468454 376260 468460
rect 376220 271046 376248 468454
rect 376208 271040 376260 271046
rect 376208 270982 376260 270988
rect 376208 252476 376260 252482
rect 376208 252418 376260 252424
rect 376220 252074 376248 252418
rect 376208 252068 376260 252074
rect 376208 252010 376260 252016
rect 376312 165617 376340 476750
rect 376760 475788 376812 475794
rect 376760 475730 376812 475736
rect 376484 471436 376536 471442
rect 376484 471378 376536 471384
rect 376392 466200 376444 466206
rect 376392 466142 376444 466148
rect 376404 271561 376432 466142
rect 376496 379846 376524 471378
rect 376576 469940 376628 469946
rect 376576 469882 376628 469888
rect 376484 379840 376536 379846
rect 376484 379782 376536 379788
rect 376496 377058 376524 379782
rect 376588 378894 376616 469882
rect 376576 378888 376628 378894
rect 376576 378830 376628 378836
rect 376484 377052 376536 377058
rect 376484 376994 376536 377000
rect 376484 376916 376536 376922
rect 376484 376858 376536 376864
rect 376390 271552 376446 271561
rect 376390 271487 376446 271496
rect 376496 270337 376524 376858
rect 376588 271289 376616 378830
rect 376668 377460 376720 377466
rect 376668 377402 376720 377408
rect 376680 377194 376708 377402
rect 376668 377188 376720 377194
rect 376668 377130 376720 377136
rect 376668 377052 376720 377058
rect 376668 376994 376720 377000
rect 376574 271280 376630 271289
rect 376574 271215 376630 271224
rect 376588 270609 376616 271215
rect 376574 270600 376630 270609
rect 376574 270535 376630 270544
rect 376482 270328 376538 270337
rect 376482 270263 376538 270272
rect 376390 270056 376446 270065
rect 376390 269991 376446 270000
rect 376298 165608 376354 165617
rect 376298 165543 376354 165552
rect 376404 164914 376432 269991
rect 376496 269929 376524 270263
rect 376680 270230 376708 376994
rect 376772 375426 376800 475730
rect 377404 470076 377456 470082
rect 377404 470018 377456 470024
rect 377312 468716 377364 468722
rect 377312 468658 377364 468664
rect 377220 417444 377272 417450
rect 377220 417386 377272 417392
rect 377232 416945 377260 417386
rect 377218 416936 377274 416945
rect 377218 416871 377274 416880
rect 376942 415304 376998 415313
rect 376942 415239 376998 415248
rect 376956 414769 376984 415239
rect 376942 414760 376998 414769
rect 376942 414695 376998 414704
rect 376956 402974 376984 414695
rect 377218 412040 377274 412049
rect 377218 411975 377274 411984
rect 377232 411942 377260 411975
rect 377220 411936 377272 411942
rect 377220 411878 377272 411884
rect 377218 410952 377274 410961
rect 377218 410887 377274 410896
rect 377232 410582 377260 410887
rect 377220 410576 377272 410582
rect 377220 410518 377272 410524
rect 376956 402946 377076 402974
rect 376944 391944 376996 391950
rect 376944 391886 376996 391892
rect 376956 390969 376984 391886
rect 376942 390960 376998 390969
rect 376942 390895 376998 390904
rect 376944 390516 376996 390522
rect 376944 390458 376996 390464
rect 376956 389337 376984 390458
rect 376942 389328 376998 389337
rect 376942 389263 376998 389272
rect 376944 389156 376996 389162
rect 376944 389098 376996 389104
rect 376956 389065 376984 389098
rect 376942 389056 376998 389065
rect 376942 388991 376998 389000
rect 376760 375420 376812 375426
rect 376760 375362 376812 375368
rect 376760 375284 376812 375290
rect 376760 375226 376812 375232
rect 376772 374921 376800 375226
rect 376758 374912 376814 374921
rect 376758 374847 376814 374856
rect 377048 373994 377076 402946
rect 377324 380662 377352 468658
rect 377416 415313 377444 470018
rect 377402 415304 377458 415313
rect 377402 415239 377458 415248
rect 377402 409184 377458 409193
rect 377402 409119 377404 409128
rect 377456 409119 377458 409128
rect 377404 409090 377456 409096
rect 377312 380656 377364 380662
rect 377312 380598 377364 380604
rect 377404 379432 377456 379438
rect 377404 379374 377456 379380
rect 377416 378826 377444 379374
rect 377404 378820 377456 378826
rect 377404 378762 377456 378768
rect 377416 378185 377444 378762
rect 377402 378176 377458 378185
rect 377402 378111 377458 378120
rect 377508 376038 377536 481102
rect 377680 470144 377732 470150
rect 377680 470086 377732 470092
rect 377588 470008 377640 470014
rect 377588 469950 377640 469956
rect 377600 413953 377628 469950
rect 377692 422294 377720 470086
rect 377692 422266 377812 422294
rect 377784 417897 377812 422266
rect 377770 417888 377826 417897
rect 377770 417823 377826 417832
rect 377586 413944 377642 413953
rect 377586 413879 377642 413888
rect 377586 412040 377642 412049
rect 377586 411975 377642 411984
rect 377496 376032 377548 376038
rect 377496 375974 377548 375980
rect 377404 375420 377456 375426
rect 377404 375362 377456 375368
rect 377416 375154 377444 375362
rect 377404 375148 377456 375154
rect 377404 375090 377456 375096
rect 377496 375080 377548 375086
rect 377496 375022 377548 375028
rect 377128 375012 377180 375018
rect 377128 374954 377180 374960
rect 376956 373966 377076 373994
rect 376956 316034 376984 373966
rect 377036 358624 377088 358630
rect 377036 358566 377088 358572
rect 376864 316006 376984 316034
rect 376864 307873 376892 316006
rect 376850 307864 376906 307873
rect 376850 307799 376906 307808
rect 376864 287054 376892 307799
rect 376942 307728 376998 307737
rect 376942 307663 376998 307672
rect 376772 287026 376892 287054
rect 376772 277394 376800 287026
rect 376852 284300 376904 284306
rect 376852 284242 376904 284248
rect 376864 284073 376892 284242
rect 376850 284064 376906 284073
rect 376850 283999 376906 284008
rect 376956 282418 376984 307663
rect 376864 282390 376984 282418
rect 376864 282076 376892 282390
rect 376942 282296 376998 282305
rect 376942 282231 376998 282240
rect 376956 282198 376984 282231
rect 376944 282192 376996 282198
rect 376944 282134 376996 282140
rect 376864 282048 376984 282076
rect 376772 277366 376892 277394
rect 376668 270224 376720 270230
rect 376668 270166 376720 270172
rect 376482 269920 376538 269929
rect 376482 269855 376538 269864
rect 376484 269748 376536 269754
rect 376484 269690 376536 269696
rect 376220 164886 376432 164914
rect 376114 164656 376170 164665
rect 376114 164591 376170 164600
rect 376220 162722 376248 164886
rect 376496 162858 376524 269690
rect 376576 268388 376628 268394
rect 376576 268330 376628 268336
rect 376484 162852 376536 162858
rect 376484 162794 376536 162800
rect 376208 162716 376260 162722
rect 376208 162658 376260 162664
rect 376116 145648 376168 145654
rect 376116 145590 376168 145596
rect 376128 144838 376156 145590
rect 376116 144832 376168 144838
rect 376116 144774 376168 144780
rect 376022 68096 376078 68105
rect 376022 68031 376078 68040
rect 375932 56092 375984 56098
rect 375932 56034 375984 56040
rect 376128 54602 376156 144774
rect 376220 59226 376248 162658
rect 376300 161900 376352 161906
rect 376300 161842 376352 161848
rect 376208 59220 376260 59226
rect 376208 59162 376260 59168
rect 376312 59090 376340 161842
rect 376588 145858 376616 268330
rect 376680 145858 376708 270166
rect 376758 269376 376814 269385
rect 376758 269311 376814 269320
rect 376772 162790 376800 269311
rect 376864 201385 376892 277366
rect 376850 201376 376906 201385
rect 376850 201311 376906 201320
rect 376956 199889 376984 282048
rect 377048 270434 377076 358566
rect 377036 270428 377088 270434
rect 377036 270370 377088 270376
rect 377140 269754 377168 374954
rect 377402 310856 377458 310865
rect 377402 310791 377458 310800
rect 377218 310040 377274 310049
rect 377218 309975 377274 309984
rect 377128 269748 377180 269754
rect 377128 269690 377180 269696
rect 377232 209774 377260 309975
rect 377310 302152 377366 302161
rect 377310 302087 377366 302096
rect 377048 209746 377260 209774
rect 377048 203017 377076 209746
rect 377218 203960 377274 203969
rect 377218 203895 377274 203904
rect 377034 203008 377090 203017
rect 377034 202943 377090 202952
rect 376942 199880 376998 199889
rect 376942 199815 376998 199824
rect 376956 180794 376984 199815
rect 376864 180766 376984 180794
rect 376864 171134 376892 180766
rect 376944 178016 376996 178022
rect 376944 177958 376996 177964
rect 376956 177041 376984 177958
rect 376942 177032 376998 177041
rect 376942 176967 376998 176976
rect 376944 175976 376996 175982
rect 376944 175918 376996 175924
rect 376956 175409 376984 175918
rect 376942 175400 376998 175409
rect 376942 175335 376998 175344
rect 376944 175228 376996 175234
rect 376944 175170 376996 175176
rect 376956 175137 376984 175170
rect 376942 175128 376998 175137
rect 376942 175063 376998 175072
rect 376864 171106 376984 171134
rect 376760 162784 376812 162790
rect 376760 162726 376812 162732
rect 376772 161906 376800 162726
rect 376760 161900 376812 161906
rect 376760 161842 376812 161848
rect 376576 145852 376628 145858
rect 376576 145794 376628 145800
rect 376668 145852 376720 145858
rect 376668 145794 376720 145800
rect 376680 142154 376708 145794
rect 376496 142126 376708 142154
rect 376300 59084 376352 59090
rect 376300 59026 376352 59032
rect 376116 54596 376168 54602
rect 376116 54538 376168 54544
rect 376496 54534 376524 142126
rect 376956 92857 376984 171106
rect 377048 95985 377076 202943
rect 377232 96937 377260 203895
rect 377324 195265 377352 302087
rect 377416 203969 377444 310791
rect 377508 268870 377536 375022
rect 377600 305017 377628 411975
rect 377680 410576 377732 410582
rect 377680 410518 377732 410524
rect 377692 306374 377720 410518
rect 377784 310865 377812 417823
rect 377954 416936 378010 416945
rect 377954 416871 378010 416880
rect 377862 413944 377918 413953
rect 377862 413879 377918 413888
rect 377770 310856 377826 310865
rect 377770 310791 377826 310800
rect 377876 307737 377904 413879
rect 377968 310049 377996 416871
rect 378046 409184 378102 409193
rect 378046 409119 378102 409128
rect 377954 310040 378010 310049
rect 377954 309975 378010 309984
rect 377862 307728 377918 307737
rect 377862 307663 377918 307672
rect 377876 306921 377904 307663
rect 377862 306912 377918 306921
rect 377862 306847 377918 306856
rect 377692 306346 377904 306374
rect 377586 305008 377642 305017
rect 377586 304943 377642 304952
rect 377600 296714 377628 304943
rect 377876 303929 377904 306346
rect 377862 303920 377918 303929
rect 377862 303855 377918 303864
rect 377600 296686 377812 296714
rect 377588 282872 377640 282878
rect 377588 282814 377640 282820
rect 377600 282169 377628 282814
rect 377586 282160 377642 282169
rect 377586 282095 377642 282104
rect 377496 268864 377548 268870
rect 377496 268806 377548 268812
rect 377680 267708 377732 267714
rect 377680 267650 377732 267656
rect 377692 267617 377720 267650
rect 377678 267608 377734 267617
rect 377678 267543 377734 267552
rect 377680 252544 377732 252550
rect 377678 252512 377680 252521
rect 377732 252512 377734 252521
rect 377678 252447 377734 252456
rect 377402 203960 377458 203969
rect 377402 203895 377458 203904
rect 377586 201376 377642 201385
rect 377586 201311 377642 201320
rect 377600 200841 377628 201311
rect 377586 200832 377642 200841
rect 377586 200767 377642 200776
rect 377310 195256 377366 195265
rect 377310 195191 377366 195200
rect 377312 145988 377364 145994
rect 377312 145930 377364 145936
rect 377218 96928 377274 96937
rect 377218 96863 377274 96872
rect 377034 95976 377090 95985
rect 377034 95911 377090 95920
rect 376942 92848 376998 92857
rect 376942 92783 376998 92792
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376666 68912 376722 68921
rect 376666 68847 376722 68856
rect 376680 57934 376708 68847
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 376668 57928 376720 57934
rect 376668 57870 376720 57876
rect 377324 54670 377352 145930
rect 377494 145752 377550 145761
rect 377494 145687 377550 145696
rect 377508 59498 377536 145687
rect 377600 93809 377628 200767
rect 377784 200114 377812 296686
rect 377692 200086 377812 200114
rect 377692 198121 377720 200086
rect 377678 198112 377734 198121
rect 377678 198047 377734 198056
rect 377586 93800 377642 93809
rect 377586 93735 377642 93744
rect 377692 91089 377720 198047
rect 377876 197033 377904 303855
rect 378060 302161 378088 409119
rect 378140 374944 378192 374950
rect 378140 374886 378192 374892
rect 378152 374678 378180 374886
rect 378140 374672 378192 374678
rect 378140 374614 378192 374620
rect 378046 302152 378102 302161
rect 378046 302087 378102 302096
rect 378152 273630 378180 374614
rect 378692 357876 378744 357882
rect 378692 357818 378744 357824
rect 378704 273630 378732 357818
rect 378140 273624 378192 273630
rect 378140 273566 378192 273572
rect 378692 273624 378744 273630
rect 378692 273566 378744 273572
rect 378152 272474 378180 273566
rect 378506 273320 378562 273329
rect 378506 273255 378562 273264
rect 378140 272468 378192 272474
rect 378140 272410 378192 272416
rect 378048 270428 378100 270434
rect 378048 270370 378100 270376
rect 377956 268864 378008 268870
rect 377956 268806 378008 268812
rect 377862 197024 377918 197033
rect 377862 196959 377918 196968
rect 377770 195256 377826 195265
rect 377770 195191 377826 195200
rect 377678 91080 377734 91089
rect 377678 91015 377734 91024
rect 377784 88233 377812 195191
rect 377876 90001 377904 196959
rect 377968 146266 377996 268806
rect 377956 146260 378008 146266
rect 377956 146202 378008 146208
rect 377968 145926 377996 146202
rect 377956 145920 378008 145926
rect 377956 145862 378008 145868
rect 378060 145314 378088 270370
rect 378416 269612 378468 269618
rect 378416 269554 378468 269560
rect 378428 146198 378456 269554
rect 378416 146192 378468 146198
rect 378416 146134 378468 146140
rect 378048 145308 378100 145314
rect 378048 145250 378100 145256
rect 377862 89992 377918 90001
rect 377862 89927 377918 89936
rect 377770 88224 377826 88233
rect 377770 88159 377826 88168
rect 377496 59492 377548 59498
rect 377496 59434 377548 59440
rect 378060 54738 378088 145250
rect 378520 57730 378548 273255
rect 378600 269544 378652 269550
rect 378600 269486 378652 269492
rect 378612 146266 378640 269486
rect 378690 269240 378746 269249
rect 378690 269175 378746 269184
rect 378704 162654 378732 269175
rect 378796 165345 378824 483618
rect 378968 482384 379020 482390
rect 378968 482326 379020 482332
rect 378876 475380 378928 475386
rect 378876 475322 378928 475328
rect 378782 165336 378838 165345
rect 378782 165271 378838 165280
rect 378888 164694 378916 475322
rect 378980 165481 379008 482326
rect 434824 480962 434852 592311
rect 434916 539345 434944 647838
rect 436100 643136 436152 643142
rect 436100 643078 436152 643084
rect 436112 620945 436140 643078
rect 457444 641776 457496 641782
rect 457444 641718 457496 641724
rect 436192 641232 436244 641238
rect 436192 641174 436244 641180
rect 436204 630465 436232 641174
rect 436190 630456 436246 630465
rect 436190 630391 436246 630400
rect 436098 620936 436154 620945
rect 436098 620871 436154 620880
rect 457456 597553 457484 641718
rect 494072 641102 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 494060 641096 494112 641102
rect 494060 641038 494112 641044
rect 457628 640960 457680 640966
rect 457628 640902 457680 640908
rect 457536 639192 457588 639198
rect 457536 639134 457588 639140
rect 457548 616865 457576 639134
rect 457640 623121 457668 640902
rect 457720 640892 457772 640898
rect 457720 640834 457772 640840
rect 457732 629241 457760 640834
rect 457812 640824 457864 640830
rect 457812 640766 457864 640772
rect 457824 634817 457852 640766
rect 471612 640756 471664 640762
rect 471612 640698 471664 640704
rect 471624 634984 471652 640698
rect 483204 640620 483256 640626
rect 483204 640562 483256 640568
rect 483216 634984 483244 640562
rect 494796 640552 494848 640558
rect 494796 640494 494848 640500
rect 494808 634984 494836 640494
rect 501236 640484 501288 640490
rect 501236 640426 501288 640432
rect 501248 634984 501276 640426
rect 512000 640416 512052 640422
rect 512000 640358 512052 640364
rect 477130 634944 477186 634953
rect 465198 634914 465488 634930
rect 465198 634908 465500 634914
rect 465198 634902 465448 634908
rect 488722 634944 488778 634953
rect 477186 634902 477434 634930
rect 477130 634879 477186 634888
rect 506754 634944 506810 634953
rect 488778 634902 489026 634930
rect 488722 634879 488778 634888
rect 506810 634902 507058 634930
rect 506754 634879 506810 634888
rect 465448 634850 465500 634856
rect 457810 634808 457866 634817
rect 457810 634743 457866 634752
rect 457718 629232 457774 629241
rect 457718 629167 457774 629176
rect 457626 623112 457682 623121
rect 457626 623047 457682 623056
rect 512012 619585 512040 640358
rect 512184 640348 512236 640354
rect 512184 640290 512236 640296
rect 512092 639056 512144 639062
rect 512092 638998 512144 639004
rect 512104 626521 512132 638998
rect 512196 631961 512224 640290
rect 580356 639260 580408 639266
rect 580356 639202 580408 639208
rect 580264 634840 580316 634846
rect 580264 634782 580316 634788
rect 512182 631952 512238 631961
rect 512182 631887 512238 631896
rect 512090 626512 512146 626521
rect 512090 626447 512146 626456
rect 511998 619576 512054 619585
rect 511998 619511 512054 619520
rect 457534 616856 457590 616865
rect 457534 616791 457590 616800
rect 511998 612776 512054 612785
rect 511998 612711 512054 612720
rect 457626 608968 457682 608977
rect 457626 608903 457682 608912
rect 457534 603120 457590 603129
rect 457534 603055 457590 603064
rect 457442 597544 457498 597553
rect 457442 597479 457498 597488
rect 436098 597136 436154 597145
rect 436098 597071 436154 597080
rect 434902 539336 434958 539345
rect 434902 539271 434958 539280
rect 436112 529718 436140 597071
rect 457442 590744 457498 590753
rect 457442 590679 457498 590688
rect 436190 582176 436246 582185
rect 436190 582111 436246 582120
rect 436204 529786 436232 582111
rect 436282 577416 436338 577425
rect 436282 577351 436338 577360
rect 436192 529780 436244 529786
rect 436192 529722 436244 529728
rect 436100 529712 436152 529718
rect 436100 529654 436152 529660
rect 436296 529514 436324 577351
rect 436374 572656 436430 572665
rect 436374 572591 436430 572600
rect 436388 529582 436416 572591
rect 436466 563136 436522 563145
rect 436466 563071 436522 563080
rect 436480 529854 436508 563071
rect 436558 558376 436614 558385
rect 436558 558311 436614 558320
rect 436468 529848 436520 529854
rect 436468 529790 436520 529796
rect 436572 529650 436600 558311
rect 436650 553616 436706 553625
rect 436650 553551 436706 553560
rect 436560 529644 436612 529650
rect 436560 529586 436612 529592
rect 436376 529576 436428 529582
rect 436376 529518 436428 529524
rect 436284 529508 436336 529514
rect 436284 529450 436336 529456
rect 436664 528086 436692 553551
rect 436742 548856 436798 548865
rect 436742 548791 436798 548800
rect 436652 528080 436704 528086
rect 436652 528022 436704 528028
rect 436756 528018 436784 548791
rect 436834 544096 436890 544105
rect 436834 544031 436890 544040
rect 436848 528154 436876 544031
rect 436926 534576 436982 534585
rect 436926 534511 436982 534520
rect 436940 528222 436968 534511
rect 457456 529922 457484 590679
rect 457444 529916 457496 529922
rect 457444 529858 457496 529864
rect 436928 528216 436980 528222
rect 436928 528158 436980 528164
rect 436836 528148 436888 528154
rect 436836 528090 436888 528096
rect 436744 528012 436796 528018
rect 436744 527954 436796 527960
rect 457548 486577 457576 603055
rect 457640 524414 457668 608903
rect 459572 585126 460046 585154
rect 465092 585126 465842 585154
rect 470612 585126 471638 585154
rect 476132 585126 477434 585154
rect 483032 585126 483230 585154
rect 488552 585126 489670 585154
rect 495466 585126 495572 585154
rect 459572 528290 459600 585126
rect 465092 528358 465120 585126
rect 465080 528352 465132 528358
rect 465080 528294 465132 528300
rect 459560 528284 459612 528290
rect 459560 528226 459612 528232
rect 470612 525638 470640 585126
rect 476132 525706 476160 585126
rect 476120 525700 476172 525706
rect 476120 525642 476172 525648
rect 470600 525632 470652 525638
rect 470600 525574 470652 525580
rect 457628 524408 457680 524414
rect 457628 524350 457680 524356
rect 457534 486568 457590 486577
rect 457534 486503 457590 486512
rect 434812 480956 434864 480962
rect 434812 480898 434864 480904
rect 379244 480072 379296 480078
rect 379244 480014 379296 480020
rect 379060 475584 379112 475590
rect 379060 475526 379112 475532
rect 379072 271114 379100 475526
rect 379152 467152 379204 467158
rect 379152 467094 379204 467100
rect 379164 271833 379192 467094
rect 379256 377482 379284 480014
rect 379336 477420 379388 477426
rect 379336 477362 379388 477368
rect 379348 378622 379376 477362
rect 483032 475425 483060 585126
rect 488552 528426 488580 585126
rect 495544 567194 495572 585126
rect 495452 567166 495572 567194
rect 500972 585126 501262 585154
rect 506492 585126 507058 585154
rect 495452 528494 495480 567166
rect 500972 529553 501000 585126
rect 500958 529544 501014 529553
rect 500958 529479 501014 529488
rect 495440 528488 495492 528494
rect 495440 528430 495492 528436
rect 488540 528420 488592 528426
rect 488540 528362 488592 528368
rect 506492 518129 506520 585126
rect 506478 518120 506534 518129
rect 506478 518055 506534 518064
rect 512012 487801 512040 612711
rect 512182 606384 512238 606393
rect 512182 606319 512238 606328
rect 512090 600400 512146 600409
rect 512090 600335 512146 600344
rect 511998 487792 512054 487801
rect 511998 487727 512054 487736
rect 512104 479505 512132 600335
rect 512196 528562 512224 606319
rect 512274 594008 512330 594017
rect 512274 593943 512330 593952
rect 512184 528556 512236 528562
rect 512184 528498 512236 528504
rect 512288 525774 512316 593943
rect 513288 586560 513340 586566
rect 513286 586528 513288 586537
rect 560944 586560 560996 586566
rect 513340 586528 513342 586537
rect 560944 586502 560996 586508
rect 513286 586463 513342 586472
rect 512276 525768 512328 525774
rect 512276 525710 512328 525716
rect 519544 524476 519596 524482
rect 519544 524418 519596 524424
rect 512090 479496 512146 479505
rect 512090 479431 512146 479440
rect 483018 475416 483074 475425
rect 483018 475351 483074 475360
rect 379980 469872 380032 469878
rect 379980 469814 380032 469820
rect 379702 382392 379758 382401
rect 379702 382327 379758 382336
rect 379520 378956 379572 378962
rect 379520 378898 379572 378904
rect 379336 378616 379388 378622
rect 379336 378558 379388 378564
rect 379532 378486 379560 378898
rect 379520 378480 379572 378486
rect 379520 378422 379572 378428
rect 379256 377454 379468 377482
rect 379336 377324 379388 377330
rect 379336 377266 379388 377272
rect 379244 358148 379296 358154
rect 379244 358090 379296 358096
rect 379150 271824 379206 271833
rect 379150 271759 379206 271768
rect 379060 271108 379112 271114
rect 379060 271050 379112 271056
rect 379256 270298 379284 358090
rect 379244 270292 379296 270298
rect 379244 270234 379296 270240
rect 379348 268802 379376 377266
rect 379440 374678 379468 377454
rect 379532 377074 379560 378422
rect 379532 377046 379652 377074
rect 379428 374672 379480 374678
rect 379428 374614 379480 374620
rect 379440 373994 379468 374614
rect 379440 373966 379560 373994
rect 379428 358012 379480 358018
rect 379428 357954 379480 357960
rect 379440 270473 379468 357954
rect 379532 357377 379560 373966
rect 379518 357368 379574 357377
rect 379518 357303 379574 357312
rect 379426 270464 379482 270473
rect 379426 270399 379482 270408
rect 379440 270298 379560 270314
rect 379428 270292 379560 270298
rect 379480 270286 379560 270292
rect 379428 270234 379480 270240
rect 379532 269822 379560 270286
rect 379520 269816 379572 269822
rect 379520 269758 379572 269764
rect 379152 268796 379204 268802
rect 379152 268738 379204 268744
rect 379336 268796 379388 268802
rect 379336 268738 379388 268744
rect 379060 266416 379112 266422
rect 379060 266358 379112 266364
rect 378966 165472 379022 165481
rect 378966 165407 379022 165416
rect 378876 164688 378928 164694
rect 378876 164630 378928 164636
rect 378692 162648 378744 162654
rect 378692 162590 378744 162596
rect 378968 162512 379020 162518
rect 378968 162454 379020 162460
rect 378980 161498 379008 162454
rect 378968 161492 379020 161498
rect 378968 161434 379020 161440
rect 378874 146296 378930 146305
rect 378600 146260 378652 146266
rect 378874 146231 378930 146240
rect 378600 146202 378652 146208
rect 378888 146033 378916 146231
rect 378874 146024 378930 146033
rect 378874 145959 378930 145968
rect 378692 145444 378744 145450
rect 378692 145386 378744 145392
rect 378704 59634 378732 145386
rect 378784 145376 378836 145382
rect 378784 145318 378836 145324
rect 378796 59702 378824 145318
rect 378784 59696 378836 59702
rect 378784 59638 378836 59644
rect 378692 59628 378744 59634
rect 378692 59570 378744 59576
rect 378508 57724 378560 57730
rect 378508 57666 378560 57672
rect 378888 57254 378916 145959
rect 378980 59566 379008 161434
rect 379072 149054 379100 266358
rect 379060 149048 379112 149054
rect 379060 148990 379112 148996
rect 379072 147801 379100 148990
rect 379058 147792 379114 147801
rect 379058 147727 379114 147736
rect 379060 146124 379112 146130
rect 379060 146066 379112 146072
rect 378968 59560 379020 59566
rect 378968 59502 379020 59508
rect 378876 57248 378928 57254
rect 378876 57190 378928 57196
rect 379072 56166 379100 146066
rect 379164 145994 379192 268738
rect 379336 147688 379388 147694
rect 379336 147630 379388 147636
rect 379244 146260 379296 146266
rect 379244 146202 379296 146208
rect 379152 145988 379204 145994
rect 379152 145930 379204 145936
rect 379256 145518 379284 146202
rect 379244 145512 379296 145518
rect 379244 145454 379296 145460
rect 379060 56160 379112 56166
rect 379060 56102 379112 56108
rect 379256 55214 379284 145454
rect 379348 56302 379376 147630
rect 379428 146192 379480 146198
rect 379428 146134 379480 146140
rect 379440 146062 379468 146134
rect 379532 146130 379560 269758
rect 379624 269618 379652 377046
rect 379716 375358 379744 382327
rect 379992 379030 380020 469814
rect 498476 466608 498528 466614
rect 498474 466576 498476 466585
rect 517796 466608 517848 466614
rect 498528 466576 498530 466585
rect 498474 466511 498530 466520
rect 499762 466576 499818 466585
rect 499762 466511 499764 466520
rect 499816 466511 499818 466520
rect 510894 466576 510950 466585
rect 517796 466550 517848 466556
rect 510894 466511 510896 466520
rect 499764 466482 499816 466488
rect 510948 466511 510950 466520
rect 517520 466540 517572 466546
rect 510896 466482 510948 466488
rect 517520 466482 517572 466488
rect 431132 380928 431184 380934
rect 431130 380896 431132 380905
rect 431184 380896 431186 380905
rect 431130 380831 431186 380840
rect 433614 380896 433670 380905
rect 433614 380831 433670 380840
rect 438490 380896 438546 380905
rect 438490 380831 438546 380840
rect 380992 380792 381044 380798
rect 380992 380734 381044 380740
rect 410706 380760 410762 380769
rect 380900 380724 380952 380730
rect 380900 380666 380952 380672
rect 380912 379710 380940 380666
rect 381004 379778 381032 380734
rect 410706 380695 410762 380704
rect 421102 380760 421158 380769
rect 421102 380695 421158 380704
rect 410720 380662 410748 380695
rect 410708 380656 410760 380662
rect 405462 380624 405518 380633
rect 410708 380598 410760 380604
rect 413466 380624 413522 380633
rect 405462 380559 405518 380568
rect 413466 380559 413522 380568
rect 419446 380624 419502 380633
rect 421116 380594 421144 380695
rect 419446 380559 419502 380568
rect 421104 380588 421156 380594
rect 405476 379846 405504 380559
rect 405464 379840 405516 379846
rect 405464 379782 405516 379788
rect 413480 379778 413508 380559
rect 380992 379772 381044 379778
rect 380992 379714 381044 379720
rect 381360 379772 381412 379778
rect 381360 379714 381412 379720
rect 413468 379772 413520 379778
rect 413468 379714 413520 379720
rect 380900 379704 380952 379710
rect 380900 379646 380952 379652
rect 380912 379250 380940 379646
rect 380912 379222 381032 379250
rect 380900 379092 380952 379098
rect 380900 379034 380952 379040
rect 379796 379024 379848 379030
rect 379796 378966 379848 378972
rect 379980 379024 380032 379030
rect 379980 378966 380032 378972
rect 379704 375352 379756 375358
rect 379704 375294 379756 375300
rect 379704 273624 379756 273630
rect 379704 273566 379756 273572
rect 379612 269612 379664 269618
rect 379612 269554 379664 269560
rect 379716 164014 379744 273566
rect 379808 271153 379836 378966
rect 379888 378616 379940 378622
rect 379888 378558 379940 378564
rect 379794 271144 379850 271153
rect 379794 271079 379850 271088
rect 379794 270464 379850 270473
rect 379794 270399 379850 270408
rect 379808 269793 379836 270399
rect 379900 270230 379928 378558
rect 380912 378554 380940 379034
rect 380900 378548 380952 378554
rect 380900 378490 380952 378496
rect 381004 378162 381032 379222
rect 381266 378856 381322 378865
rect 381266 378791 381322 378800
rect 381082 378720 381138 378729
rect 381082 378655 381138 378664
rect 380912 378134 381032 378162
rect 379980 375964 380032 375970
rect 379980 375906 380032 375912
rect 379888 270224 379940 270230
rect 379888 270166 379940 270172
rect 379794 269784 379850 269793
rect 379794 269719 379850 269728
rect 379704 164008 379756 164014
rect 379704 163950 379756 163956
rect 379612 162852 379664 162858
rect 379612 162794 379664 162800
rect 379624 162178 379652 162794
rect 379612 162172 379664 162178
rect 379612 162114 379664 162120
rect 379520 146124 379572 146130
rect 379520 146066 379572 146072
rect 379428 146056 379480 146062
rect 379428 145998 379480 146004
rect 379336 56296 379388 56302
rect 379336 56238 379388 56244
rect 379440 56030 379468 145998
rect 379624 59362 379652 162114
rect 379612 59356 379664 59362
rect 379612 59298 379664 59304
rect 379428 56024 379480 56030
rect 379428 55966 379480 55972
rect 379244 55208 379296 55214
rect 379244 55150 379296 55156
rect 379716 54806 379744 163950
rect 379808 148918 379836 269719
rect 379900 269550 379928 270166
rect 379888 269544 379940 269550
rect 379888 269486 379940 269492
rect 379992 269006 380020 375906
rect 380912 357882 380940 378134
rect 380992 377188 381044 377194
rect 380992 377130 381044 377136
rect 381004 358154 381032 377130
rect 380992 358148 381044 358154
rect 380992 358090 381044 358096
rect 381096 358086 381124 378655
rect 381176 378548 381228 378554
rect 381176 378490 381228 378496
rect 381188 358630 381216 378490
rect 381176 358624 381228 358630
rect 381176 358566 381228 358572
rect 381084 358080 381136 358086
rect 381084 358022 381136 358028
rect 381280 358018 381308 378791
rect 381372 377194 381400 379714
rect 419460 379642 419488 380559
rect 421104 380530 421156 380536
rect 433628 380526 433656 380831
rect 436006 380760 436062 380769
rect 436006 380695 436062 380704
rect 434350 380624 434406 380633
rect 434350 380559 434406 380568
rect 433616 380520 433668 380526
rect 426438 380488 426494 380497
rect 433616 380462 433668 380468
rect 426438 380423 426494 380432
rect 426452 379710 426480 380423
rect 426440 379704 426492 379710
rect 426440 379646 426492 379652
rect 419448 379636 419500 379642
rect 419448 379578 419500 379584
rect 434364 379574 434392 380559
rect 436020 380458 436048 380695
rect 436008 380452 436060 380458
rect 436008 380394 436060 380400
rect 438504 380390 438532 380831
rect 440882 380760 440938 380769
rect 440882 380695 440938 380704
rect 443458 380760 443514 380769
rect 443458 380695 443514 380704
rect 438492 380384 438544 380390
rect 438492 380326 438544 380332
rect 440896 380322 440924 380695
rect 440884 380316 440936 380322
rect 440884 380258 440936 380264
rect 443472 380254 443500 380695
rect 485962 380624 486018 380633
rect 485962 380559 486018 380568
rect 443460 380248 443512 380254
rect 443460 380190 443512 380196
rect 485976 380186 486004 380559
rect 485964 380180 486016 380186
rect 485964 380122 486016 380128
rect 434352 379568 434404 379574
rect 434352 379510 434404 379516
rect 408316 379500 408368 379506
rect 408316 379442 408368 379448
rect 408328 379409 408356 379442
rect 396078 379400 396134 379409
rect 396078 379335 396134 379344
rect 397090 379400 397146 379409
rect 397090 379335 397146 379344
rect 405830 379400 405886 379409
rect 405830 379335 405886 379344
rect 407578 379400 407634 379409
rect 407578 379335 407634 379344
rect 408314 379400 408370 379409
rect 408314 379335 408370 379344
rect 411258 379400 411314 379409
rect 411258 379335 411314 379344
rect 412362 379400 412418 379409
rect 412362 379335 412418 379344
rect 415674 379400 415730 379409
rect 415674 379335 415730 379344
rect 425978 379400 426034 379409
rect 425978 379335 426034 379344
rect 435178 379400 435234 379409
rect 435178 379335 435234 379344
rect 437846 379400 437902 379409
rect 437846 379335 437902 379344
rect 445850 379400 445906 379409
rect 445850 379335 445906 379344
rect 447506 379400 447562 379409
rect 447506 379335 447562 379344
rect 451002 379400 451058 379409
rect 451002 379335 451058 379344
rect 453026 379400 453082 379409
rect 453026 379335 453082 379344
rect 455510 379400 455566 379409
rect 455510 379335 455566 379344
rect 458362 379400 458418 379409
rect 458362 379335 458418 379344
rect 460938 379400 460994 379409
rect 460938 379335 460994 379344
rect 474830 379400 474886 379409
rect 474830 379335 474886 379344
rect 396092 378894 396120 379335
rect 397104 379030 397132 379335
rect 399482 379264 399538 379273
rect 399482 379199 399538 379208
rect 400402 379264 400458 379273
rect 400402 379199 400458 379208
rect 402978 379264 403034 379273
rect 402978 379199 403034 379208
rect 397092 379024 397144 379030
rect 397092 378966 397144 378972
rect 396080 378888 396132 378894
rect 396080 378830 396132 378836
rect 399496 378690 399524 379199
rect 400416 378758 400444 379199
rect 400404 378752 400456 378758
rect 400404 378694 400456 378700
rect 399484 378684 399536 378690
rect 399484 378626 399536 378632
rect 402992 377262 403020 379199
rect 405844 378622 405872 379335
rect 405832 378616 405884 378622
rect 405832 378558 405884 378564
rect 407592 378418 407620 379335
rect 409970 379264 410026 379273
rect 409970 379199 410026 379208
rect 407580 378412 407632 378418
rect 407580 378354 407632 378360
rect 408682 378176 408738 378185
rect 408682 378111 408738 378120
rect 402980 377256 403032 377262
rect 402980 377198 403032 377204
rect 381360 377188 381412 377194
rect 381360 377130 381412 377136
rect 408696 375086 408724 378111
rect 409984 377330 410012 379199
rect 411272 378486 411300 379335
rect 412376 378554 412404 379335
rect 413282 378584 413338 378593
rect 412364 378548 412416 378554
rect 413282 378519 413338 378528
rect 414570 378584 414626 378593
rect 414570 378519 414626 378528
rect 412364 378490 412416 378496
rect 411260 378480 411312 378486
rect 411260 378422 411312 378428
rect 409972 377324 410024 377330
rect 409972 377266 410024 377272
rect 413296 376106 413324 378519
rect 413284 376100 413336 376106
rect 413284 376042 413336 376048
rect 414584 375970 414612 378519
rect 415688 377534 415716 379335
rect 415858 379264 415914 379273
rect 415858 379199 415914 379208
rect 416870 379264 416926 379273
rect 416870 379199 416926 379208
rect 422850 379264 422906 379273
rect 422850 379199 422906 379208
rect 415676 377528 415728 377534
rect 415676 377470 415728 377476
rect 415872 377398 415900 379199
rect 416884 377466 416912 379199
rect 418434 378584 418490 378593
rect 418434 378519 418490 378528
rect 418158 378176 418214 378185
rect 418158 378111 418214 378120
rect 416872 377460 416924 377466
rect 416872 377402 416924 377408
rect 415860 377392 415912 377398
rect 415860 377334 415912 377340
rect 414572 375964 414624 375970
rect 414572 375906 414624 375912
rect 408684 375080 408736 375086
rect 408684 375022 408736 375028
rect 418172 375018 418200 378111
rect 418448 376038 418476 378519
rect 420642 378176 420698 378185
rect 420642 378111 420698 378120
rect 421194 378176 421250 378185
rect 421194 378111 421250 378120
rect 422666 378176 422722 378185
rect 422666 378111 422722 378120
rect 418436 376032 418488 376038
rect 418436 375974 418488 375980
rect 420656 375154 420684 378111
rect 421208 375222 421236 378111
rect 421196 375216 421248 375222
rect 421196 375158 421248 375164
rect 420644 375148 420696 375154
rect 420644 375090 420696 375096
rect 418160 375012 418212 375018
rect 418160 374954 418212 374960
rect 422680 374882 422708 378111
rect 422864 376174 422892 379199
rect 423954 378176 424010 378185
rect 423954 378111 424010 378120
rect 425150 378176 425206 378185
rect 425150 378111 425206 378120
rect 422852 376168 422904 376174
rect 422852 376110 422904 376116
rect 423968 374950 423996 378111
rect 425164 375290 425192 378111
rect 425992 377602 426020 379335
rect 430670 378856 430726 378865
rect 430670 378791 430726 378800
rect 428554 378176 428610 378185
rect 428554 378111 428610 378120
rect 429658 378176 429714 378185
rect 429658 378111 429714 378120
rect 425980 377596 426032 377602
rect 425980 377538 426032 377544
rect 425152 375284 425204 375290
rect 425152 375226 425204 375232
rect 423956 374944 424008 374950
rect 423956 374886 424008 374892
rect 422668 374876 422720 374882
rect 422668 374818 422720 374824
rect 428568 374746 428596 378111
rect 429672 374814 429700 378111
rect 430684 376310 430712 378791
rect 435192 378350 435220 379335
rect 437860 378826 437888 379335
rect 437848 378820 437900 378826
rect 437848 378762 437900 378768
rect 436190 378720 436246 378729
rect 436190 378655 436246 378664
rect 435180 378344 435232 378350
rect 432234 378312 432290 378321
rect 435180 378286 435232 378292
rect 432234 378247 432290 378256
rect 430672 376304 430724 376310
rect 430672 376246 430724 376252
rect 432248 375358 432276 378247
rect 436204 376242 436232 378655
rect 439042 378176 439098 378185
rect 439042 378111 439098 378120
rect 436192 376236 436244 376242
rect 436192 376178 436244 376184
rect 432236 375352 432288 375358
rect 432236 375294 432288 375300
rect 429660 374808 429712 374814
rect 429660 374750 429712 374756
rect 428556 374740 428608 374746
rect 428556 374682 428608 374688
rect 439056 374678 439084 378111
rect 445864 377942 445892 379335
rect 445852 377936 445904 377942
rect 445852 377878 445904 377884
rect 447520 377670 447548 379335
rect 451016 377874 451044 379335
rect 451004 377868 451056 377874
rect 451004 377810 451056 377816
rect 453040 377806 453068 379335
rect 453028 377800 453080 377806
rect 453028 377742 453080 377748
rect 455524 377738 455552 379335
rect 458376 378010 458404 379335
rect 460952 378078 460980 379335
rect 463514 379264 463570 379273
rect 463514 379199 463570 379208
rect 473450 379264 473506 379273
rect 473450 379199 473506 379208
rect 460940 378072 460992 378078
rect 460940 378014 460992 378020
rect 458364 378004 458416 378010
rect 458364 377946 458416 377952
rect 455512 377732 455564 377738
rect 455512 377674 455564 377680
rect 447508 377664 447560 377670
rect 447508 377606 447560 377612
rect 463528 376514 463556 379199
rect 465170 378992 465226 379001
rect 465170 378927 465226 378936
rect 465184 376689 465212 378927
rect 470782 378856 470838 378865
rect 470782 378791 470838 378800
rect 467930 378720 467986 378729
rect 467930 378655 467986 378664
rect 465170 376680 465226 376689
rect 465170 376615 465226 376624
rect 463516 376508 463568 376514
rect 463516 376450 463568 376456
rect 467944 376378 467972 378655
rect 470796 376446 470824 378791
rect 473464 376582 473492 379199
rect 474844 378146 474872 379335
rect 503074 379264 503130 379273
rect 503074 379199 503130 379208
rect 503534 379264 503590 379273
rect 503534 379199 503590 379208
rect 477590 378992 477646 379001
rect 477590 378927 477646 378936
rect 474832 378140 474884 378146
rect 474832 378082 474884 378088
rect 477604 376718 477632 378927
rect 483386 378856 483442 378865
rect 483386 378791 483442 378800
rect 477592 376712 477644 376718
rect 477592 376654 477644 376660
rect 483400 376650 483428 378791
rect 503088 378282 503116 379199
rect 503076 378276 503128 378282
rect 503076 378218 503128 378224
rect 503548 378214 503576 379199
rect 503536 378208 503588 378214
rect 503536 378150 503588 378156
rect 483388 376644 483440 376650
rect 483388 376586 483440 376592
rect 473452 376576 473504 376582
rect 473452 376518 473504 376524
rect 470784 376440 470836 376446
rect 470784 376382 470836 376388
rect 467932 376372 467984 376378
rect 467932 376314 467984 376320
rect 439044 374672 439096 374678
rect 439044 374614 439096 374620
rect 500408 359644 500460 359650
rect 500408 359586 500460 359592
rect 498936 359576 498988 359582
rect 498936 359518 498988 359524
rect 498948 358873 498976 359518
rect 500420 358873 500448 359586
rect 498934 358864 498990 358873
rect 498934 358799 498990 358808
rect 500406 358864 500462 358873
rect 500406 358799 500462 358808
rect 510894 358864 510950 358873
rect 517532 358834 517560 466482
rect 517612 378276 517664 378282
rect 517612 378218 517664 378224
rect 510894 358799 510896 358808
rect 510948 358799 510950 358808
rect 517520 358828 517572 358834
rect 510896 358770 510948 358776
rect 517520 358770 517572 358776
rect 381268 358012 381320 358018
rect 381268 357954 381320 357960
rect 380900 357876 380952 357882
rect 380900 357818 380952 357824
rect 426438 273864 426494 273873
rect 426438 273799 426494 273808
rect 426452 273630 426480 273799
rect 426440 273624 426492 273630
rect 421102 273592 421158 273601
rect 426440 273566 426492 273572
rect 431130 273592 431186 273601
rect 421102 273527 421104 273536
rect 421156 273527 421158 273536
rect 431130 273527 431186 273536
rect 433338 273592 433394 273601
rect 433338 273527 433394 273536
rect 453394 273592 453450 273601
rect 453394 273527 453450 273536
rect 421104 273498 421156 273504
rect 431144 273494 431172 273527
rect 431132 273488 431184 273494
rect 430946 273456 431002 273465
rect 431132 273430 431184 273436
rect 433352 273426 433380 273527
rect 430946 273391 431002 273400
rect 433340 273420 433392 273426
rect 430960 273358 430988 273391
rect 433340 273362 433392 273368
rect 430948 273352 431000 273358
rect 430948 273294 431000 273300
rect 453408 273290 453436 273527
rect 453396 273284 453448 273290
rect 453396 273226 453448 273232
rect 422852 273216 422904 273222
rect 422666 273184 422722 273193
rect 422666 273119 422722 273128
rect 422850 273184 422852 273193
rect 422904 273184 422906 273193
rect 422850 273119 422906 273128
rect 423402 273184 423458 273193
rect 423402 273119 423458 273128
rect 425978 273184 426034 273193
rect 425978 273119 425980 273128
rect 422680 272921 422708 273119
rect 423416 273086 423444 273119
rect 426032 273119 426034 273128
rect 425980 273090 426032 273096
rect 423404 273080 423456 273086
rect 423404 273022 423456 273028
rect 468482 273048 468538 273057
rect 468482 272983 468484 272992
rect 468536 272983 468538 272992
rect 470874 273048 470930 273057
rect 470874 272983 470930 272992
rect 468484 272954 468536 272960
rect 470888 272950 470916 272983
rect 470876 272944 470928 272950
rect 422666 272912 422722 272921
rect 470876 272886 470928 272892
rect 473450 272912 473506 272921
rect 422666 272847 422722 272856
rect 473450 272847 473452 272856
rect 473504 272847 473506 272856
rect 475842 272912 475898 272921
rect 475842 272847 475898 272856
rect 473452 272818 473504 272824
rect 475856 272814 475884 272847
rect 475844 272808 475896 272814
rect 475844 272750 475896 272756
rect 478418 272776 478474 272785
rect 478418 272711 478420 272720
rect 478472 272711 478474 272720
rect 480810 272776 480866 272785
rect 480810 272711 480866 272720
rect 478420 272682 478472 272688
rect 480824 272678 480852 272711
rect 480812 272672 480864 272678
rect 380070 272640 380126 272649
rect 480812 272614 480864 272620
rect 483202 272640 483258 272649
rect 380070 272575 380126 272584
rect 483202 272575 483204 272584
rect 379980 269000 380032 269006
rect 379980 268942 380032 268948
rect 379992 258074 380020 268942
rect 380084 267646 380112 272575
rect 483256 272575 483258 272584
rect 485962 272640 486018 272649
rect 485962 272575 486018 272584
rect 483204 272546 483256 272552
rect 485976 272542 486004 272575
rect 485964 272536 486016 272542
rect 423770 272504 423826 272513
rect 485964 272478 486016 272484
rect 423770 272439 423772 272448
rect 423824 272439 423826 272448
rect 423772 272410 423824 272416
rect 401690 272232 401746 272241
rect 401690 272167 401746 272176
rect 415858 272232 415914 272241
rect 415858 272167 415914 272176
rect 416042 272232 416098 272241
rect 416042 272167 416098 272176
rect 455786 272232 455842 272241
rect 455786 272167 455842 272176
rect 396724 271924 396776 271930
rect 396724 271866 396776 271872
rect 380162 271144 380218 271153
rect 380162 271079 380218 271088
rect 380176 269686 380204 271079
rect 380532 270428 380584 270434
rect 380532 270370 380584 270376
rect 380164 269680 380216 269686
rect 380164 269622 380216 269628
rect 380544 269618 380572 270370
rect 391940 269748 391992 269754
rect 391940 269690 391992 269696
rect 380532 269612 380584 269618
rect 380532 269554 380584 269560
rect 387890 269376 387946 269385
rect 387890 269311 387946 269320
rect 387904 268938 387932 269311
rect 390558 269240 390614 269249
rect 390558 269175 390614 269184
rect 387892 268932 387944 268938
rect 387892 268874 387944 268880
rect 390572 268734 390600 269175
rect 390560 268728 390612 268734
rect 390560 268670 390612 268676
rect 391952 268666 391980 269690
rect 391940 268660 391992 268666
rect 391940 268602 391992 268608
rect 380072 267640 380124 267646
rect 380072 267582 380124 267588
rect 380084 266422 380112 267582
rect 380072 266416 380124 266422
rect 380072 266358 380124 266364
rect 379900 258046 380020 258074
rect 379796 148912 379848 148918
rect 379796 148854 379848 148860
rect 379808 147694 379836 148854
rect 379796 147688 379848 147694
rect 379796 147630 379848 147636
rect 379900 146266 379928 258046
rect 396736 252550 396764 271866
rect 397458 270600 397514 270609
rect 397458 270535 397514 270544
rect 398838 270600 398894 270609
rect 398838 270535 398894 270544
rect 400218 270600 400274 270609
rect 400218 270535 400274 270544
rect 397472 270026 397500 270535
rect 398852 270162 398880 270535
rect 398840 270156 398892 270162
rect 398840 270098 398892 270104
rect 400232 270094 400260 270535
rect 401704 270366 401732 272167
rect 415872 271930 415900 272167
rect 415860 271924 415912 271930
rect 415860 271866 415912 271872
rect 416056 271182 416084 272167
rect 427084 271992 427136 271998
rect 427084 271934 427136 271940
rect 436100 271992 436152 271998
rect 436100 271934 436152 271940
rect 425704 271924 425756 271930
rect 425704 271866 425756 271872
rect 416044 271176 416096 271182
rect 409878 271144 409934 271153
rect 409878 271079 409934 271088
rect 412730 271144 412786 271153
rect 416044 271118 416096 271124
rect 418158 271144 418214 271153
rect 412730 271079 412786 271088
rect 418158 271079 418160 271088
rect 409892 270978 409920 271079
rect 412744 271046 412772 271079
rect 418212 271079 418214 271088
rect 418160 271050 418212 271056
rect 412732 271040 412784 271046
rect 412732 270982 412784 270988
rect 409880 270972 409932 270978
rect 409880 270914 409932 270920
rect 405738 270872 405794 270881
rect 405738 270807 405794 270816
rect 402978 270600 403034 270609
rect 402978 270535 403034 270544
rect 403346 270600 403402 270609
rect 403346 270535 403402 270544
rect 404358 270600 404414 270609
rect 404358 270535 404414 270544
rect 401692 270360 401744 270366
rect 401692 270302 401744 270308
rect 400220 270088 400272 270094
rect 400220 270030 400272 270036
rect 397460 270020 397512 270026
rect 397460 269962 397512 269968
rect 402992 268394 403020 270535
rect 403360 269958 403388 270535
rect 404372 270298 404400 270535
rect 404360 270292 404412 270298
rect 404360 270234 404412 270240
rect 405752 270230 405780 270807
rect 411350 270736 411406 270745
rect 411350 270671 411406 270680
rect 407118 270600 407174 270609
rect 407118 270535 407174 270544
rect 408498 270600 408554 270609
rect 408498 270535 408554 270544
rect 409878 270600 409934 270609
rect 409878 270535 409934 270544
rect 411258 270600 411314 270609
rect 411258 270535 411314 270544
rect 405740 270224 405792 270230
rect 405740 270166 405792 270172
rect 403348 269952 403400 269958
rect 403348 269894 403400 269900
rect 407132 269890 407160 270535
rect 407120 269884 407172 269890
rect 407120 269826 407172 269832
rect 408512 268870 408540 270535
rect 408500 268864 408552 268870
rect 408500 268806 408552 268812
rect 409892 268802 409920 270535
rect 411272 270502 411300 270535
rect 411260 270496 411312 270502
rect 411260 270438 411312 270444
rect 411364 270434 411392 270671
rect 413006 270600 413062 270609
rect 413006 270535 413062 270544
rect 414018 270600 414074 270609
rect 414018 270535 414074 270544
rect 416778 270600 416834 270609
rect 416778 270535 416834 270544
rect 418158 270600 418214 270609
rect 418158 270535 418214 270544
rect 419538 270600 419594 270609
rect 419538 270535 419594 270544
rect 420918 270600 420974 270609
rect 420918 270535 420974 270544
rect 411352 270428 411404 270434
rect 411352 270370 411404 270376
rect 413020 269822 413048 270535
rect 413008 269816 413060 269822
rect 413008 269758 413060 269764
rect 414032 269006 414060 270535
rect 416792 269074 416820 270535
rect 416780 269068 416832 269074
rect 416780 269010 416832 269016
rect 414020 269000 414072 269006
rect 414020 268942 414072 268948
rect 409880 268796 409932 268802
rect 409880 268738 409932 268744
rect 418172 268666 418200 270535
rect 419552 268734 419580 270535
rect 420932 268938 420960 270535
rect 420920 268932 420972 268938
rect 420920 268874 420972 268880
rect 419540 268728 419592 268734
rect 419540 268670 419592 268676
rect 418160 268660 418212 268666
rect 418160 268602 418212 268608
rect 402980 268388 403032 268394
rect 402980 268330 403032 268336
rect 396724 252544 396776 252550
rect 396724 252486 396776 252492
rect 425716 252006 425744 271866
rect 427096 252074 427124 271934
rect 427820 271924 427872 271930
rect 427820 271866 427872 271872
rect 427832 271833 427860 271866
rect 436112 271833 436140 271934
rect 455800 271862 455828 272167
rect 455788 271856 455840 271862
rect 427818 271824 427874 271833
rect 427818 271759 427874 271768
rect 433338 271824 433394 271833
rect 433338 271759 433394 271768
rect 436098 271824 436154 271833
rect 436098 271759 436154 271768
rect 437478 271824 437534 271833
rect 437478 271759 437534 271768
rect 442998 271824 443054 271833
rect 442998 271759 443054 271768
rect 445758 271824 445814 271833
rect 445758 271759 445814 271768
rect 447138 271824 447194 271833
rect 447138 271759 447194 271768
rect 449898 271824 449954 271833
rect 455788 271798 455840 271804
rect 458178 271824 458234 271833
rect 449898 271759 449954 271768
rect 458178 271759 458180 271768
rect 433352 271386 433380 271759
rect 437492 271522 437520 271759
rect 443012 271590 443040 271759
rect 443000 271584 443052 271590
rect 443000 271526 443052 271532
rect 437480 271516 437532 271522
rect 437480 271458 437532 271464
rect 445772 271454 445800 271759
rect 447152 271726 447180 271759
rect 447140 271720 447192 271726
rect 447140 271662 447192 271668
rect 449912 271658 449940 271759
rect 458232 271759 458234 271768
rect 458180 271730 458232 271736
rect 503626 271688 503682 271697
rect 449900 271652 449952 271658
rect 503626 271623 503682 271632
rect 449900 271594 449952 271600
rect 445760 271448 445812 271454
rect 440238 271416 440294 271425
rect 433340 271380 433392 271386
rect 445760 271390 445812 271396
rect 440238 271351 440294 271360
rect 433340 271322 433392 271328
rect 440252 271318 440280 271351
rect 503640 271318 503668 271623
rect 440240 271312 440292 271318
rect 434718 271280 434774 271289
rect 503628 271312 503680 271318
rect 440240 271254 440292 271260
rect 503534 271280 503590 271289
rect 434718 271215 434720 271224
rect 434772 271215 434774 271224
rect 503628 271254 503680 271260
rect 503534 271215 503590 271224
rect 434720 271186 434772 271192
rect 503548 271182 503576 271215
rect 503536 271176 503588 271182
rect 503536 271118 503588 271124
rect 431958 270872 432014 270881
rect 431958 270807 432014 270816
rect 433338 270872 433394 270881
rect 433338 270807 433394 270816
rect 437478 270872 437534 270881
rect 437478 270807 437534 270816
rect 438858 270872 438914 270881
rect 438858 270807 438914 270816
rect 429198 270736 429254 270745
rect 429198 270671 429254 270680
rect 427084 252068 427136 252074
rect 427084 252010 427136 252016
rect 425704 252000 425756 252006
rect 425704 251942 425756 251948
rect 429212 251938 429240 270671
rect 429200 251932 429252 251938
rect 429200 251874 429252 251880
rect 431972 251870 432000 270807
rect 433352 267578 433380 270807
rect 437492 267714 437520 270807
rect 437480 267708 437532 267714
rect 437480 267650 437532 267656
rect 438872 267646 438900 270807
rect 438860 267640 438912 267646
rect 438860 267582 438912 267588
rect 433340 267572 433392 267578
rect 433340 267514 433392 267520
rect 500868 253360 500920 253366
rect 500866 253328 500868 253337
rect 500920 253328 500922 253337
rect 499212 253292 499264 253298
rect 500866 253263 500922 253272
rect 499212 253234 499264 253240
rect 499224 252793 499252 253234
rect 499210 252784 499266 252793
rect 499210 252719 499266 252728
rect 510894 252648 510950 252657
rect 517532 252618 517560 358770
rect 517624 271318 517652 378218
rect 517704 378208 517756 378214
rect 517704 378150 517756 378156
rect 517716 271862 517744 378150
rect 517808 359582 517836 466550
rect 517888 466472 517940 466478
rect 517888 466414 517940 466420
rect 517900 364334 517928 466414
rect 518900 465112 518952 465118
rect 518900 465054 518952 465060
rect 518912 459649 518940 465054
rect 519556 460222 519584 524418
rect 560956 511970 560984 586502
rect 580276 577697 580304 634782
rect 580368 630873 580396 639202
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580264 515432 580316 515438
rect 580264 515374 580316 515380
rect 560944 511964 560996 511970
rect 560944 511906 560996 511912
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 520924 495508 520976 495514
rect 520924 495450 520976 495456
rect 519544 460216 519596 460222
rect 519544 460158 519596 460164
rect 518898 459640 518954 459649
rect 518898 459575 518954 459584
rect 519450 459640 519506 459649
rect 519450 459575 519506 459584
rect 519082 400344 519138 400353
rect 519082 400279 519138 400288
rect 518990 398168 519046 398177
rect 518990 398103 519046 398112
rect 519004 364334 519032 398103
rect 519096 366382 519124 400279
rect 519358 396808 519414 396817
rect 519358 396743 519414 396752
rect 519174 395312 519230 395321
rect 519174 395247 519230 395256
rect 519188 369170 519216 395247
rect 519266 394088 519322 394097
rect 519266 394023 519322 394032
rect 519176 369164 519228 369170
rect 519176 369106 519228 369112
rect 519084 366376 519136 366382
rect 519084 366318 519136 366324
rect 517900 364306 518020 364334
rect 517992 359650 518020 364306
rect 518912 364306 519032 364334
rect 518912 363730 518940 364306
rect 518900 363724 518952 363730
rect 518900 363666 518952 363672
rect 517980 359644 518032 359650
rect 517980 359586 518032 359592
rect 517796 359576 517848 359582
rect 517796 359518 517848 359524
rect 517704 271856 517756 271862
rect 517704 271798 517756 271804
rect 517612 271312 517664 271318
rect 517612 271254 517664 271260
rect 510894 252583 510896 252592
rect 510948 252583 510950 252592
rect 517520 252612 517572 252618
rect 510896 252554 510948 252560
rect 517520 252554 517572 252560
rect 431960 251864 432012 251870
rect 431960 251806 432012 251812
rect 421012 167000 421064 167006
rect 421012 166942 421064 166948
rect 418436 166864 418488 166870
rect 418434 166832 418436 166841
rect 421024 166841 421052 166942
rect 423404 166932 423456 166938
rect 423404 166874 423456 166880
rect 423416 166841 423444 166874
rect 418488 166832 418490 166841
rect 418434 166767 418490 166776
rect 421010 166832 421066 166841
rect 421010 166767 421066 166776
rect 423402 166832 423458 166841
rect 423402 166767 423458 166776
rect 428186 166832 428242 166841
rect 428186 166767 428188 166776
rect 428240 166767 428242 166776
rect 445850 166832 445906 166841
rect 445850 166767 445906 166776
rect 470966 166832 471022 166841
rect 470966 166767 471022 166776
rect 475842 166832 475898 166841
rect 475842 166767 475898 166776
rect 478418 166832 478474 166841
rect 478418 166767 478474 166776
rect 480902 166832 480958 166841
rect 480902 166767 480958 166776
rect 428188 166738 428240 166744
rect 445864 166734 445892 166767
rect 445852 166728 445904 166734
rect 445852 166670 445904 166676
rect 470980 166666 471008 166767
rect 470968 166660 471020 166666
rect 470968 166602 471020 166608
rect 475856 166598 475884 166767
rect 475844 166592 475896 166598
rect 475844 166534 475896 166540
rect 478432 166530 478460 166767
rect 478420 166524 478472 166530
rect 478420 166466 478472 166472
rect 480916 166462 480944 166767
rect 483386 166696 483442 166705
rect 483386 166631 483442 166640
rect 485962 166696 486018 166705
rect 485962 166631 486018 166640
rect 480904 166456 480956 166462
rect 480904 166398 480956 166404
rect 483400 166326 483428 166631
rect 485976 166394 486004 166631
rect 503258 166560 503314 166569
rect 503258 166495 503314 166504
rect 485964 166388 486016 166394
rect 485964 166330 486016 166336
rect 483388 166320 483440 166326
rect 483388 166262 483440 166268
rect 436100 165640 436152 165646
rect 380530 165608 380586 165617
rect 380530 165543 380586 165552
rect 397458 165608 397514 165617
rect 397458 165543 397514 165552
rect 401598 165608 401654 165617
rect 401598 165543 401654 165552
rect 404358 165608 404414 165617
rect 404358 165543 404414 165552
rect 409878 165608 409934 165617
rect 409878 165543 409934 165552
rect 415490 165608 415546 165617
rect 415490 165543 415546 165552
rect 416042 165608 416098 165617
rect 416042 165543 416098 165552
rect 418526 165608 418582 165617
rect 418526 165543 418582 165552
rect 423770 165608 423826 165617
rect 423770 165543 423826 165552
rect 433430 165608 433486 165617
rect 433430 165543 433486 165552
rect 434718 165608 434774 165617
rect 434718 165543 434774 165552
rect 436098 165608 436100 165617
rect 436152 165608 436154 165617
rect 436098 165543 436154 165552
rect 437754 165608 437810 165617
rect 437754 165543 437810 165552
rect 438030 165608 438086 165617
rect 438030 165543 438086 165552
rect 440146 165608 440202 165617
rect 442998 165608 443054 165617
rect 440202 165566 440280 165594
rect 440146 165543 440202 165552
rect 380544 165345 380572 165543
rect 380530 165336 380586 165345
rect 380530 165271 380586 165280
rect 396170 164384 396226 164393
rect 396170 164319 396226 164328
rect 396078 164248 396134 164257
rect 396078 164183 396134 164192
rect 396092 163878 396120 164183
rect 396184 163946 396212 164319
rect 396172 163940 396224 163946
rect 396172 163882 396224 163888
rect 396080 163872 396132 163878
rect 396080 163814 396132 163820
rect 379980 162852 380032 162858
rect 379980 162794 380032 162800
rect 379992 162586 380020 162794
rect 379980 162580 380032 162586
rect 379980 162522 380032 162528
rect 379980 148368 380032 148374
rect 379980 148310 380032 148316
rect 379888 146260 379940 146266
rect 379888 146202 379940 146208
rect 379900 56234 379928 146202
rect 379888 56228 379940 56234
rect 379888 56170 379940 56176
rect 379992 54874 380020 148310
rect 396092 145382 396120 163814
rect 396184 145450 396212 163882
rect 396724 161492 396776 161498
rect 396724 161434 396776 161440
rect 396736 146198 396764 161434
rect 397472 148850 397500 165543
rect 398838 164248 398894 164257
rect 398838 164183 398894 164192
rect 400218 164248 400274 164257
rect 400218 164183 400274 164192
rect 397460 148844 397512 148850
rect 397460 148786 397512 148792
rect 398852 148510 398880 164183
rect 400232 148578 400260 164183
rect 400220 148572 400272 148578
rect 400220 148514 400272 148520
rect 398840 148504 398892 148510
rect 398840 148446 398892 148452
rect 401612 148442 401640 165543
rect 402978 164384 403034 164393
rect 402978 164319 403034 164328
rect 401600 148436 401652 148442
rect 401600 148378 401652 148384
rect 396724 146192 396776 146198
rect 396724 146134 396776 146140
rect 402992 145722 403020 164319
rect 403070 164248 403126 164257
rect 403070 164183 403126 164192
rect 403084 145790 403112 164183
rect 404372 145858 404400 165543
rect 407118 164928 407174 164937
rect 409892 164898 409920 165543
rect 407118 164863 407174 164872
rect 409880 164892 409932 164898
rect 407132 164830 407160 164863
rect 409880 164834 409932 164840
rect 407120 164824 407172 164830
rect 407120 164766 407172 164772
rect 412638 164792 412694 164801
rect 412638 164727 412640 164736
rect 412692 164727 412694 164736
rect 412640 164698 412692 164704
rect 411258 164384 411314 164393
rect 411258 164319 411314 164328
rect 405738 164248 405794 164257
rect 405738 164183 405794 164192
rect 407210 164248 407266 164257
rect 407210 164183 407266 164192
rect 408498 164248 408554 164257
rect 408498 164183 408554 164192
rect 409878 164248 409934 164257
rect 409878 164183 409934 164192
rect 404360 145852 404412 145858
rect 404360 145794 404412 145800
rect 403072 145784 403124 145790
rect 403072 145726 403124 145732
rect 402980 145716 403032 145722
rect 402980 145658 403032 145664
rect 405752 145518 405780 164183
rect 407224 145654 407252 164183
rect 408512 145926 408540 164183
rect 409892 145994 409920 164183
rect 409880 145988 409932 145994
rect 409880 145930 409932 145936
rect 408500 145920 408552 145926
rect 408500 145862 408552 145868
rect 407212 145648 407264 145654
rect 407212 145590 407264 145596
rect 405740 145512 405792 145518
rect 405740 145454 405792 145460
rect 396172 145444 396224 145450
rect 396172 145386 396224 145392
rect 396080 145376 396132 145382
rect 396080 145318 396132 145324
rect 411272 145314 411300 164319
rect 411350 164248 411406 164257
rect 411350 164183 411406 164192
rect 412730 164248 412786 164257
rect 412730 164183 412786 164192
rect 414018 164248 414074 164257
rect 414018 164183 414074 164192
rect 411364 146062 411392 164183
rect 412744 146130 412772 164183
rect 414032 146266 414060 164183
rect 414020 146260 414072 146266
rect 414020 146202 414072 146208
rect 412732 146124 412784 146130
rect 412732 146066 412784 146072
rect 411352 146056 411404 146062
rect 415504 146033 415532 165543
rect 416056 164694 416084 165543
rect 416044 164688 416096 164694
rect 416044 164630 416096 164636
rect 416778 164248 416834 164257
rect 416778 164183 416834 164192
rect 418158 164248 418214 164257
rect 418158 164183 418214 164192
rect 416792 146198 416820 164183
rect 418172 162178 418200 164183
rect 418540 162722 418568 165543
rect 419264 165096 419316 165102
rect 419264 165038 419316 165044
rect 419276 164898 419304 165038
rect 419264 164892 419316 164898
rect 419264 164834 419316 164840
rect 420918 164792 420974 164801
rect 420918 164727 420974 164736
rect 419538 164248 419594 164257
rect 419538 164183 419594 164192
rect 418528 162716 418580 162722
rect 418528 162658 418580 162664
rect 419552 162654 419580 164183
rect 420932 162790 420960 164727
rect 423586 164248 423642 164257
rect 423642 164206 423720 164234
rect 423586 164183 423642 164192
rect 420920 162784 420972 162790
rect 420920 162726 420972 162732
rect 419540 162648 419592 162654
rect 419540 162590 419592 162596
rect 418160 162172 418212 162178
rect 418160 162114 418212 162120
rect 416780 146192 416832 146198
rect 416780 146134 416832 146140
rect 411352 145998 411404 146004
rect 415490 146024 415546 146033
rect 415490 145959 415546 145968
rect 423692 145897 423720 164206
rect 423678 145888 423734 145897
rect 423678 145823 423734 145832
rect 423784 145761 423812 165543
rect 433338 164928 433394 164937
rect 433338 164863 433340 164872
rect 433392 164863 433394 164872
rect 433340 164834 433392 164840
rect 433444 164830 433472 165543
rect 434732 164966 434760 165543
rect 434720 164960 434772 164966
rect 434720 164902 434772 164908
rect 428924 164824 428976 164830
rect 433432 164824 433484 164830
rect 428924 164766 428976 164772
rect 430670 164792 430726 164801
rect 426530 164384 426586 164393
rect 426530 164319 426586 164328
rect 426346 164248 426402 164257
rect 426402 164206 426480 164234
rect 426346 164183 426402 164192
rect 423770 145752 423826 145761
rect 423770 145687 423826 145696
rect 426452 145625 426480 164206
rect 426544 164014 426572 164319
rect 427726 164248 427782 164257
rect 427782 164206 427860 164234
rect 427726 164183 427782 164192
rect 426532 164008 426584 164014
rect 426532 163950 426584 163956
rect 427832 148918 427860 164206
rect 428936 162858 428964 164766
rect 433432 164766 433484 164772
rect 430670 164727 430726 164736
rect 429290 164384 429346 164393
rect 429290 164319 429346 164328
rect 429106 164248 429162 164257
rect 429162 164206 429240 164234
rect 429106 164183 429162 164192
rect 428924 162852 428976 162858
rect 428924 162794 428976 162800
rect 427820 148912 427872 148918
rect 427820 148854 427872 148860
rect 429212 148374 429240 164206
rect 429304 163606 429332 164319
rect 430578 164248 430634 164257
rect 430578 164183 430580 164192
rect 430632 164183 430634 164192
rect 430580 164154 430632 164160
rect 429292 163600 429344 163606
rect 429292 163542 429344 163548
rect 430684 163538 430712 164727
rect 431958 164248 432014 164257
rect 431958 164183 432014 164192
rect 434626 164248 434682 164257
rect 434810 164248 434866 164257
rect 434682 164206 434760 164234
rect 434626 164183 434682 164192
rect 431972 164082 432000 164183
rect 431960 164076 432012 164082
rect 431960 164018 432012 164024
rect 430672 163532 430724 163538
rect 430672 163474 430724 163480
rect 434732 148986 434760 164206
rect 434810 164183 434866 164192
rect 434824 164150 434852 164183
rect 434812 164144 434864 164150
rect 434812 164086 434864 164092
rect 437768 162761 437796 165543
rect 438044 165170 438072 165543
rect 438032 165164 438084 165170
rect 438032 165106 438084 165112
rect 437754 162752 437810 162761
rect 437754 162687 437810 162696
rect 440252 149054 440280 165566
rect 442998 165543 443054 165552
rect 447322 165608 447378 165617
rect 447322 165543 447378 165552
rect 449898 165608 449954 165617
rect 449898 165543 449954 165552
rect 452658 165608 452714 165617
rect 452658 165543 452714 165552
rect 455418 165608 455474 165617
rect 455418 165543 455420 165552
rect 443012 165442 443040 165543
rect 443000 165436 443052 165442
rect 443000 165378 443052 165384
rect 447336 165238 447364 165543
rect 449912 165306 449940 165543
rect 452672 165374 452700 165543
rect 455472 165543 455474 165552
rect 458362 165608 458418 165617
rect 458362 165543 458418 165552
rect 455420 165514 455472 165520
rect 458376 165510 458404 165543
rect 458364 165504 458416 165510
rect 458364 165446 458416 165452
rect 452660 165368 452712 165374
rect 452660 165310 452712 165316
rect 449900 165300 449952 165306
rect 449900 165242 449952 165248
rect 447324 165232 447376 165238
rect 447324 165174 447376 165180
rect 503272 165102 503300 166495
rect 503350 165608 503406 165617
rect 503350 165543 503406 165552
rect 503260 165096 503312 165102
rect 440330 165064 440386 165073
rect 503260 165038 503312 165044
rect 440330 164999 440332 165008
rect 440384 164999 440386 165008
rect 440332 164970 440384 164976
rect 503364 164966 503392 165543
rect 517532 164966 517560 252554
rect 517624 165918 517652 271254
rect 517704 253360 517756 253366
rect 517704 253302 517756 253308
rect 517716 253230 517744 253302
rect 517808 253298 517836 359518
rect 517888 271856 517940 271862
rect 517888 271798 517940 271804
rect 517900 271182 517928 271798
rect 517888 271176 517940 271182
rect 517888 271118 517940 271124
rect 517796 253292 517848 253298
rect 517796 253234 517848 253240
rect 517704 253224 517756 253230
rect 517704 253166 517756 253172
rect 517612 165912 517664 165918
rect 517612 165854 517664 165860
rect 517612 165572 517664 165578
rect 517612 165514 517664 165520
rect 503352 164960 503404 164966
rect 503352 164902 503404 164908
rect 510528 164960 510580 164966
rect 510528 164902 510580 164908
rect 517520 164960 517572 164966
rect 517520 164902 517572 164908
rect 440240 149048 440292 149054
rect 440240 148990 440292 148996
rect 434720 148980 434772 148986
rect 434720 148922 434772 148928
rect 429200 148368 429252 148374
rect 429200 148310 429252 148316
rect 500224 146192 500276 146198
rect 500224 146134 500276 146140
rect 498660 146124 498712 146130
rect 498660 146066 498712 146072
rect 426438 145616 426494 145625
rect 426438 145551 426494 145560
rect 411260 145308 411312 145314
rect 411260 145250 411312 145256
rect 498672 144945 498700 146066
rect 500236 144945 500264 146134
rect 510540 145586 510568 164902
rect 517624 164898 517652 165514
rect 517612 164892 517664 164898
rect 517612 164834 517664 164840
rect 517520 146124 517572 146130
rect 517520 146066 517572 146072
rect 517532 145654 517560 146066
rect 517520 145648 517572 145654
rect 517520 145590 517572 145596
rect 510528 145580 510580 145586
rect 510528 145522 510580 145528
rect 510540 145466 510568 145522
rect 510618 145480 510674 145489
rect 510540 145438 510618 145466
rect 510618 145415 510674 145424
rect 498658 144936 498714 144945
rect 498658 144871 498714 144880
rect 500222 144936 500278 144945
rect 500222 144871 500278 144880
rect 396078 59800 396134 59809
rect 396078 59735 396134 59744
rect 397090 59800 397146 59809
rect 397090 59735 397146 59744
rect 416962 59800 417018 59809
rect 416962 59735 417018 59744
rect 423494 59800 423550 59809
rect 423494 59735 423550 59744
rect 423954 59800 424010 59809
rect 423954 59735 424010 59744
rect 396092 59702 396120 59735
rect 396080 59696 396132 59702
rect 396080 59638 396132 59644
rect 397104 59634 397132 59735
rect 403070 59664 403126 59673
rect 397092 59628 397144 59634
rect 403070 59599 403126 59608
rect 404174 59664 404230 59673
rect 404174 59599 404230 59608
rect 412546 59664 412602 59673
rect 412546 59599 412602 59608
rect 416042 59664 416098 59673
rect 416042 59599 416098 59608
rect 397092 59570 397144 59576
rect 403084 58478 403112 59599
rect 404188 58614 404216 59599
rect 410706 59528 410762 59537
rect 410706 59463 410762 59472
rect 410720 59294 410748 59463
rect 410708 59288 410760 59294
rect 410708 59230 410760 59236
rect 404176 58608 404228 58614
rect 404176 58550 404228 58556
rect 403072 58472 403124 58478
rect 403072 58414 403124 58420
rect 397458 57896 397514 57905
rect 397458 57831 397514 57840
rect 399482 57896 399538 57905
rect 399482 57831 399538 57840
rect 400218 57896 400274 57905
rect 400218 57831 400274 57840
rect 401690 57896 401746 57905
rect 401690 57831 401746 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407210 57896 407266 57905
rect 407210 57831 407266 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 379980 54868 380032 54874
rect 379980 54810 380032 54816
rect 379704 54800 379756 54806
rect 379704 54742 379756 54748
rect 378048 54732 378100 54738
rect 378048 54674 378100 54680
rect 377312 54664 377364 54670
rect 377312 54606 377364 54612
rect 376484 54528 376536 54534
rect 376484 54470 376536 54476
rect 375564 54460 375616 54466
rect 375564 54402 375616 54408
rect 374276 54392 374328 54398
rect 374276 54334 374328 54340
rect 397472 54330 397500 57831
rect 399496 55894 399524 57831
rect 399484 55888 399536 55894
rect 399484 55830 399536 55836
rect 400232 55146 400260 57831
rect 401704 55962 401732 57831
rect 401692 55956 401744 55962
rect 401692 55898 401744 55904
rect 400220 55140 400272 55146
rect 400220 55082 400272 55088
rect 404372 54534 404400 57831
rect 405844 55214 405872 57831
rect 405832 55208 405884 55214
rect 405832 55150 405884 55156
rect 407224 54602 407252 57831
rect 408328 56574 408356 57831
rect 408316 56568 408368 56574
rect 408316 56510 408368 56516
rect 408696 56098 408724 57831
rect 408684 56092 408736 56098
rect 408684 56034 408736 56040
rect 409892 54670 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 56030 411300 56879
rect 411260 56024 411312 56030
rect 411260 55966 411312 55972
rect 411364 54738 411392 57831
rect 412560 56953 412588 59599
rect 416056 59022 416084 59599
rect 416976 59566 417004 59735
rect 419446 59664 419502 59673
rect 419446 59599 419502 59608
rect 421746 59664 421802 59673
rect 421746 59599 421802 59608
rect 416964 59560 417016 59566
rect 416964 59502 417016 59508
rect 418158 59528 418214 59537
rect 418158 59463 418214 59472
rect 418172 59362 418200 59463
rect 418160 59356 418212 59362
rect 418160 59298 418212 59304
rect 419460 59226 419488 59599
rect 420642 59528 420698 59537
rect 420642 59463 420698 59472
rect 419448 59220 419500 59226
rect 419448 59162 419500 59168
rect 420656 59158 420684 59463
rect 420644 59152 420696 59158
rect 420644 59094 420696 59100
rect 421760 59090 421788 59599
rect 423508 59430 423536 59735
rect 423968 59498 423996 59735
rect 458454 59664 458510 59673
rect 458454 59599 458510 59608
rect 503258 59664 503314 59673
rect 503258 59599 503314 59608
rect 423956 59492 424008 59498
rect 423956 59434 424008 59440
rect 423496 59424 423548 59430
rect 423496 59366 423548 59372
rect 425978 59392 426034 59401
rect 425978 59327 426034 59336
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 453394 59392 453450 59401
rect 453394 59327 453450 59336
rect 421748 59084 421800 59090
rect 421748 59026 421800 59032
rect 416044 59016 416096 59022
rect 416044 58958 416096 58964
rect 425992 58954 426020 59327
rect 425980 58948 426032 58954
rect 425980 58890 426032 58896
rect 428200 58682 428228 59327
rect 453408 58818 453436 59327
rect 458468 58886 458496 59599
rect 475842 58984 475898 58993
rect 475842 58919 475898 58928
rect 458456 58880 458508 58886
rect 458456 58822 458508 58828
rect 453396 58812 453448 58818
rect 453396 58754 453448 58760
rect 475856 58750 475884 58919
rect 475844 58744 475896 58750
rect 475844 58686 475896 58692
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 485964 57928 486016 57934
rect 414570 57896 414626 57905
rect 414570 57831 414626 57840
rect 415490 57896 415546 57905
rect 415490 57831 415546 57840
rect 426530 57896 426586 57905
rect 426530 57831 426586 57840
rect 427634 57896 427690 57905
rect 427634 57831 427690 57840
rect 427818 57896 427874 57905
rect 427818 57831 427874 57840
rect 429198 57896 429254 57905
rect 429198 57831 429254 57840
rect 430578 57896 430634 57905
rect 430578 57831 430634 57840
rect 432234 57896 432290 57905
rect 432234 57831 432290 57840
rect 434442 57896 434498 57905
rect 434442 57831 434498 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 436282 57896 436338 57905
rect 436282 57831 436338 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 445850 57896 445906 57905
rect 445850 57831 445906 57840
rect 451002 57896 451058 57905
rect 451002 57831 451058 57840
rect 460938 57896 460994 57905
rect 460938 57831 460994 57840
rect 465906 57896 465962 57905
rect 465906 57831 465962 57840
rect 470874 57896 470930 57905
rect 470874 57831 470876 57840
rect 412546 56944 412602 56953
rect 412546 56879 412602 56888
rect 412638 56808 412694 56817
rect 412638 56743 412694 56752
rect 412652 56166 412680 56743
rect 414584 56234 414612 57831
rect 415504 57254 415532 57831
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 414572 56228 414624 56234
rect 414572 56170 414624 56176
rect 412640 56160 412692 56166
rect 412640 56102 412692 56108
rect 426544 54806 426572 57831
rect 427648 56302 427676 57831
rect 427636 56296 427688 56302
rect 427636 56238 427688 56244
rect 427832 54874 427860 57831
rect 429212 54942 429240 57831
rect 430592 55010 430620 57831
rect 430948 57452 431000 57458
rect 430948 57394 431000 57400
rect 430960 57225 430988 57394
rect 430946 57216 431002 57225
rect 430946 57151 431002 57160
rect 432248 56370 432276 57831
rect 433154 57624 433210 57633
rect 433154 57559 433210 57568
rect 433430 57624 433486 57633
rect 433430 57559 433486 57568
rect 433168 57225 433196 57559
rect 433154 57216 433210 57225
rect 433154 57151 433210 57160
rect 432236 56364 432288 56370
rect 432236 56306 432288 56312
rect 433444 55078 433472 57559
rect 434456 56438 434484 57831
rect 434718 57624 434774 57633
rect 434718 57559 434774 57568
rect 434444 56432 434496 56438
rect 434444 56374 434496 56380
rect 433432 55072 433484 55078
rect 433432 55014 433484 55020
rect 430580 55004 430632 55010
rect 430580 54946 430632 54952
rect 429200 54936 429252 54942
rect 429200 54878 429252 54884
rect 427820 54868 427872 54874
rect 427820 54810 427872 54816
rect 426532 54800 426584 54806
rect 426532 54742 426584 54748
rect 411352 54732 411404 54738
rect 411352 54674 411404 54680
rect 409880 54664 409932 54670
rect 409880 54606 409932 54612
rect 407212 54596 407264 54602
rect 407212 54538 407264 54544
rect 404360 54528 404412 54534
rect 404360 54470 404412 54476
rect 434732 54398 434760 57559
rect 435928 57390 435956 57831
rect 435916 57384 435968 57390
rect 435916 57326 435968 57332
rect 436296 56506 436324 57831
rect 437478 57624 437534 57633
rect 437478 57559 437534 57568
rect 436284 56500 436336 56506
rect 436284 56442 436336 56448
rect 437492 54466 437520 57559
rect 438504 57322 438532 57831
rect 445864 57526 445892 57831
rect 451016 57594 451044 57831
rect 460952 57662 460980 57831
rect 465920 57798 465948 57831
rect 470928 57831 470930 57840
rect 478418 57896 478474 57905
rect 478418 57831 478474 57840
rect 485962 57896 485964 57905
rect 486016 57896 486018 57905
rect 503272 57866 503300 59599
rect 517624 57934 517652 164834
rect 517716 146198 517744 253166
rect 517704 146192 517756 146198
rect 517704 146134 517756 146140
rect 517716 145586 517744 146134
rect 517808 146130 517836 253234
rect 517900 165578 517928 271118
rect 517992 253230 518020 359586
rect 518912 292505 518940 363666
rect 519084 362228 519136 362234
rect 519084 362170 519136 362176
rect 519096 296714 519124 362170
rect 519004 296686 519124 296714
rect 518898 292496 518954 292505
rect 518898 292431 518954 292440
rect 519004 287609 519032 296686
rect 519188 288833 519216 369106
rect 519280 362234 519308 394023
rect 519372 371958 519400 396743
rect 519360 371952 519412 371958
rect 519360 371894 519412 371900
rect 519360 366376 519412 366382
rect 519360 366318 519412 366324
rect 519268 362228 519320 362234
rect 519268 362170 519320 362176
rect 519266 352880 519322 352889
rect 519266 352815 519322 352824
rect 519174 288824 519230 288833
rect 519174 288759 519230 288768
rect 518990 287600 519046 287609
rect 518990 287535 519046 287544
rect 519004 287094 519032 287535
rect 518992 287088 519044 287094
rect 518992 287030 519044 287036
rect 517980 253224 518032 253230
rect 517980 253166 518032 253172
rect 518898 186416 518954 186425
rect 518898 186351 518954 186360
rect 517980 165912 518032 165918
rect 517980 165854 518032 165860
rect 517888 165572 517940 165578
rect 517888 165514 517940 165520
rect 517992 165102 518020 165854
rect 517980 165096 518032 165102
rect 517980 165038 518032 165044
rect 517796 146124 517848 146130
rect 517796 146066 517848 146072
rect 517704 145580 517756 145586
rect 517704 145522 517756 145528
rect 503352 57928 503404 57934
rect 503350 57896 503352 57905
rect 517612 57928 517664 57934
rect 503404 57896 503406 57905
rect 485962 57831 486018 57840
rect 503260 57860 503312 57866
rect 470876 57802 470928 57808
rect 465908 57792 465960 57798
rect 465908 57734 465960 57740
rect 478432 57730 478460 57831
rect 517612 57870 517664 57876
rect 517992 57866 518020 165038
rect 518912 79937 518940 186351
rect 519004 180713 519032 287030
rect 519084 183592 519136 183598
rect 519084 183534 519136 183540
rect 518990 180704 519046 180713
rect 518990 180639 519046 180648
rect 518898 79928 518954 79937
rect 518898 79863 518954 79872
rect 519004 74225 519032 180639
rect 519096 78305 519124 183534
rect 519188 181937 519216 288759
rect 519280 246265 519308 352815
rect 519372 293865 519400 366318
rect 519464 352889 519492 459575
rect 520936 396778 520964 495450
rect 580276 458153 580304 515374
rect 580356 460216 580408 460222
rect 580356 460158 580408 460164
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 580368 404977 580396 460158
rect 580354 404968 580410 404977
rect 580354 404903 580410 404912
rect 520924 396772 520976 396778
rect 520924 396714 520976 396720
rect 580356 396772 580408 396778
rect 580356 396714 580408 396720
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580264 378276 580316 378282
rect 580264 378218 580316 378224
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 519544 371952 519596 371958
rect 519544 371894 519596 371900
rect 519450 352880 519506 352889
rect 519450 352815 519506 352824
rect 519358 293856 519414 293865
rect 519358 293791 519414 293800
rect 519266 246256 519322 246265
rect 519266 246191 519322 246200
rect 519174 181928 519230 181937
rect 519174 181863 519230 181872
rect 519280 139369 519308 246191
rect 519372 186425 519400 293791
rect 519556 290329 519584 371894
rect 580276 325281 580304 378218
rect 580368 351937 580396 396714
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 519634 292496 519690 292505
rect 519634 292431 519690 292440
rect 519542 290320 519598 290329
rect 519542 290255 519598 290264
rect 519556 277394 519584 290255
rect 519464 277366 519584 277394
rect 519358 186416 519414 186425
rect 519358 186351 519414 186360
rect 519464 183433 519492 277366
rect 519648 184793 519676 292431
rect 520186 288824 520242 288833
rect 520186 288759 520242 288768
rect 520200 288454 520228 288759
rect 520188 288448 520240 288454
rect 520188 288390 520240 288396
rect 580264 288448 580316 288454
rect 580264 288390 580316 288396
rect 580276 232393 580304 288390
rect 580356 287088 580408 287094
rect 580356 287030 580408 287036
rect 580368 272241 580396 287030
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 519634 184784 519690 184793
rect 519634 184719 519690 184728
rect 520186 184784 520242 184793
rect 520186 184719 520242 184728
rect 520200 183598 520228 184719
rect 520188 183592 520240 183598
rect 520188 183534 520240 183540
rect 580264 183592 580316 183598
rect 580264 183534 580316 183540
rect 520096 183524 520148 183530
rect 520096 183466 520148 183472
rect 520108 183433 520136 183466
rect 519450 183424 519506 183433
rect 519450 183359 519506 183368
rect 520094 183424 520150 183433
rect 520094 183359 520150 183368
rect 519358 181928 519414 181937
rect 519358 181863 519414 181872
rect 519266 139360 519322 139369
rect 519266 139295 519322 139304
rect 519082 78296 519138 78305
rect 519082 78231 519138 78240
rect 519372 75449 519400 181863
rect 519464 76809 519492 183359
rect 580276 152697 580304 183534
rect 580368 183530 580396 192471
rect 580356 183524 580408 183530
rect 580356 183466 580408 183472
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580356 145648 580408 145654
rect 580356 145590 580408 145596
rect 580264 145580 580316 145586
rect 580264 145522 580316 145528
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519450 76800 519506 76809
rect 519450 76735 519506 76744
rect 519358 75440 519414 75449
rect 519358 75375 519414 75384
rect 518990 74216 519046 74225
rect 518990 74151 519046 74160
rect 503350 57831 503406 57840
rect 517980 57860 518032 57866
rect 503260 57802 503312 57808
rect 517980 57802 518032 57808
rect 478420 57724 478472 57730
rect 478420 57666 478472 57672
rect 460940 57656 460992 57662
rect 460940 57598 460992 57604
rect 451004 57588 451056 57594
rect 451004 57530 451056 57536
rect 445852 57520 445904 57526
rect 445852 57462 445904 57468
rect 438492 57316 438544 57322
rect 438492 57258 438544 57264
rect 437480 54460 437532 54466
rect 437480 54402 437532 54408
rect 434720 54392 434772 54398
rect 434720 54334 434772 54340
rect 213276 54324 213328 54330
rect 213276 54266 213328 54272
rect 237380 54324 237432 54330
rect 237380 54266 237432 54272
rect 373724 54324 373776 54330
rect 373724 54266 373776 54272
rect 397460 54324 397512 54330
rect 397460 54266 397512 54272
rect 580276 33153 580304 145522
rect 580368 73001 580396 145590
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 140042 4040 140098 4049
rect 140042 3975 140098 3984
rect 129370 3904 129426 3913
rect 129370 3839 129426 3848
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 584 480 612 3402
rect 125876 2848 125928 2854
rect 125876 2790 125928 2796
rect 125888 480 125916 2790
rect 129384 480 129412 3839
rect 136454 3496 136510 3505
rect 136454 3431 136510 3440
rect 132958 3360 133014 3369
rect 132958 3295 133014 3304
rect 132972 480 133000 3295
rect 136468 480 136496 3431
rect 140056 480 140084 3975
rect 147126 3768 147182 3777
rect 147126 3703 147182 3712
rect 143538 3224 143594 3233
rect 143538 3159 143594 3168
rect 143552 480 143580 3159
rect 147140 480 147168 3703
rect 150622 3632 150678 3641
rect 150622 3567 150678 3576
rect 150636 480 150664 3567
rect 365718 3224 365774 3233
rect 365718 3159 365774 3168
rect 365732 2854 365760 3159
rect 365720 2848 365772 2854
rect 365720 2790 365772 2796
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 684256 3570 684312
rect 2962 410488 3018 410544
rect 3514 632032 3570 632088
rect 3514 547984 3570 548040
rect 3514 514800 3570 514856
rect 3514 482160 3570 482216
rect 3422 201864 3478 201920
rect 2778 97552 2834 97608
rect 3790 579944 3846 580000
rect 3790 462576 3846 462632
rect 3698 358400 3754 358456
rect 3606 306176 3662 306232
rect 3514 58520 3570 58576
rect 57610 635568 57666 635624
rect 57518 626728 57574 626784
rect 57426 604968 57482 605024
rect 57242 598848 57298 598904
rect 57150 596128 57206 596184
rect 57058 590008 57114 590064
rect 57334 586608 57390 586664
rect 57702 614488 57758 614544
rect 57702 602248 57758 602304
rect 57702 580488 57758 580544
rect 59082 632848 59138 632904
rect 58898 623328 58954 623384
rect 57886 611088 57942 611144
rect 58806 608368 58862 608424
rect 58714 592728 58770 592784
rect 58530 583888 58586 583944
rect 58990 617208 59046 617264
rect 59266 629448 59322 629504
rect 59174 620608 59230 620664
rect 120814 613264 120870 613320
rect 59542 577732 59598 577788
rect 120722 576816 120778 576872
rect 121090 598168 121146 598224
rect 121734 628768 121790 628824
rect 121642 622648 121698 622704
rect 121826 616528 121882 616584
rect 122010 601568 122066 601624
rect 121918 579808 121974 579864
rect 122102 595448 122158 595504
rect 122194 592048 122250 592104
rect 122286 589328 122342 589384
rect 122930 634888 122986 634944
rect 123022 632168 123078 632224
rect 123114 626048 123170 626104
rect 123206 619928 123262 619984
rect 123390 610408 123446 610464
rect 123482 607688 123538 607744
rect 124126 604288 124182 604344
rect 123482 585928 123538 585984
rect 123574 583208 123630 583264
rect 147126 635568 147182 635624
rect 146298 626728 146354 626784
rect 146298 623328 146354 623384
rect 147218 614488 147274 614544
rect 146206 611088 146262 611144
rect 146298 604968 146354 605024
rect 147126 602248 147182 602304
rect 146298 592728 146354 592784
rect 146298 590008 146354 590064
rect 146298 586608 146354 586664
rect 147034 583888 147090 583944
rect 147218 596128 147274 596184
rect 147494 629448 147550 629504
rect 147402 620608 147458 620664
rect 148598 632848 148654 632904
rect 148414 608368 148470 608424
rect 148506 598848 148562 598904
rect 148690 617208 148746 617264
rect 149610 577732 149666 577788
rect 149794 580452 149850 580508
rect 211158 635160 211214 635216
rect 210790 585384 210846 585440
rect 210882 580080 210938 580136
rect 210974 576816 211030 576872
rect 212538 628224 212594 628280
rect 211250 625640 211306 625696
rect 211434 619656 211490 619712
rect 211342 615984 211398 616040
rect 211710 601024 211766 601080
rect 211618 597624 211674 597680
rect 211526 594904 211582 594960
rect 211802 592320 211858 592376
rect 212814 632440 212870 632496
rect 212722 622376 212778 622432
rect 213090 613264 213146 613320
rect 212906 610000 212962 610056
rect 212998 607280 213054 607336
rect 213182 589600 213238 589656
rect 213274 582664 213330 582720
rect 214010 603744 214066 603800
rect 237378 635704 237434 635760
rect 237378 629448 237434 629504
rect 237378 626728 237434 626784
rect 237378 623328 237434 623384
rect 237378 620608 237434 620664
rect 237378 617208 237434 617264
rect 238022 611088 238078 611144
rect 237378 608368 237434 608424
rect 237378 604968 237434 605024
rect 237378 602248 237434 602304
rect 237378 598848 237434 598904
rect 237378 596128 237434 596184
rect 237378 592728 237434 592784
rect 237378 590008 237434 590064
rect 237378 586608 237434 586664
rect 237378 583888 237434 583944
rect 237378 580488 237434 580544
rect 237378 577768 237434 577824
rect 238298 632848 238354 632904
rect 238942 614488 238998 614544
rect 300858 635160 300914 635216
rect 300674 576816 300730 576872
rect 238666 550024 238722 550080
rect 248694 549616 248750 549672
rect 255134 549752 255190 549808
rect 300950 632440 301006 632496
rect 302238 628224 302294 628280
rect 301042 625640 301098 625696
rect 301134 619656 301190 619712
rect 301318 610000 301374 610056
rect 301226 601024 301282 601080
rect 294510 549480 294566 549536
rect 293130 549344 293186 549400
rect 301410 592320 301466 592376
rect 301502 589600 301558 589656
rect 301594 582664 301650 582720
rect 302330 622376 302386 622432
rect 302422 615984 302478 616040
rect 302514 613264 302570 613320
rect 302698 607280 302754 607336
rect 302606 597624 302662 597680
rect 302882 603744 302938 603800
rect 303158 603764 303214 603800
rect 303158 603744 303160 603764
rect 303160 603744 303212 603764
rect 303212 603744 303214 603764
rect 302790 594904 302846 594960
rect 302974 585384 303030 585440
rect 303066 580080 303122 580136
rect 298098 549888 298154 549944
rect 300398 549616 300454 549672
rect 301686 550024 301742 550080
rect 301502 549344 301558 549400
rect 300398 528400 300454 528456
rect 301686 528264 301742 528320
rect 302790 540368 302846 540424
rect 302882 525408 302938 525464
rect 57886 517928 57942 517984
rect 42246 479440 42302 479496
rect 42338 476720 42394 476776
rect 42246 271496 42302 271552
rect 42614 479984 42670 480040
rect 43534 476856 43590 476912
rect 42706 467064 42762 467120
rect 50618 484472 50674 484528
rect 50894 484472 50950 484528
rect 43810 479576 43866 479632
rect 44086 467200 44142 467256
rect 46110 379208 46166 379264
rect 46846 482296 46902 482352
rect 46386 268504 46442 268560
rect 46478 268368 46534 268424
rect 47398 379344 47454 379400
rect 47766 378936 47822 378992
rect 47674 271768 47730 271824
rect 47950 482432 48006 482488
rect 47766 271632 47822 271688
rect 47582 271360 47638 271416
rect 48042 271768 48098 271824
rect 48134 271088 48190 271144
rect 48042 270952 48098 271008
rect 50342 479712 50398 479768
rect 49146 271360 49202 271416
rect 49514 467880 49570 467936
rect 49330 165416 49386 165472
rect 49606 380840 49662 380896
rect 50710 467880 50766 467936
rect 50986 379480 51042 379536
rect 50894 165280 50950 165336
rect 51538 380024 51594 380080
rect 51538 379072 51594 379128
rect 51998 465840 52054 465896
rect 51814 270272 51870 270328
rect 53562 471552 53618 471608
rect 52274 465160 52330 465216
rect 52366 380568 52422 380624
rect 52274 379480 52330 379536
rect 52366 282240 52422 282296
rect 53286 271768 53342 271824
rect 53654 471280 53710 471336
rect 304262 527040 304318 527096
rect 303342 510448 303398 510504
rect 302238 495508 302294 495544
rect 302238 495488 302240 495508
rect 302240 495488 302292 495508
rect 302292 495488 302294 495508
rect 53746 388456 53802 388512
rect 53838 272756 53840 272776
rect 53840 272756 53892 272776
rect 53892 272756 53894 272776
rect 53838 272720 53894 272756
rect 54206 272720 54262 272776
rect 54206 146240 54262 146296
rect 55034 471144 55090 471200
rect 56322 471416 56378 471472
rect 56046 165008 56102 165064
rect 56690 410352 56746 410408
rect 57058 417832 57114 417888
rect 57058 414160 57114 414216
rect 57242 416880 57298 416936
rect 57242 413208 57298 413264
rect 57242 411440 57298 411496
rect 57242 408584 57298 408640
rect 57242 391584 57298 391640
rect 57150 389036 57152 389056
rect 57152 389036 57204 389056
rect 57204 389036 57206 389056
rect 57150 389000 57206 389036
rect 56874 309848 56930 309904
rect 56782 301552 56838 301608
rect 56874 203360 56930 203416
rect 57518 389272 57574 389328
rect 57426 309032 57482 309088
rect 57426 307808 57482 307864
rect 57242 282512 57298 282568
rect 57058 195200 57114 195256
rect 57058 175072 57114 175128
rect 54758 146240 54814 146296
rect 56138 146104 56194 146160
rect 57242 204176 57298 204232
rect 57610 311072 57666 311128
rect 57518 304952 57574 305008
rect 57518 303612 57574 303648
rect 57518 303592 57520 303612
rect 57520 303592 57572 303612
rect 57572 303592 57574 303612
rect 57886 309848 57942 309904
rect 57794 309032 57850 309088
rect 57702 306720 57758 306776
rect 57610 204176 57666 204232
rect 57518 203360 57574 203416
rect 57426 198736 57482 198792
rect 57334 196968 57390 197024
rect 57242 97416 57298 97472
rect 57610 200776 57666 200832
rect 57518 96464 57574 96520
rect 57794 304952 57850 305008
rect 57702 199824 57758 199880
rect 57702 198736 57758 198792
rect 57886 282512 57942 282568
rect 57702 198056 57758 198112
rect 57610 93744 57666 93800
rect 57426 93336 57482 93392
rect 57794 195200 57850 195256
rect 57702 91024 57758 91080
rect 57334 90480 57390 90536
rect 58622 284144 58678 284200
rect 58530 272448 58586 272504
rect 58714 281968 58770 282024
rect 57886 175752 57942 175808
rect 57794 88168 57850 88224
rect 57610 70080 57666 70136
rect 58162 164076 58218 164112
rect 58162 164056 58164 164076
rect 58164 164056 58216 164076
rect 58216 164056 58218 164076
rect 58806 177520 58862 177576
rect 58070 147736 58126 147792
rect 58714 145696 58770 145752
rect 57886 68856 57942 68912
rect 3422 19352 3478 19408
rect 58898 145560 58954 145616
rect 59542 388456 59598 388512
rect 59542 377984 59598 378040
rect 59818 272584 59874 272640
rect 59818 271088 59874 271144
rect 59818 270544 59874 270600
rect 63222 485288 63278 485344
rect 63222 484744 63278 484800
rect 65430 485560 65486 485616
rect 65430 485288 65486 485344
rect 66350 482704 66406 482760
rect 68926 484880 68982 484936
rect 67822 468288 67878 468344
rect 69110 468968 69166 469024
rect 69202 468832 69258 468888
rect 69018 466384 69074 466440
rect 70490 467064 70546 467120
rect 72514 485560 72570 485616
rect 71870 467200 71926 467256
rect 71778 466248 71834 466304
rect 73342 485560 73398 485616
rect 73250 485424 73306 485480
rect 73802 485288 73858 485344
rect 73158 469104 73214 469160
rect 74262 484744 74318 484800
rect 74630 466112 74686 466168
rect 74538 465840 74594 465896
rect 76010 485696 76066 485752
rect 77758 485424 77814 485480
rect 77298 485152 77354 485208
rect 78678 485560 78734 485616
rect 78678 468696 78734 468752
rect 80518 479984 80574 480040
rect 78862 468560 78918 468616
rect 84290 471552 84346 471608
rect 81530 469784 81586 469840
rect 85762 471280 85818 471336
rect 88522 471416 88578 471472
rect 88430 471144 88486 471200
rect 76010 465976 76066 466032
rect 91374 485016 91430 485072
rect 74722 465704 74778 465760
rect 67638 465568 67694 465624
rect 94042 468424 94098 468480
rect 118698 479848 118754 479904
rect 121366 482568 121422 482624
rect 120446 482432 120502 482488
rect 118790 479576 118846 479632
rect 121918 479712 121974 479768
rect 122378 479440 122434 479496
rect 124218 477128 124274 477184
rect 124954 476856 125010 476912
rect 124494 476720 124550 476776
rect 125782 476992 125838 477048
rect 127070 482296 127126 482352
rect 128358 477264 128414 477320
rect 145654 485288 145710 485344
rect 145470 485016 145526 485072
rect 144366 483656 144422 483712
rect 145746 472504 145802 472560
rect 147586 485152 147642 485208
rect 146666 479576 146722 479632
rect 147770 478080 147826 478136
rect 147678 472640 147734 472696
rect 152738 479440 152794 479496
rect 151818 478216 151874 478272
rect 151358 476720 151414 476776
rect 150438 474000 150494 474056
rect 155866 483792 155922 483848
rect 155222 482296 155278 482352
rect 154486 480800 154542 480856
rect 157522 476856 157578 476912
rect 156786 475496 156842 475552
rect 155958 474136 156014 474192
rect 160098 468696 160154 468752
rect 163686 485424 163742 485480
rect 162490 471144 162546 471200
rect 161478 468560 161534 468616
rect 153198 467064 153254 467120
rect 165618 465976 165674 466032
rect 171138 485560 171194 485616
rect 170310 478352 170366 478408
rect 169850 472776 169906 472832
rect 169758 468832 169814 468888
rect 168378 468424 168434 468480
rect 172426 480936 172482 480992
rect 171230 471552 171286 471608
rect 171138 468968 171194 469024
rect 170402 466112 170458 466168
rect 172702 471280 172758 471336
rect 172610 467200 172666 467256
rect 174818 471688 174874 471744
rect 178682 479712 178738 479768
rect 178038 466556 178040 466576
rect 178040 466556 178092 466576
rect 178092 466556 178094 466576
rect 178038 466520 178094 466556
rect 180154 466928 180210 466984
rect 166998 465840 167054 465896
rect 162858 465704 162914 465760
rect 182270 471416 182326 471472
rect 185674 484880 185730 484936
rect 187054 485696 187110 485752
rect 190918 466520 190974 466576
rect 187698 464344 187754 464400
rect 110970 380704 111026 380760
rect 113546 380704 113602 380760
rect 116030 380704 116086 380760
rect 118422 380704 118478 380760
rect 120998 380704 121054 380760
rect 123482 380704 123538 380760
rect 125966 380704 126022 380760
rect 131026 380704 131082 380760
rect 133510 380704 133566 380760
rect 140962 380704 141018 380760
rect 143538 380704 143594 380760
rect 146022 380704 146078 380760
rect 155958 380724 156014 380760
rect 155958 380704 155960 380724
rect 155960 380704 156012 380724
rect 156012 380704 156014 380724
rect 158534 380704 158590 380760
rect 160926 380704 160982 380760
rect 163410 380704 163466 380760
rect 165986 380704 166042 380760
rect 128358 380196 128360 380216
rect 128360 380196 128412 380216
rect 128412 380196 128414 380216
rect 128358 380160 128414 380196
rect 85486 379344 85542 379400
rect 86590 379344 86646 379400
rect 87878 379344 87934 379400
rect 88338 379380 88340 379400
rect 88340 379380 88392 379400
rect 88392 379380 88394 379400
rect 88338 379344 88394 379380
rect 88798 379364 88854 379400
rect 88798 379344 88800 379364
rect 88800 379344 88852 379364
rect 88852 379344 88854 379364
rect 80426 379208 80482 379264
rect 77206 378936 77262 378992
rect 83278 378800 83334 378856
rect 80426 378256 80482 378312
rect 90086 379344 90142 379400
rect 90638 379344 90694 379400
rect 91374 379344 91430 379400
rect 92386 379380 92388 379400
rect 92388 379380 92440 379400
rect 92440 379380 92442 379400
rect 92386 379344 92442 379380
rect 93582 379344 93638 379400
rect 96066 379344 96122 379400
rect 98274 379344 98330 379400
rect 98458 379344 98514 379400
rect 101034 379344 101090 379400
rect 103518 379344 103574 379400
rect 104898 379344 104954 379400
rect 108210 379344 108266 379400
rect 108854 379344 108910 379400
rect 111338 379344 111394 379400
rect 112350 379344 112406 379400
rect 113454 379344 113510 379400
rect 114466 379344 114522 379400
rect 115846 379344 115902 379400
rect 135902 379344 135958 379400
rect 138478 379344 138534 379400
rect 150990 379344 151046 379400
rect 154026 379344 154082 379400
rect 93490 379208 93546 379264
rect 95974 379208 96030 379264
rect 94686 378936 94742 378992
rect 84382 378120 84438 378176
rect 97814 378528 97870 378584
rect 99470 379208 99526 379264
rect 102966 379208 103022 379264
rect 100850 378528 100906 378584
rect 101862 378120 101918 378176
rect 105726 378392 105782 378448
rect 106462 378120 106518 378176
rect 107566 378120 107622 378176
rect 148690 378936 148746 378992
rect 183466 378936 183522 378992
rect 182270 378392 182326 378448
rect 178590 358828 178646 358864
rect 178590 358808 178592 358828
rect 178592 358808 178644 358828
rect 178644 358808 178646 358828
rect 180154 358808 180210 358864
rect 197358 484880 197414 484936
rect 197450 484744 197506 484800
rect 190918 358808 190974 358864
rect 113362 273808 113418 273864
rect 61566 273264 61622 273320
rect 61106 272992 61162 273048
rect 60922 272584 60978 272640
rect 60738 272448 60794 272504
rect 60738 252456 60794 252512
rect 61474 272892 61476 272912
rect 61476 272892 61528 272912
rect 61528 272892 61530 272912
rect 61474 272856 61530 272892
rect 61106 271496 61162 271552
rect 76010 273128 76066 273184
rect 77114 273128 77170 273184
rect 83002 273128 83058 273184
rect 90730 273128 90786 273184
rect 93674 273128 93730 273184
rect 95882 273128 95938 273184
rect 95882 272720 95938 272776
rect 96066 273128 96122 273184
rect 96066 272720 96122 272776
rect 98458 272720 98514 272776
rect 87602 272312 87658 272368
rect 94410 272332 94466 272368
rect 94410 272312 94412 272332
rect 94412 272312 94464 272332
rect 94464 272312 94466 272332
rect 61566 271088 61622 271144
rect 62118 271088 62174 271144
rect 84198 271768 84254 271824
rect 77298 270972 77354 271008
rect 77298 270952 77300 270972
rect 77300 270952 77352 270972
rect 77352 270952 77354 270972
rect 62210 270544 62266 270600
rect 84658 271632 84714 271688
rect 77390 268504 77446 268560
rect 85578 270544 85634 270600
rect 96618 271768 96674 271824
rect 99378 272196 99434 272232
rect 99378 272176 99380 272196
rect 99380 272176 99432 272196
rect 99432 272176 99434 272196
rect 100758 271768 100814 271824
rect 106278 271768 106334 271824
rect 106554 271768 106610 271824
rect 112350 271768 112406 271824
rect 98090 271632 98146 271688
rect 107658 271632 107714 271688
rect 88338 271224 88394 271280
rect 88338 270816 88394 270872
rect 89718 270680 89774 270736
rect 92478 270680 92534 270736
rect 91098 270544 91154 270600
rect 85762 268368 85818 268424
rect 100758 271496 100814 271552
rect 104898 271360 104954 271416
rect 103518 271224 103574 271280
rect 109222 271360 109278 271416
rect 113270 271360 113326 271416
rect 104898 270680 104954 270736
rect 107658 270544 107714 270600
rect 110418 271224 110474 271280
rect 113178 271244 113234 271280
rect 113178 271224 113180 271244
rect 113180 271224 113232 271244
rect 113232 271224 113234 271244
rect 110418 270544 110474 270600
rect 133418 273672 133474 273728
rect 135902 273556 135958 273592
rect 135902 273536 135904 273556
rect 135904 273536 135956 273556
rect 135956 273536 135958 273556
rect 138478 273536 138534 273592
rect 140870 273536 140926 273592
rect 143538 273536 143594 273592
rect 145930 273536 145986 273592
rect 123114 271804 123116 271824
rect 123116 271804 123168 271824
rect 123168 271804 123170 271824
rect 123114 271768 123170 271804
rect 125598 271768 125654 271824
rect 128358 271788 128414 271824
rect 128358 271768 128360 271788
rect 128360 271768 128412 271788
rect 128412 271768 128414 271788
rect 151358 271788 151414 271824
rect 151358 271768 151360 271788
rect 151360 271768 151412 271788
rect 151412 271768 151414 271788
rect 154486 271804 154488 271824
rect 154488 271804 154540 271824
rect 154540 271804 154542 271824
rect 154486 271768 154542 271804
rect 157246 271768 157302 271824
rect 115938 271632 115994 271688
rect 117318 271632 117374 271688
rect 120078 271652 120134 271688
rect 120078 271632 120080 271652
rect 120080 271632 120132 271652
rect 120132 271632 120134 271652
rect 115846 271496 115902 271552
rect 158626 271652 158682 271688
rect 158626 271632 158628 271652
rect 158628 271632 158680 271652
rect 158680 271632 158682 271652
rect 161294 271632 161350 271688
rect 164146 271632 164202 271688
rect 183466 271360 183522 271416
rect 183466 271124 183468 271144
rect 183468 271124 183520 271144
rect 183520 271124 183522 271144
rect 183466 271088 183522 271124
rect 129738 270952 129794 271008
rect 147678 270680 147734 270736
rect 191746 253680 191802 253736
rect 179326 253172 179328 253192
rect 179328 253172 179380 253192
rect 179380 253172 179382 253192
rect 179326 253136 179382 253172
rect 180522 253136 180578 253192
rect 98458 166776 98514 166832
rect 101034 166776 101090 166832
rect 105818 166812 105820 166832
rect 105820 166812 105872 166832
rect 105872 166812 105874 166832
rect 105818 166776 105874 166812
rect 108210 166796 108266 166832
rect 108210 166776 108212 166796
rect 108212 166776 108264 166796
rect 108264 166776 108266 166796
rect 138478 166776 138534 166832
rect 140870 166776 140926 166832
rect 145930 166776 145986 166832
rect 163318 166640 163374 166696
rect 165894 166640 165950 166696
rect 114374 166504 114430 166560
rect 116950 166504 117006 166560
rect 148506 166524 148562 166560
rect 148506 166504 148508 166524
rect 148508 166504 148560 166524
rect 148560 166504 148562 166524
rect 96066 166252 96122 166288
rect 96066 166232 96068 166252
rect 96068 166232 96120 166252
rect 96120 166232 96122 166252
rect 153290 166504 153346 166560
rect 183282 166504 183338 166560
rect 81438 165552 81494 165608
rect 84198 165552 84254 165608
rect 89994 165552 90050 165608
rect 91098 165552 91154 165608
rect 95238 165552 95294 165608
rect 99378 165552 99434 165608
rect 103518 165552 103574 165608
rect 109498 165552 109554 165608
rect 110878 165552 110934 165608
rect 111154 165552 111210 165608
rect 113178 165552 113234 165608
rect 113546 165552 113602 165608
rect 115938 165552 115994 165608
rect 117962 165552 118018 165608
rect 118330 165552 118386 165608
rect 118974 165552 119030 165608
rect 120906 165552 120962 165608
rect 123482 165552 123538 165608
rect 125874 165552 125930 165608
rect 128358 165552 128414 165608
rect 129738 165552 129794 165608
rect 132498 165572 132554 165608
rect 132498 165552 132500 165572
rect 132500 165552 132552 165572
rect 132552 165552 132554 165572
rect 59910 165144 59966 165200
rect 76010 164328 76066 164384
rect 75918 164192 75974 164248
rect 59726 146104 59782 146160
rect 59358 140800 59414 140856
rect 77298 164192 77354 164248
rect 78678 164192 78734 164248
rect 80058 164192 80114 164248
rect 82818 164192 82874 164248
rect 88338 164872 88394 164928
rect 89902 164328 89958 164384
rect 84290 164192 84346 164248
rect 85578 164192 85634 164248
rect 86958 164192 87014 164248
rect 88430 164192 88486 164248
rect 91190 164192 91246 164248
rect 92478 164192 92534 164248
rect 93858 164192 93914 164248
rect 96618 164192 96674 164248
rect 97998 164192 98054 164248
rect 92478 145696 92534 145752
rect 107658 164872 107714 164928
rect 106278 164736 106334 164792
rect 100758 164484 100814 164520
rect 100758 164464 100760 164484
rect 100760 164464 100812 164484
rect 100812 164464 100814 164484
rect 100022 164192 100078 164248
rect 102138 164192 102194 164248
rect 103518 164192 103574 164248
rect 106186 164192 106242 164248
rect 106370 164192 106426 164248
rect 114558 164464 114614 164520
rect 115938 164464 115994 164520
rect 183374 165552 183430 165608
rect 200486 485288 200542 485344
rect 198830 400868 198832 400888
rect 198832 400868 198884 400888
rect 198884 400868 198886 400888
rect 198830 400832 198886 400868
rect 198830 351872 198886 351928
rect 198738 289720 198794 289776
rect 198738 288768 198794 288824
rect 100022 146240 100078 146296
rect 99378 146104 99434 146160
rect 98642 145560 98698 145616
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 191286 144880 191342 144936
rect 77114 59744 77170 59800
rect 83094 59744 83150 59800
rect 94502 59744 94558 59800
rect 101770 59744 101826 59800
rect 102782 59744 102838 59800
rect 113546 59744 113602 59800
rect 89994 59472 90050 59528
rect 95882 59472 95938 59528
rect 96986 59472 97042 59528
rect 98090 59472 98146 59528
rect 100758 59508 100760 59528
rect 100760 59508 100812 59528
rect 100812 59508 100814 59528
rect 100758 59472 100814 59508
rect 107566 59608 107622 59664
rect 110970 59336 111026 59392
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 84198 57976 84254 58032
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 78678 57840 78734 57896
rect 80426 57840 80482 57896
rect 81438 57840 81494 57896
rect 85394 57840 85450 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88338 57840 88394 57896
rect 88706 57840 88762 57896
rect 90730 57840 90786 57896
rect 91098 57840 91154 57896
rect 91466 57840 91522 57896
rect 93306 57840 93362 57896
rect 93674 57840 93730 57896
rect 99378 57840 99434 57896
rect 103794 57840 103850 57896
rect 106278 57840 106334 57896
rect 108210 57840 108266 57896
rect 109038 57840 109094 57896
rect 111154 57840 111210 57896
rect 112074 57840 112130 57896
rect 113178 57840 113234 57896
rect 115754 57840 115810 57896
rect 115938 57840 115994 57896
rect 119066 57840 119122 57896
rect 130842 57840 130898 57896
rect 133418 57840 133474 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 113270 57296 113326 57352
rect 115846 57568 115902 57624
rect 116122 57568 116178 57624
rect 115846 57296 115902 57352
rect 153290 57840 153346 57896
rect 183466 57860 183522 57896
rect 183466 57840 183468 57860
rect 183468 57840 183520 57860
rect 183520 57840 183522 57860
rect 122838 57568 122894 57624
rect 119066 56072 119122 56128
rect 199014 460128 199070 460184
rect 199474 398112 199530 398168
rect 199382 397296 199438 397352
rect 199290 394576 199346 394632
rect 199566 395256 199622 395312
rect 199014 353096 199070 353152
rect 199014 351872 199070 351928
rect 199290 292712 199346 292768
rect 199014 291624 199070 291680
rect 198830 246200 198886 246256
rect 198738 181872 198794 181928
rect 199198 290944 199254 291000
rect 199106 288360 199162 288416
rect 199106 287544 199162 287600
rect 198830 139168 198886 139224
rect 199014 184864 199070 184920
rect 199014 183504 199070 183560
rect 198922 77696 198978 77752
rect 199842 397296 199898 397352
rect 199566 292712 199622 292768
rect 199474 291624 199530 291680
rect 199382 289720 199438 289776
rect 199750 290944 199806 291000
rect 199658 288360 199714 288416
rect 201498 485188 201500 485208
rect 201500 485188 201552 485208
rect 201552 485188 201554 485208
rect 201498 485152 201554 485188
rect 202878 485016 202934 485072
rect 199290 186360 199346 186416
rect 199198 183504 199254 183560
rect 199198 180648 199254 180704
rect 199014 76336 199070 76392
rect 198738 74840 198794 74896
rect 202786 380704 202842 380760
rect 199290 79328 199346 79384
rect 199198 73616 199254 73672
rect 202970 380432 203026 380488
rect 202970 379208 203026 379264
rect 202970 378528 203026 378584
rect 204258 485152 204314 485208
rect 204258 484880 204314 484936
rect 203614 471144 203670 471200
rect 203706 465976 203762 466032
rect 205638 484744 205694 484800
rect 205178 380704 205234 380760
rect 205270 379208 205326 379264
rect 205362 379072 205418 379128
rect 205362 378392 205418 378448
rect 183190 57740 183192 57760
rect 183192 57740 183244 57760
rect 183244 57740 183246 57760
rect 183190 57704 183246 57740
rect 160098 57568 160154 57624
rect 162858 57568 162914 57624
rect 165618 57568 165674 57624
rect 153290 56208 153346 56264
rect 206190 378800 206246 378856
rect 206926 415248 206982 415304
rect 206190 270408 206246 270464
rect 206742 270408 206798 270464
rect 207018 379344 207074 379400
rect 207018 378528 207074 378584
rect 208214 378528 208270 378584
rect 208122 378256 208178 378312
rect 208122 269728 208178 269784
rect 208490 485288 208546 485344
rect 208398 380704 208454 380760
rect 208398 380296 208454 380352
rect 208398 379072 208454 379128
rect 208398 378664 208454 378720
rect 208306 378120 208362 378176
rect 208306 377984 208362 378040
rect 208858 379480 208914 379536
rect 209410 381520 209466 381576
rect 209686 380704 209742 380760
rect 209502 379072 209558 379128
rect 209410 270408 209466 270464
rect 209502 269864 209558 269920
rect 210238 378664 210294 378720
rect 211158 485288 211214 485344
rect 211158 484780 211160 484800
rect 211160 484780 211212 484800
rect 211212 484780 211214 484800
rect 211158 484744 211214 484780
rect 212538 485424 212594 485480
rect 210698 270952 210754 271008
rect 210974 269728 211030 269784
rect 211986 471280 212042 471336
rect 212078 271632 212134 271688
rect 212446 377984 212502 378040
rect 213182 271496 213238 271552
rect 213826 380432 213882 380488
rect 213642 271496 213698 271552
rect 213550 269864 213606 269920
rect 213274 145696 213330 145752
rect 165618 55120 165674 55176
rect 162858 54984 162914 55040
rect 160098 54848 160154 54904
rect 213826 377984 213882 378040
rect 214010 376216 214066 376272
rect 214470 376488 214526 376544
rect 214838 484472 214894 484528
rect 215206 377984 215262 378040
rect 215114 376624 215170 376680
rect 214470 145560 214526 145616
rect 214470 55120 214526 55176
rect 215482 377848 215538 377904
rect 215850 271768 215906 271824
rect 216034 465704 216090 465760
rect 216310 379208 216366 379264
rect 216218 271768 216274 271824
rect 216218 271224 216274 271280
rect 216678 417832 216734 417888
rect 216862 413752 216918 413808
rect 216678 410896 216734 410952
rect 216678 409148 216734 409184
rect 216678 409128 216680 409148
rect 216680 409128 216732 409148
rect 216732 409128 216734 409148
rect 216678 390904 216734 390960
rect 216678 389272 216734 389328
rect 216678 380840 216734 380896
rect 216678 380432 216734 380488
rect 217230 416880 217286 416936
rect 217138 414704 217194 414760
rect 216954 409128 217010 409184
rect 216954 380840 217010 380896
rect 217322 411984 217378 412040
rect 217322 411304 217378 411360
rect 217322 380840 217378 380896
rect 216954 380568 217010 380624
rect 217138 380568 217194 380624
rect 216586 375400 216642 375456
rect 215850 145968 215906 146024
rect 216862 309984 216918 310040
rect 216678 284008 216734 284064
rect 216678 282240 216734 282296
rect 216770 282104 216826 282160
rect 217046 309984 217102 310040
rect 216954 303864 217010 303920
rect 216954 302096 217010 302152
rect 216862 202952 216918 203008
rect 216862 198736 216918 198792
rect 217874 417832 217930 417888
rect 217782 411304 217838 411360
rect 217690 389000 217746 389056
rect 217598 380568 217654 380624
rect 217598 380024 217654 380080
rect 217598 307808 217654 307864
rect 217506 303864 217562 303920
rect 217322 302096 217378 302152
rect 216954 195200 217010 195256
rect 216770 176976 216826 177032
rect 216678 175344 216734 175400
rect 217046 175072 217102 175128
rect 217414 203904 217470 203960
rect 216862 92792 216918 92848
rect 216678 69944 216734 70000
rect 216678 68312 216734 68368
rect 217322 146240 217378 146296
rect 217782 380432 217838 380488
rect 217690 306720 217746 306776
rect 217598 200776 217654 200832
rect 217506 196968 217562 197024
rect 217414 96872 217470 96928
rect 218150 378528 218206 378584
rect 217966 377848 218022 377904
rect 217874 310936 217930 310992
rect 217782 304952 217838 305008
rect 217690 199824 217746 199880
rect 217690 198736 217746 198792
rect 218426 273400 218482 273456
rect 217966 252476 218022 252512
rect 217966 252456 217968 252476
rect 217968 252456 218020 252476
rect 218020 252456 218022 252476
rect 217874 203904 217930 203960
rect 217874 202952 217930 203008
rect 217782 198056 217838 198112
rect 217690 195200 217746 195256
rect 217598 93744 217654 93800
rect 217506 89936 217562 89992
rect 217966 162716 218022 162752
rect 217966 162696 217968 162716
rect 217968 162696 218020 162716
rect 218020 162696 218022 162716
rect 218242 146240 218298 146296
rect 217874 95920 217930 95976
rect 217782 91024 217838 91080
rect 217690 88168 217746 88224
rect 217966 68312 218022 68368
rect 218702 60560 218758 60616
rect 219622 270000 219678 270056
rect 219898 377848 219954 377904
rect 219438 145968 219494 146024
rect 219254 60560 219310 60616
rect 219898 146240 219954 146296
rect 219898 146104 219954 146160
rect 226154 485016 226210 485072
rect 224866 484472 224922 484528
rect 223670 479576 223726 479632
rect 223578 474000 223634 474056
rect 226338 472640 226394 472696
rect 228454 483792 228510 483848
rect 228546 478216 228602 478272
rect 231398 483656 231454 483712
rect 232318 485016 232374 485072
rect 232134 480800 232190 480856
rect 233238 485424 233294 485480
rect 234342 485152 234398 485208
rect 235814 485560 235870 485616
rect 235906 485288 235962 485344
rect 236550 482296 236606 482352
rect 234618 476720 234674 476776
rect 232410 475496 232466 475552
rect 229098 472504 229154 472560
rect 240322 478080 240378 478136
rect 252650 472912 252706 472968
rect 256238 482432 256294 482488
rect 270498 475632 270554 475688
rect 248418 465704 248474 465760
rect 286138 479712 286194 479768
rect 277398 465840 277454 465896
rect 295522 471144 295578 471200
rect 320822 639240 320878 639296
rect 321558 634480 321614 634536
rect 321558 629720 321614 629776
rect 321558 624960 321614 625016
rect 321558 620200 321614 620256
rect 321558 615440 321614 615496
rect 321558 610680 321614 610736
rect 321558 605920 321614 605976
rect 321558 596400 321614 596456
rect 321558 591640 321614 591696
rect 321558 586880 321614 586936
rect 321558 581440 321614 581496
rect 321006 576680 321062 576736
rect 321558 571920 321614 571976
rect 321558 567196 321560 567216
rect 321560 567196 321612 567216
rect 321612 567196 321614 567216
rect 321558 567160 321614 567196
rect 321558 562400 321614 562456
rect 321558 557640 321614 557696
rect 321558 552880 321614 552936
rect 322202 549888 322258 549944
rect 321558 548120 321614 548176
rect 321558 543360 321614 543416
rect 321558 538600 321614 538656
rect 322202 547984 322258 548040
rect 322110 533840 322166 533896
rect 321190 526904 321246 526960
rect 322202 526768 322258 526824
rect 324778 641688 324834 641744
rect 324226 601160 324282 601216
rect 323950 549752 324006 549808
rect 323950 528128 324006 528184
rect 423862 641688 423918 641744
rect 333058 639512 333114 639568
rect 433338 626184 433394 626240
rect 433338 615848 433394 615904
rect 324042 526632 324098 526688
rect 342718 526632 342774 526688
rect 360750 526768 360806 526824
rect 424506 527040 424562 527096
rect 429198 526904 429254 526960
rect 433430 601568 433486 601624
rect 433522 567432 433578 567488
rect 434626 529760 434682 529816
rect 434810 635160 434866 635216
rect 434810 592320 434866 592376
rect 397458 523640 397514 523696
rect 318062 482160 318118 482216
rect 296810 471280 296866 471336
rect 296718 468424 296774 468480
rect 338486 466556 338488 466576
rect 338488 466556 338540 466576
rect 338540 466556 338542 466576
rect 338486 466520 338542 466556
rect 339774 466540 339830 466576
rect 339774 466520 339776 466540
rect 339776 466520 339828 466540
rect 339828 466520 339830 466540
rect 350998 466520 351054 466576
rect 248234 380876 248236 380896
rect 248236 380876 248288 380896
rect 248288 380876 248290 380896
rect 248234 380840 248290 380876
rect 235998 380568 236054 380624
rect 237102 380568 237158 380624
rect 243082 380568 243138 380624
rect 245382 380568 245438 380624
rect 247590 380568 247646 380624
rect 254490 380568 254546 380624
rect 255870 380568 255926 380624
rect 256974 380568 257030 380624
rect 258078 380568 258134 380624
rect 259458 380568 259514 380624
rect 265254 380568 265310 380624
rect 265530 380568 265586 380624
rect 270958 380568 271014 380624
rect 246210 379344 246266 379400
rect 248602 379344 248658 379400
rect 250074 379344 250130 379400
rect 251178 379344 251234 379400
rect 252282 379344 252338 379400
rect 253386 379344 253442 379400
rect 261666 379344 261722 379400
rect 263874 379344 263930 379400
rect 253110 379072 253166 379128
rect 253110 378392 253166 378448
rect 244278 378256 244334 378312
rect 250626 378256 250682 378312
rect 239126 375944 239182 376000
rect 253570 378528 253626 378584
rect 255962 378528 256018 378584
rect 258354 378528 258410 378584
rect 260930 378528 260986 378584
rect 263598 378528 263654 378584
rect 262770 378256 262826 378312
rect 268658 379344 268714 379400
rect 265898 378528 265954 378584
rect 268106 378528 268162 378584
rect 265530 378392 265586 378448
rect 266358 378256 266414 378312
rect 267554 378256 267610 378312
rect 271050 379344 271106 379400
rect 272154 379344 272210 379400
rect 273258 379364 273314 379400
rect 273258 379344 273260 379364
rect 273260 379344 273312 379364
rect 273312 379344 273314 379364
rect 274362 379380 274364 379400
rect 274364 379380 274416 379400
rect 274416 379380 274418 379400
rect 274362 379344 274418 379380
rect 275650 379344 275706 379400
rect 276110 379344 276166 379400
rect 277030 379344 277086 379400
rect 278226 379344 278282 379400
rect 285954 379344 286010 379400
rect 287610 379344 287666 379400
rect 290922 379344 290978 379400
rect 292670 379344 292726 379400
rect 273442 378528 273498 378584
rect 276018 378120 276074 378176
rect 280250 379208 280306 379264
rect 283378 379208 283434 379264
rect 295430 379344 295486 379400
rect 298466 379344 298522 379400
rect 300858 379344 300914 379400
rect 303250 379344 303306 379400
rect 305826 379344 305882 379400
rect 307850 379344 307906 379400
rect 310978 379364 311034 379400
rect 310978 379344 310980 379364
rect 310980 379344 311032 379364
rect 311032 379344 311034 379364
rect 313370 379344 313426 379400
rect 315762 379380 315764 379400
rect 315764 379380 315816 379400
rect 315816 379380 315818 379400
rect 315762 379344 315818 379380
rect 317418 379344 317474 379400
rect 325882 379208 325938 379264
rect 320914 378528 320970 378584
rect 343178 378392 343234 378448
rect 343546 378256 343602 378312
rect 338486 358808 338542 358864
rect 340050 358808 340106 358864
rect 351734 358808 351790 358864
rect 266358 273536 266414 273592
rect 283470 273536 283526 273592
rect 273258 273400 273314 273456
rect 285954 272856 286010 272912
rect 288162 272856 288218 272912
rect 290922 272876 290978 272912
rect 290922 272856 290924 272876
rect 290924 272856 290976 272876
rect 290976 272856 290978 272876
rect 295890 272892 295892 272912
rect 295892 272892 295944 272912
rect 295944 272892 295946 272912
rect 295890 272856 295946 272892
rect 303434 272856 303490 272912
rect 298466 272740 298522 272776
rect 298466 272720 298468 272740
rect 298468 272720 298520 272740
rect 298520 272720 298522 272740
rect 300858 272720 300914 272776
rect 305826 272604 305882 272640
rect 305826 272584 305828 272604
rect 305828 272584 305880 272604
rect 305880 272584 305882 272604
rect 320914 272584 320970 272640
rect 265162 272176 265218 272232
rect 263598 271768 263654 271824
rect 264978 271768 265034 271824
rect 258262 271224 258318 271280
rect 260838 271244 260894 271280
rect 260838 271224 260840 271244
rect 260840 271224 260892 271244
rect 260892 271224 260894 271244
rect 247038 271088 247094 271144
rect 252558 271108 252614 271144
rect 252558 271088 252560 271108
rect 252560 271088 252612 271108
rect 252612 271088 252614 271108
rect 255318 271088 255374 271144
rect 253938 270816 253994 270872
rect 244370 270680 244426 270736
rect 251270 270680 251326 270736
rect 237378 270544 237434 270600
rect 242898 270544 242954 270600
rect 244278 270544 244334 270600
rect 220726 270000 220782 270056
rect 245658 270544 245714 270600
rect 247038 270544 247094 270600
rect 248510 270544 248566 270600
rect 249798 270544 249854 270600
rect 251178 270544 251234 270600
rect 252558 270544 252614 270600
rect 255318 270680 255374 270736
rect 259550 270680 259606 270736
rect 256698 270544 256754 270600
rect 258078 270544 258134 270600
rect 259458 270544 259514 270600
rect 260838 270544 260894 270600
rect 262218 270544 262274 270600
rect 263598 270544 263654 270600
rect 268014 271768 268070 271824
rect 270498 271768 270554 271824
rect 271878 271768 271934 271824
rect 276018 271768 276074 271824
rect 277950 271768 278006 271824
rect 280066 271768 280122 271824
rect 280250 271768 280306 271824
rect 307758 271788 307814 271824
rect 307758 271768 307760 271788
rect 307760 271768 307812 271788
rect 307812 271768 307814 271788
rect 270498 271224 270554 271280
rect 267922 270816 267978 270872
rect 266358 270544 266414 270600
rect 269118 270544 269174 270600
rect 277214 271496 277270 271552
rect 313278 271804 313280 271824
rect 313280 271804 313332 271824
rect 313332 271804 313334 271824
rect 313278 271768 313334 271804
rect 343546 271496 343602 271552
rect 343454 271360 343510 271416
rect 277398 270816 277454 270872
rect 273166 270544 273222 270600
rect 274638 270544 274694 270600
rect 339406 253544 339462 253600
rect 351826 253172 351828 253192
rect 351828 253172 351880 253192
rect 351880 253172 351882 253192
rect 351826 253136 351882 253172
rect 340786 253000 340842 253056
rect 303526 166640 303582 166696
rect 285954 166524 286010 166560
rect 285954 166504 285956 166524
rect 285956 166504 286008 166524
rect 286008 166504 286010 166524
rect 288254 166504 288310 166560
rect 293406 166540 293408 166560
rect 293408 166540 293460 166560
rect 293460 166540 293462 166560
rect 293406 166504 293462 166540
rect 295890 166504 295946 166560
rect 260930 166368 260986 166424
rect 265898 166368 265954 166424
rect 235998 165552 236054 165608
rect 238758 165552 238814 165608
rect 242898 165552 242954 165608
rect 247038 165552 247094 165608
rect 247682 165552 247738 165608
rect 249798 165552 249854 165608
rect 252558 165552 252614 165608
rect 258078 165552 258134 165608
rect 260838 165552 260894 165608
rect 264978 165552 265034 165608
rect 267738 165552 267794 165608
rect 271878 165552 271934 165608
rect 273442 165552 273498 165608
rect 275926 165552 275982 165608
rect 236090 164192 236146 164248
rect 237378 164192 237434 164248
rect 220818 146104 220874 146160
rect 240138 164192 240194 164248
rect 241518 164192 241574 164248
rect 244370 164464 244426 164520
rect 244278 164192 244334 164248
rect 237378 145696 237434 145752
rect 245658 164192 245714 164248
rect 251270 164464 251326 164520
rect 259550 164464 259606 164520
rect 248418 164192 248474 164248
rect 249798 164192 249854 164248
rect 251178 164192 251234 164248
rect 252558 164192 252614 164248
rect 253938 164192 253994 164248
rect 255318 164192 255374 164248
rect 256698 164192 256754 164248
rect 258078 164192 258134 164248
rect 259458 164192 259514 164248
rect 263506 164192 263562 164248
rect 263782 164192 263838 164248
rect 266358 164600 266414 164656
rect 267646 164464 267702 164520
rect 267830 164192 267886 164248
rect 269118 164192 269174 164248
rect 270498 164192 270554 164248
rect 267738 146240 267794 146296
rect 267830 146104 267886 146160
rect 263598 145968 263654 146024
rect 274454 164464 274510 164520
rect 274546 164192 274602 164248
rect 276018 164192 276074 164248
rect 276202 165552 276258 165608
rect 277398 165552 277454 165608
rect 280066 165552 280122 165608
rect 280250 165552 280306 165608
rect 283378 165552 283434 165608
rect 300858 165572 300914 165608
rect 300858 165552 300860 165572
rect 300860 165552 300912 165572
rect 300912 165552 300914 165572
rect 277398 164192 277454 164248
rect 323306 165552 323362 165608
rect 343454 165552 343510 165608
rect 343546 165416 343602 165472
rect 269118 145560 269174 145616
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 237102 59744 237158 59800
rect 255870 59744 255926 59800
rect 256974 59744 257030 59800
rect 262862 59744 262918 59800
rect 263874 59744 263930 59800
rect 258078 59608 258134 59664
rect 260654 59608 260710 59664
rect 261758 59608 261814 59664
rect 308494 59608 308550 59664
rect 315854 59608 315910 59664
rect 279238 59336 279294 59392
rect 290922 59200 290978 59256
rect 300858 59200 300914 59256
rect 320914 59200 320970 59256
rect 325882 59200 325938 59256
rect 357438 380160 357494 380216
rect 235998 57840 236054 57896
rect 237378 57840 237434 57896
rect 239218 57840 239274 57896
rect 240138 57840 240194 57896
rect 241610 57840 241666 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 245290 57840 245346 57896
rect 245658 57840 245714 57896
rect 247038 57840 247094 57896
rect 248234 57840 248290 57896
rect 248602 57840 248658 57896
rect 249798 57840 249854 57896
rect 251178 57840 251234 57896
rect 251362 57840 251418 57896
rect 253386 57840 253442 57896
rect 253938 57840 253994 57896
rect 258354 57840 258410 57896
rect 264978 57840 265034 57896
rect 266450 57840 266506 57896
rect 268106 57840 268162 57896
rect 268934 57840 268990 57896
rect 271050 57840 271106 57896
rect 271878 57840 271934 57896
rect 273258 57840 273314 57896
rect 275098 57840 275154 57896
rect 276938 57840 276994 57896
rect 278318 57840 278374 57896
rect 295890 57840 295946 57896
rect 298098 57840 298154 57896
rect 303434 57840 303490 57896
rect 305826 57840 305882 57896
rect 310978 57840 311034 57896
rect 313370 57860 313426 57896
rect 313370 57840 313372 57860
rect 313372 57840 313424 57860
rect 313424 57840 313426 57860
rect 266358 57296 266414 57352
rect 268934 57568 268990 57624
rect 269118 57568 269174 57624
rect 269118 55120 269174 55176
rect 273350 57568 273406 57624
rect 277398 57568 277454 57624
rect 318246 57840 318302 57896
rect 323306 57876 323308 57896
rect 323308 57876 323360 57896
rect 323360 57876 323362 57896
rect 323306 57840 323362 57876
rect 343178 57876 343180 57896
rect 343180 57876 343232 57896
rect 343232 57876 343234 57896
rect 343178 57840 343234 57876
rect 343454 57860 343510 57896
rect 358910 460128 358966 460184
rect 359002 400288 359058 400344
rect 359094 398112 359150 398168
rect 359186 395256 359242 395312
rect 359278 394032 359334 394088
rect 359738 396752 359794 396808
rect 358910 353096 358966 353152
rect 359094 291760 359150 291816
rect 359002 290944 359058 291000
rect 359002 289720 359058 289776
rect 359002 288768 359058 288824
rect 358910 246200 358966 246256
rect 358818 186360 358874 186416
rect 359278 292712 359334 292768
rect 359186 287544 359242 287600
rect 359094 184864 359150 184920
rect 359002 182008 359058 182064
rect 358910 139304 358966 139360
rect 358818 79872 358874 79928
rect 359370 290944 359426 291000
rect 359278 186360 359334 186416
rect 359554 292712 359610 292768
rect 359646 291760 359702 291816
rect 359462 289720 359518 289776
rect 359370 183368 359426 183424
rect 359278 182008 359334 182064
rect 359186 180648 359242 180704
rect 359094 78240 359150 78296
rect 359370 76880 359426 76936
rect 359278 75384 359334 75440
rect 359186 74024 359242 74080
rect 361486 377984 361542 378040
rect 343454 57840 343456 57860
rect 343456 57840 343508 57860
rect 343508 57840 343510 57860
rect 363510 377984 363566 378040
rect 370962 379072 371018 379128
rect 370870 378936 370926 378992
rect 371146 377848 371202 377904
rect 369766 145832 369822 145888
rect 371054 145696 371110 145752
rect 371790 380160 371846 380216
rect 371698 273264 371754 273320
rect 371698 145560 371754 145616
rect 372710 378800 372766 378856
rect 372526 270000 372582 270056
rect 372986 269184 373042 269240
rect 373538 270952 373594 271008
rect 375102 378664 375158 378720
rect 375286 378700 375288 378720
rect 375288 378700 375340 378720
rect 375340 378700 375342 378720
rect 375286 378664 375342 378700
rect 374918 269864 374974 269920
rect 375746 270544 375802 270600
rect 375562 164056 375618 164112
rect 375838 269320 375894 269376
rect 376390 271496 376446 271552
rect 376574 271224 376630 271280
rect 376574 270544 376630 270600
rect 376482 270272 376538 270328
rect 376390 270000 376446 270056
rect 376298 165552 376354 165608
rect 377218 416880 377274 416936
rect 376942 415248 376998 415304
rect 376942 414704 376998 414760
rect 377218 411984 377274 412040
rect 377218 410896 377274 410952
rect 376942 390904 376998 390960
rect 376942 389272 376998 389328
rect 376942 389000 376998 389056
rect 376758 374856 376814 374912
rect 377402 415248 377458 415304
rect 377402 409148 377458 409184
rect 377402 409128 377404 409148
rect 377404 409128 377456 409148
rect 377456 409128 377458 409148
rect 377402 378120 377458 378176
rect 377770 417832 377826 417888
rect 377586 413888 377642 413944
rect 377586 411984 377642 412040
rect 376850 307808 376906 307864
rect 376942 307672 376998 307728
rect 376850 284008 376906 284064
rect 376942 282240 376998 282296
rect 376482 269864 376538 269920
rect 376114 164600 376170 164656
rect 376022 68040 376078 68096
rect 376758 269320 376814 269376
rect 376850 201320 376906 201376
rect 377402 310800 377458 310856
rect 377218 309984 377274 310040
rect 377310 302096 377366 302152
rect 377218 203904 377274 203960
rect 377034 202952 377090 203008
rect 376942 199824 376998 199880
rect 376942 176976 376998 177032
rect 376942 175344 376998 175400
rect 376942 175072 376998 175128
rect 377954 416880 378010 416936
rect 377862 413888 377918 413944
rect 377770 310800 377826 310856
rect 378046 409128 378102 409184
rect 377954 309984 378010 310040
rect 377862 307672 377918 307728
rect 377862 306856 377918 306912
rect 377586 304952 377642 305008
rect 377862 303864 377918 303920
rect 377586 282104 377642 282160
rect 377678 267552 377734 267608
rect 377678 252492 377680 252512
rect 377680 252492 377732 252512
rect 377732 252492 377734 252512
rect 377678 252456 377734 252492
rect 377402 203904 377458 203960
rect 377586 201320 377642 201376
rect 377586 200776 377642 200832
rect 377310 195200 377366 195256
rect 377218 96872 377274 96928
rect 377034 95920 377090 95976
rect 376942 92792 376998 92848
rect 376942 69944 376998 70000
rect 376666 68856 376722 68912
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 377494 145696 377550 145752
rect 377678 198056 377734 198112
rect 377586 93744 377642 93800
rect 378046 302096 378102 302152
rect 378506 273264 378562 273320
rect 377862 196968 377918 197024
rect 377770 195200 377826 195256
rect 377678 91024 377734 91080
rect 377862 89936 377918 89992
rect 377770 88168 377826 88224
rect 378690 269184 378746 269240
rect 378782 165280 378838 165336
rect 436190 630400 436246 630456
rect 436098 620880 436154 620936
rect 580170 683848 580226 683904
rect 477130 634888 477186 634944
rect 488722 634888 488778 634944
rect 506754 634888 506810 634944
rect 457810 634752 457866 634808
rect 457718 629176 457774 629232
rect 457626 623056 457682 623112
rect 512182 631896 512238 631952
rect 512090 626456 512146 626512
rect 511998 619520 512054 619576
rect 457534 616800 457590 616856
rect 511998 612720 512054 612776
rect 457626 608912 457682 608968
rect 457534 603064 457590 603120
rect 457442 597488 457498 597544
rect 436098 597080 436154 597136
rect 434902 539280 434958 539336
rect 457442 590688 457498 590744
rect 436190 582120 436246 582176
rect 436282 577360 436338 577416
rect 436374 572600 436430 572656
rect 436466 563080 436522 563136
rect 436558 558320 436614 558376
rect 436650 553560 436706 553616
rect 436742 548800 436798 548856
rect 436834 544040 436890 544096
rect 436926 534520 436982 534576
rect 457534 486512 457590 486568
rect 500958 529488 501014 529544
rect 506478 518064 506534 518120
rect 512182 606328 512238 606384
rect 512090 600344 512146 600400
rect 511998 487736 512054 487792
rect 512274 593952 512330 594008
rect 513286 586508 513288 586528
rect 513288 586508 513340 586528
rect 513340 586508 513342 586528
rect 513286 586472 513342 586508
rect 512090 479440 512146 479496
rect 483018 475360 483074 475416
rect 379702 382336 379758 382392
rect 379150 271768 379206 271824
rect 379518 357312 379574 357368
rect 379426 270408 379482 270464
rect 378966 165416 379022 165472
rect 378874 146240 378930 146296
rect 378874 145968 378930 146024
rect 379058 147736 379114 147792
rect 498474 466556 498476 466576
rect 498476 466556 498528 466576
rect 498528 466556 498530 466576
rect 498474 466520 498530 466556
rect 499762 466540 499818 466576
rect 499762 466520 499764 466540
rect 499764 466520 499816 466540
rect 499816 466520 499818 466540
rect 510894 466540 510950 466576
rect 510894 466520 510896 466540
rect 510896 466520 510948 466540
rect 510948 466520 510950 466540
rect 431130 380876 431132 380896
rect 431132 380876 431184 380896
rect 431184 380876 431186 380896
rect 431130 380840 431186 380876
rect 433614 380840 433670 380896
rect 438490 380840 438546 380896
rect 410706 380704 410762 380760
rect 421102 380704 421158 380760
rect 405462 380568 405518 380624
rect 413466 380568 413522 380624
rect 419446 380568 419502 380624
rect 379794 271088 379850 271144
rect 379794 270408 379850 270464
rect 381266 378800 381322 378856
rect 381082 378664 381138 378720
rect 379794 269728 379850 269784
rect 436006 380704 436062 380760
rect 434350 380568 434406 380624
rect 426438 380432 426494 380488
rect 440882 380704 440938 380760
rect 443458 380704 443514 380760
rect 485962 380568 486018 380624
rect 396078 379344 396134 379400
rect 397090 379344 397146 379400
rect 405830 379344 405886 379400
rect 407578 379344 407634 379400
rect 408314 379344 408370 379400
rect 411258 379344 411314 379400
rect 412362 379344 412418 379400
rect 415674 379344 415730 379400
rect 425978 379344 426034 379400
rect 435178 379344 435234 379400
rect 437846 379344 437902 379400
rect 445850 379344 445906 379400
rect 447506 379344 447562 379400
rect 451002 379344 451058 379400
rect 453026 379344 453082 379400
rect 455510 379344 455566 379400
rect 458362 379344 458418 379400
rect 460938 379344 460994 379400
rect 474830 379344 474886 379400
rect 399482 379208 399538 379264
rect 400402 379208 400458 379264
rect 402978 379208 403034 379264
rect 409970 379208 410026 379264
rect 408682 378120 408738 378176
rect 413282 378528 413338 378584
rect 414570 378528 414626 378584
rect 415858 379208 415914 379264
rect 416870 379208 416926 379264
rect 422850 379208 422906 379264
rect 418434 378528 418490 378584
rect 418158 378120 418214 378176
rect 420642 378120 420698 378176
rect 421194 378120 421250 378176
rect 422666 378120 422722 378176
rect 423954 378120 424010 378176
rect 425150 378120 425206 378176
rect 430670 378800 430726 378856
rect 428554 378120 428610 378176
rect 429658 378120 429714 378176
rect 436190 378664 436246 378720
rect 432234 378256 432290 378312
rect 439042 378120 439098 378176
rect 463514 379208 463570 379264
rect 473450 379208 473506 379264
rect 465170 378936 465226 378992
rect 470782 378800 470838 378856
rect 467930 378664 467986 378720
rect 465170 376624 465226 376680
rect 503074 379208 503130 379264
rect 503534 379208 503590 379264
rect 477590 378936 477646 378992
rect 483386 378800 483442 378856
rect 498934 358808 498990 358864
rect 500406 358808 500462 358864
rect 510894 358828 510950 358864
rect 510894 358808 510896 358828
rect 510896 358808 510948 358828
rect 510948 358808 510950 358828
rect 426438 273808 426494 273864
rect 421102 273556 421158 273592
rect 421102 273536 421104 273556
rect 421104 273536 421156 273556
rect 421156 273536 421158 273556
rect 431130 273536 431186 273592
rect 433338 273536 433394 273592
rect 453394 273536 453450 273592
rect 430946 273400 431002 273456
rect 422666 273128 422722 273184
rect 422850 273164 422852 273184
rect 422852 273164 422904 273184
rect 422904 273164 422906 273184
rect 422850 273128 422906 273164
rect 423402 273128 423458 273184
rect 425978 273148 426034 273184
rect 425978 273128 425980 273148
rect 425980 273128 426032 273148
rect 426032 273128 426034 273148
rect 468482 273012 468538 273048
rect 468482 272992 468484 273012
rect 468484 272992 468536 273012
rect 468536 272992 468538 273012
rect 470874 272992 470930 273048
rect 422666 272856 422722 272912
rect 473450 272876 473506 272912
rect 473450 272856 473452 272876
rect 473452 272856 473504 272876
rect 473504 272856 473506 272876
rect 475842 272856 475898 272912
rect 478418 272740 478474 272776
rect 478418 272720 478420 272740
rect 478420 272720 478472 272740
rect 478472 272720 478474 272740
rect 480810 272720 480866 272776
rect 380070 272584 380126 272640
rect 483202 272604 483258 272640
rect 483202 272584 483204 272604
rect 483204 272584 483256 272604
rect 483256 272584 483258 272604
rect 485962 272584 486018 272640
rect 423770 272468 423826 272504
rect 423770 272448 423772 272468
rect 423772 272448 423824 272468
rect 423824 272448 423826 272468
rect 401690 272176 401746 272232
rect 415858 272176 415914 272232
rect 416042 272176 416098 272232
rect 455786 272176 455842 272232
rect 380162 271088 380218 271144
rect 387890 269320 387946 269376
rect 390558 269184 390614 269240
rect 397458 270544 397514 270600
rect 398838 270544 398894 270600
rect 400218 270544 400274 270600
rect 409878 271088 409934 271144
rect 412730 271088 412786 271144
rect 418158 271108 418214 271144
rect 418158 271088 418160 271108
rect 418160 271088 418212 271108
rect 418212 271088 418214 271108
rect 405738 270816 405794 270872
rect 402978 270544 403034 270600
rect 403346 270544 403402 270600
rect 404358 270544 404414 270600
rect 411350 270680 411406 270736
rect 407118 270544 407174 270600
rect 408498 270544 408554 270600
rect 409878 270544 409934 270600
rect 411258 270544 411314 270600
rect 413006 270544 413062 270600
rect 414018 270544 414074 270600
rect 416778 270544 416834 270600
rect 418158 270544 418214 270600
rect 419538 270544 419594 270600
rect 420918 270544 420974 270600
rect 427818 271768 427874 271824
rect 433338 271768 433394 271824
rect 436098 271768 436154 271824
rect 437478 271768 437534 271824
rect 442998 271768 443054 271824
rect 445758 271768 445814 271824
rect 447138 271768 447194 271824
rect 449898 271768 449954 271824
rect 458178 271788 458234 271824
rect 458178 271768 458180 271788
rect 458180 271768 458232 271788
rect 458232 271768 458234 271788
rect 503626 271632 503682 271688
rect 440238 271360 440294 271416
rect 434718 271244 434774 271280
rect 434718 271224 434720 271244
rect 434720 271224 434772 271244
rect 434772 271224 434774 271244
rect 503534 271224 503590 271280
rect 431958 270816 432014 270872
rect 433338 270816 433394 270872
rect 437478 270816 437534 270872
rect 438858 270816 438914 270872
rect 429198 270680 429254 270736
rect 500866 253308 500868 253328
rect 500868 253308 500920 253328
rect 500920 253308 500922 253328
rect 500866 253272 500922 253308
rect 499210 252728 499266 252784
rect 510894 252612 510950 252648
rect 580354 630808 580410 630864
rect 580262 577632 580318 577688
rect 580170 511264 580226 511320
rect 518898 459584 518954 459640
rect 519450 459584 519506 459640
rect 519082 400288 519138 400344
rect 518990 398112 519046 398168
rect 519358 396752 519414 396808
rect 519174 395256 519230 395312
rect 519266 394032 519322 394088
rect 510894 252592 510896 252612
rect 510896 252592 510948 252612
rect 510948 252592 510950 252612
rect 418434 166812 418436 166832
rect 418436 166812 418488 166832
rect 418488 166812 418490 166832
rect 418434 166776 418490 166812
rect 421010 166776 421066 166832
rect 423402 166776 423458 166832
rect 428186 166796 428242 166832
rect 428186 166776 428188 166796
rect 428188 166776 428240 166796
rect 428240 166776 428242 166796
rect 445850 166776 445906 166832
rect 470966 166776 471022 166832
rect 475842 166776 475898 166832
rect 478418 166776 478474 166832
rect 480902 166776 480958 166832
rect 483386 166640 483442 166696
rect 485962 166640 486018 166696
rect 503258 166504 503314 166560
rect 380530 165552 380586 165608
rect 397458 165552 397514 165608
rect 401598 165552 401654 165608
rect 404358 165552 404414 165608
rect 409878 165552 409934 165608
rect 415490 165552 415546 165608
rect 416042 165552 416098 165608
rect 418526 165552 418582 165608
rect 423770 165552 423826 165608
rect 433430 165552 433486 165608
rect 434718 165552 434774 165608
rect 436098 165588 436100 165608
rect 436100 165588 436152 165608
rect 436152 165588 436154 165608
rect 436098 165552 436154 165588
rect 437754 165552 437810 165608
rect 438030 165552 438086 165608
rect 440146 165552 440202 165608
rect 380530 165280 380586 165336
rect 396170 164328 396226 164384
rect 396078 164192 396134 164248
rect 398838 164192 398894 164248
rect 400218 164192 400274 164248
rect 402978 164328 403034 164384
rect 403070 164192 403126 164248
rect 407118 164872 407174 164928
rect 412638 164756 412694 164792
rect 412638 164736 412640 164756
rect 412640 164736 412692 164756
rect 412692 164736 412694 164756
rect 411258 164328 411314 164384
rect 405738 164192 405794 164248
rect 407210 164192 407266 164248
rect 408498 164192 408554 164248
rect 409878 164192 409934 164248
rect 411350 164192 411406 164248
rect 412730 164192 412786 164248
rect 414018 164192 414074 164248
rect 416778 164192 416834 164248
rect 418158 164192 418214 164248
rect 420918 164736 420974 164792
rect 419538 164192 419594 164248
rect 423586 164192 423642 164248
rect 415490 145968 415546 146024
rect 423678 145832 423734 145888
rect 433338 164892 433394 164928
rect 433338 164872 433340 164892
rect 433340 164872 433392 164892
rect 433392 164872 433394 164892
rect 426530 164328 426586 164384
rect 426346 164192 426402 164248
rect 423770 145696 423826 145752
rect 427726 164192 427782 164248
rect 430670 164736 430726 164792
rect 429290 164328 429346 164384
rect 429106 164192 429162 164248
rect 430578 164212 430634 164248
rect 430578 164192 430580 164212
rect 430580 164192 430632 164212
rect 430632 164192 430634 164212
rect 431958 164192 432014 164248
rect 434626 164192 434682 164248
rect 434810 164192 434866 164248
rect 437754 162696 437810 162752
rect 442998 165552 443054 165608
rect 447322 165552 447378 165608
rect 449898 165552 449954 165608
rect 452658 165552 452714 165608
rect 455418 165572 455474 165608
rect 455418 165552 455420 165572
rect 455420 165552 455472 165572
rect 455472 165552 455474 165572
rect 458362 165552 458418 165608
rect 503350 165552 503406 165608
rect 440330 165028 440386 165064
rect 440330 165008 440332 165028
rect 440332 165008 440384 165028
rect 440384 165008 440386 165028
rect 426438 145560 426494 145616
rect 510618 145424 510674 145480
rect 498658 144880 498714 144936
rect 500222 144880 500278 144936
rect 396078 59744 396134 59800
rect 397090 59744 397146 59800
rect 416962 59744 417018 59800
rect 423494 59744 423550 59800
rect 423954 59744 424010 59800
rect 403070 59608 403126 59664
rect 404174 59608 404230 59664
rect 412546 59608 412602 59664
rect 416042 59608 416098 59664
rect 410706 59472 410762 59528
rect 397458 57840 397514 57896
rect 399482 57840 399538 57896
rect 400218 57840 400274 57896
rect 401690 57840 401746 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407210 57840 407266 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 411258 56888 411314 56944
rect 419446 59608 419502 59664
rect 421746 59608 421802 59664
rect 418158 59472 418214 59528
rect 420642 59472 420698 59528
rect 458454 59608 458510 59664
rect 503258 59608 503314 59664
rect 425978 59336 426034 59392
rect 428186 59336 428242 59392
rect 453394 59336 453450 59392
rect 475842 58928 475898 58984
rect 414570 57840 414626 57896
rect 415490 57840 415546 57896
rect 426530 57840 426586 57896
rect 427634 57840 427690 57896
rect 427818 57840 427874 57896
rect 429198 57840 429254 57896
rect 430578 57840 430634 57896
rect 432234 57840 432290 57896
rect 434442 57840 434498 57896
rect 435914 57840 435970 57896
rect 436282 57840 436338 57896
rect 438490 57840 438546 57896
rect 445850 57840 445906 57896
rect 451002 57840 451058 57896
rect 460938 57840 460994 57896
rect 465906 57840 465962 57896
rect 470874 57860 470930 57896
rect 470874 57840 470876 57860
rect 470876 57840 470928 57860
rect 470928 57840 470930 57860
rect 412546 56888 412602 56944
rect 412638 56752 412694 56808
rect 430946 57160 431002 57216
rect 433154 57568 433210 57624
rect 433430 57568 433486 57624
rect 433154 57160 433210 57216
rect 434718 57568 434774 57624
rect 437478 57568 437534 57624
rect 478418 57840 478474 57896
rect 485962 57876 485964 57896
rect 485964 57876 486016 57896
rect 486016 57876 486018 57896
rect 485962 57840 486018 57876
rect 518898 292440 518954 292496
rect 519266 352824 519322 352880
rect 519174 288768 519230 288824
rect 518990 287544 519046 287600
rect 518898 186360 518954 186416
rect 503350 57876 503352 57896
rect 503352 57876 503404 57896
rect 503404 57876 503406 57896
rect 503350 57840 503406 57876
rect 518990 180648 519046 180704
rect 518898 79872 518954 79928
rect 580262 458088 580318 458144
rect 580354 404912 580410 404968
rect 580170 378392 580226 378448
rect 519450 352824 519506 352880
rect 519358 293800 519414 293856
rect 519266 246200 519322 246256
rect 519174 181872 519230 181928
rect 580354 351872 580410 351928
rect 580262 325216 580318 325272
rect 519634 292440 519690 292496
rect 519542 290264 519598 290320
rect 519358 186360 519414 186416
rect 520186 288768 520242 288824
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 519634 184728 519690 184784
rect 520186 184728 520242 184784
rect 519450 183368 519506 183424
rect 520094 183368 520150 183424
rect 519358 181872 519414 181928
rect 519266 139304 519322 139360
rect 519082 78240 519138 78296
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519450 76744 519506 76800
rect 519358 75384 519414 75440
rect 518990 74160 519046 74216
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
rect 140042 3984 140098 4040
rect 129370 3848 129426 3904
rect 136454 3440 136510 3496
rect 132958 3304 133014 3360
rect 147126 3712 147182 3768
rect 143538 3168 143594 3224
rect 150622 3576 150678 3632
rect 365718 3168 365774 3224
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 324773 641746 324839 641749
rect 423857 641746 423923 641749
rect 324773 641744 423923 641746
rect 324773 641688 324778 641744
rect 324834 641688 423862 641744
rect 423918 641688 423923 641744
rect 324773 641686 423923 641688
rect 324773 641683 324839 641686
rect 423857 641683 423923 641686
rect 333053 639570 333119 639573
rect 315990 639568 333119 639570
rect 315990 639512 333058 639568
rect 333114 639512 333119 639568
rect 315990 639510 333119 639512
rect 54334 639372 54340 639436
rect 54404 639434 54410 639436
rect 315990 639434 316050 639510
rect 333053 639507 333119 639510
rect 54404 639374 316050 639434
rect 54404 639372 54410 639374
rect 320817 639298 320883 639301
rect 320817 639296 325036 639298
rect 320817 639240 320822 639296
rect 320878 639240 325036 639296
rect 320817 639238 325036 639240
rect 320817 639235 320883 639238
rect 238710 635838 240426 635898
rect 237373 635762 237439 635765
rect 238710 635762 238770 635838
rect 237373 635760 238770 635762
rect 237373 635704 237378 635760
rect 237434 635704 238770 635760
rect 237373 635702 238770 635704
rect 237373 635699 237439 635702
rect 57605 635626 57671 635629
rect 147121 635626 147187 635629
rect 57605 635624 60076 635626
rect 57605 635568 57610 635624
rect 57666 635568 60076 635624
rect 57605 635566 60076 635568
rect 147121 635624 150052 635626
rect 147121 635568 147126 635624
rect 147182 635568 150052 635624
rect 240366 635596 240426 635838
rect 147121 635566 150052 635568
rect 57605 635563 57671 635566
rect 147121 635563 147187 635566
rect 211153 635218 211219 635221
rect 300853 635218 300919 635221
rect 434805 635218 434871 635221
rect 210558 635216 211219 635218
rect 210558 635160 211158 635216
rect 211214 635160 211219 635216
rect 210558 635158 211219 635160
rect 122925 634946 122991 634949
rect 120796 634944 122991 634946
rect 120796 634888 122930 634944
rect 122986 634888 122991 634944
rect 210558 634916 210618 635158
rect 211153 635155 211219 635158
rect 300718 635216 300919 635218
rect 300718 635160 300858 635216
rect 300914 635160 300919 635216
rect 300718 635158 300919 635160
rect 433780 635216 434871 635218
rect 433780 635160 434810 635216
rect 434866 635160 434871 635216
rect 433780 635158 434871 635160
rect 300718 634916 300778 635158
rect 300853 635155 300919 635158
rect 434805 635155 434871 635158
rect 120796 634886 122991 634888
rect 122925 634883 122991 634886
rect 476062 634884 476068 634948
rect 476132 634946 476138 634948
rect 477125 634946 477191 634949
rect 476132 634944 477191 634946
rect 476132 634888 477130 634944
rect 477186 634888 477191 634944
rect 476132 634886 477191 634888
rect 476132 634884 476138 634886
rect 477125 634883 477191 634886
rect 488574 634884 488580 634948
rect 488644 634946 488650 634948
rect 488717 634946 488783 634949
rect 488644 634944 488783 634946
rect 488644 634888 488722 634944
rect 488778 634888 488783 634944
rect 488644 634886 488783 634888
rect 488644 634884 488650 634886
rect 488717 634883 488783 634886
rect 506606 634884 506612 634948
rect 506676 634946 506682 634948
rect 506749 634946 506815 634949
rect 506676 634944 506815 634946
rect 506676 634888 506754 634944
rect 506810 634888 506815 634944
rect 506676 634886 506815 634888
rect 506676 634884 506682 634886
rect 506749 634883 506815 634886
rect 457805 634810 457871 634813
rect 457805 634808 460122 634810
rect 457805 634752 457810 634808
rect 457866 634752 460122 634808
rect 457805 634750 460122 634752
rect 457805 634747 457871 634750
rect 460062 634712 460122 634750
rect 321553 634538 321619 634541
rect 321553 634536 325036 634538
rect 321553 634480 321558 634536
rect 321614 634480 325036 634536
rect 321553 634478 325036 634480
rect 321553 634475 321619 634478
rect 59077 632906 59143 632909
rect 148593 632906 148659 632909
rect 238293 632906 238359 632909
rect 59077 632904 60076 632906
rect 59077 632848 59082 632904
rect 59138 632848 60076 632904
rect 59077 632846 60076 632848
rect 148593 632904 150052 632906
rect 148593 632848 148598 632904
rect 148654 632848 150052 632904
rect 148593 632846 150052 632848
rect 238293 632904 240032 632906
rect 238293 632848 238298 632904
rect 238354 632848 240032 632904
rect 238293 632846 240032 632848
rect 59077 632843 59143 632846
rect 148593 632843 148659 632846
rect 238293 632843 238359 632846
rect 212809 632498 212875 632501
rect 300945 632498 301011 632501
rect 210558 632496 212875 632498
rect 210558 632440 212814 632496
rect 212870 632440 212875 632496
rect 210558 632438 212875 632440
rect 123017 632226 123083 632229
rect 120796 632224 123083 632226
rect -960 632090 480 632180
rect 120796 632168 123022 632224
rect 123078 632168 123083 632224
rect 210558 632196 210618 632438
rect 212809 632435 212875 632438
rect 300718 632496 301011 632498
rect 300718 632440 300950 632496
rect 301006 632440 301011 632496
rect 300718 632438 301011 632440
rect 300718 632196 300778 632438
rect 300945 632435 301011 632438
rect 120796 632166 123083 632168
rect 123017 632163 123083 632166
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 509926 631954 509986 631992
rect 512177 631954 512243 631957
rect 509926 631952 512243 631954
rect 509926 631896 512182 631952
rect 512238 631896 512243 631952
rect 509926 631894 512243 631896
rect 512177 631891 512243 631894
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect 436185 630458 436251 630461
rect 433780 630456 436251 630458
rect 433780 630400 436190 630456
rect 436246 630400 436251 630456
rect 433780 630398 436251 630400
rect 436185 630395 436251 630398
rect 321553 629778 321619 629781
rect 321553 629776 325036 629778
rect 321553 629720 321558 629776
rect 321614 629720 325036 629776
rect 321553 629718 325036 629720
rect 321553 629715 321619 629718
rect 59261 629506 59327 629509
rect 147489 629506 147555 629509
rect 237373 629506 237439 629509
rect 59261 629504 60076 629506
rect 59261 629448 59266 629504
rect 59322 629448 60076 629504
rect 59261 629446 60076 629448
rect 147489 629504 150052 629506
rect 147489 629448 147494 629504
rect 147550 629448 150052 629504
rect 147489 629446 150052 629448
rect 237373 629504 240032 629506
rect 237373 629448 237378 629504
rect 237434 629448 240032 629504
rect 237373 629446 240032 629448
rect 59261 629443 59327 629446
rect 147489 629443 147555 629446
rect 237373 629443 237439 629446
rect 457713 629234 457779 629237
rect 457713 629232 460122 629234
rect 457713 629176 457718 629232
rect 457774 629176 460122 629232
rect 457713 629174 460122 629176
rect 457713 629171 457779 629174
rect 121729 628826 121795 628829
rect 120796 628824 121795 628826
rect 120796 628768 121734 628824
rect 121790 628768 121795 628824
rect 120796 628766 121795 628768
rect 121729 628763 121795 628766
rect 210742 628282 210802 628796
rect 212533 628282 212599 628285
rect 210742 628280 212599 628282
rect 210742 628224 212538 628280
rect 212594 628224 212599 628280
rect 210742 628222 212599 628224
rect 300718 628282 300778 628796
rect 460062 628592 460122 629174
rect 302233 628282 302299 628285
rect 300718 628280 302299 628282
rect 300718 628224 302238 628280
rect 302294 628224 302299 628280
rect 300718 628222 302299 628224
rect 212533 628219 212599 628222
rect 302233 628219 302299 628222
rect 57513 626786 57579 626789
rect 146293 626786 146359 626789
rect 237373 626786 237439 626789
rect 57513 626784 60076 626786
rect 57513 626728 57518 626784
rect 57574 626728 60076 626784
rect 57513 626726 60076 626728
rect 146293 626784 150052 626786
rect 146293 626728 146298 626784
rect 146354 626728 150052 626784
rect 146293 626726 150052 626728
rect 237373 626784 240032 626786
rect 237373 626728 237378 626784
rect 237434 626728 240032 626784
rect 237373 626726 240032 626728
rect 57513 626723 57579 626726
rect 146293 626723 146359 626726
rect 237373 626723 237439 626726
rect 512085 626514 512151 626517
rect 509926 626512 512151 626514
rect 509926 626456 512090 626512
rect 512146 626456 512151 626512
rect 509926 626454 512151 626456
rect 433333 626242 433399 626245
rect 433333 626240 433442 626242
rect 433333 626184 433338 626240
rect 433394 626184 433442 626240
rect 433333 626179 433442 626184
rect 123109 626106 123175 626109
rect 120796 626104 123175 626106
rect 120796 626048 123114 626104
rect 123170 626048 123175 626104
rect 120796 626046 123175 626048
rect 123109 626043 123175 626046
rect 210742 625698 210802 626076
rect 211245 625698 211311 625701
rect 210742 625696 211311 625698
rect 210742 625640 211250 625696
rect 211306 625640 211311 625696
rect 210742 625638 211311 625640
rect 300718 625698 300778 626076
rect 301037 625698 301103 625701
rect 300718 625696 301103 625698
rect 300718 625640 301042 625696
rect 301098 625640 301103 625696
rect 433382 625668 433442 626179
rect 509926 625872 509986 626454
rect 512085 626451 512151 626454
rect 300718 625638 301103 625640
rect 211245 625635 211311 625638
rect 301037 625635 301103 625638
rect 321553 625018 321619 625021
rect 321553 625016 325036 625018
rect 321553 624960 321558 625016
rect 321614 624960 325036 625016
rect 321553 624958 325036 624960
rect 321553 624955 321619 624958
rect 58893 623386 58959 623389
rect 146293 623386 146359 623389
rect 237373 623386 237439 623389
rect 58893 623384 60076 623386
rect 58893 623328 58898 623384
rect 58954 623328 60076 623384
rect 58893 623326 60076 623328
rect 146293 623384 150052 623386
rect 146293 623328 146298 623384
rect 146354 623328 150052 623384
rect 146293 623326 150052 623328
rect 237373 623384 240032 623386
rect 237373 623328 237378 623384
rect 237434 623328 240032 623384
rect 237373 623326 240032 623328
rect 58893 623323 58959 623326
rect 146293 623323 146359 623326
rect 237373 623323 237439 623326
rect 457621 623114 457687 623117
rect 457621 623112 460122 623114
rect 457621 623056 457626 623112
rect 457682 623056 460122 623112
rect 457621 623054 460122 623056
rect 457621 623051 457687 623054
rect 121637 622706 121703 622709
rect 120796 622704 121703 622706
rect 120796 622648 121642 622704
rect 121698 622648 121703 622704
rect 120796 622646 121703 622648
rect 121637 622643 121703 622646
rect 210742 622434 210802 622676
rect 212717 622434 212783 622437
rect 210742 622432 212783 622434
rect 210742 622376 212722 622432
rect 212778 622376 212783 622432
rect 210742 622374 212783 622376
rect 300718 622434 300778 622676
rect 460062 622472 460122 623054
rect 302325 622434 302391 622437
rect 300718 622432 302391 622434
rect 300718 622376 302330 622432
rect 302386 622376 302391 622432
rect 300718 622374 302391 622376
rect 212717 622371 212783 622374
rect 302325 622371 302391 622374
rect 436093 620938 436159 620941
rect 433780 620936 436159 620938
rect 433780 620880 436098 620936
rect 436154 620880 436159 620936
rect 433780 620878 436159 620880
rect 436093 620875 436159 620878
rect 59169 620666 59235 620669
rect 147397 620666 147463 620669
rect 237373 620666 237439 620669
rect 59169 620664 60076 620666
rect 59169 620608 59174 620664
rect 59230 620608 60076 620664
rect 59169 620606 60076 620608
rect 147397 620664 150052 620666
rect 147397 620608 147402 620664
rect 147458 620608 150052 620664
rect 147397 620606 150052 620608
rect 237373 620664 240032 620666
rect 237373 620608 237378 620664
rect 237434 620608 240032 620664
rect 237373 620606 240032 620608
rect 59169 620603 59235 620606
rect 147397 620603 147463 620606
rect 237373 620603 237439 620606
rect 321553 620258 321619 620261
rect 321553 620256 325036 620258
rect 321553 620200 321558 620256
rect 321614 620200 325036 620256
rect 321553 620198 325036 620200
rect 321553 620195 321619 620198
rect 123201 619986 123267 619989
rect 120796 619984 123267 619986
rect 120796 619928 123206 619984
rect 123262 619928 123267 619984
rect 120796 619926 123267 619928
rect 123201 619923 123267 619926
rect 210742 619714 210802 619956
rect 211429 619714 211495 619717
rect 210742 619712 211495 619714
rect 210742 619656 211434 619712
rect 211490 619656 211495 619712
rect 210742 619654 211495 619656
rect 300718 619714 300778 619956
rect 301129 619714 301195 619717
rect 300718 619712 301195 619714
rect 300718 619656 301134 619712
rect 301190 619656 301195 619712
rect 300718 619654 301195 619656
rect 211429 619651 211495 619654
rect 301129 619651 301195 619654
rect 511993 619578 512059 619581
rect 509926 619576 512059 619578
rect 509926 619520 511998 619576
rect 512054 619520 512059 619576
rect 509926 619518 512059 619520
rect -960 619020 480 619260
rect 509926 619072 509986 619518
rect 511993 619515 512059 619518
rect 583520 617388 584960 617628
rect 58985 617266 59051 617269
rect 148685 617266 148751 617269
rect 237373 617266 237439 617269
rect 58985 617264 60076 617266
rect 58985 617208 58990 617264
rect 59046 617208 60076 617264
rect 58985 617206 60076 617208
rect 148685 617264 150052 617266
rect 148685 617208 148690 617264
rect 148746 617208 150052 617264
rect 148685 617206 150052 617208
rect 237373 617264 240032 617266
rect 237373 617208 237378 617264
rect 237434 617208 240032 617264
rect 237373 617206 240032 617208
rect 58985 617203 59051 617206
rect 148685 617203 148751 617206
rect 237373 617203 237439 617206
rect 457529 616858 457595 616861
rect 457529 616856 460122 616858
rect 457529 616800 457534 616856
rect 457590 616800 460122 616856
rect 457529 616798 460122 616800
rect 457529 616795 457595 616798
rect 121821 616586 121887 616589
rect 120796 616584 121887 616586
rect 120796 616528 121826 616584
rect 121882 616528 121887 616584
rect 120796 616526 121887 616528
rect 121821 616523 121887 616526
rect 210742 616042 210802 616556
rect 211337 616042 211403 616045
rect 210742 616040 211403 616042
rect 210742 615984 211342 616040
rect 211398 615984 211403 616040
rect 210742 615982 211403 615984
rect 300718 616042 300778 616556
rect 460062 616352 460122 616798
rect 302417 616042 302483 616045
rect 300718 616040 302483 616042
rect 300718 615984 302422 616040
rect 302478 615984 302483 616040
rect 300718 615982 302483 615984
rect 211337 615979 211403 615982
rect 302417 615979 302483 615982
rect 433382 615909 433442 616148
rect 433333 615904 433442 615909
rect 433333 615848 433338 615904
rect 433394 615848 433442 615904
rect 433333 615846 433442 615848
rect 433333 615843 433399 615846
rect 321553 615498 321619 615501
rect 321553 615496 325036 615498
rect 321553 615440 321558 615496
rect 321614 615440 325036 615496
rect 321553 615438 325036 615440
rect 321553 615435 321619 615438
rect 57697 614546 57763 614549
rect 147213 614546 147279 614549
rect 238937 614546 239003 614549
rect 57697 614544 60076 614546
rect 57697 614488 57702 614544
rect 57758 614488 60076 614544
rect 57697 614486 60076 614488
rect 147213 614544 150052 614546
rect 147213 614488 147218 614544
rect 147274 614488 150052 614544
rect 147213 614486 150052 614488
rect 238937 614544 240032 614546
rect 238937 614488 238942 614544
rect 238998 614488 240032 614544
rect 238937 614486 240032 614488
rect 57697 614483 57763 614486
rect 147213 614483 147279 614486
rect 238937 614483 239003 614486
rect 120766 613325 120826 613836
rect 120766 613320 120875 613325
rect 120766 613264 120814 613320
rect 120870 613264 120875 613320
rect 120766 613262 120875 613264
rect 210742 613322 210802 613836
rect 213085 613322 213151 613325
rect 210742 613320 213151 613322
rect 210742 613264 213090 613320
rect 213146 613264 213151 613320
rect 210742 613262 213151 613264
rect 300718 613322 300778 613836
rect 302509 613322 302575 613325
rect 300718 613320 302575 613322
rect 300718 613264 302514 613320
rect 302570 613264 302575 613320
rect 300718 613262 302575 613264
rect 120809 613259 120875 613262
rect 213085 613259 213151 613262
rect 302509 613259 302575 613262
rect 509926 612778 509986 612952
rect 511993 612778 512059 612781
rect 509926 612776 512059 612778
rect 509926 612720 511998 612776
rect 512054 612720 512059 612776
rect 509926 612718 512059 612720
rect 511993 612715 512059 612718
rect 436134 611418 436140 611420
rect 433780 611358 436140 611418
rect 436134 611356 436140 611358
rect 436204 611356 436210 611420
rect 57881 611146 57947 611149
rect 146201 611146 146267 611149
rect 238017 611146 238083 611149
rect 57881 611144 60076 611146
rect 57881 611088 57886 611144
rect 57942 611088 60076 611144
rect 57881 611086 60076 611088
rect 146201 611144 150052 611146
rect 146201 611088 146206 611144
rect 146262 611088 150052 611144
rect 146201 611086 150052 611088
rect 238017 611144 240032 611146
rect 238017 611088 238022 611144
rect 238078 611088 240032 611144
rect 238017 611086 240032 611088
rect 57881 611083 57947 611086
rect 146201 611083 146267 611086
rect 238017 611083 238083 611086
rect 321553 610738 321619 610741
rect 321553 610736 325036 610738
rect 321553 610680 321558 610736
rect 321614 610680 325036 610736
rect 321553 610678 325036 610680
rect 321553 610675 321619 610678
rect 123385 610466 123451 610469
rect 120796 610464 123451 610466
rect 120796 610408 123390 610464
rect 123446 610408 123451 610464
rect 120796 610406 123451 610408
rect 123385 610403 123451 610406
rect 210742 610058 210802 610436
rect 212901 610058 212967 610061
rect 210742 610056 212967 610058
rect 210742 610000 212906 610056
rect 212962 610000 212967 610056
rect 210742 609998 212967 610000
rect 300718 610058 300778 610436
rect 301313 610058 301379 610061
rect 300718 610056 301379 610058
rect 300718 610000 301318 610056
rect 301374 610000 301379 610056
rect 300718 609998 301379 610000
rect 212901 609995 212967 609998
rect 301313 609995 301379 609998
rect 457621 608970 457687 608973
rect 460062 608970 460122 609552
rect 457621 608968 460122 608970
rect 457621 608912 457626 608968
rect 457682 608912 460122 608968
rect 457621 608910 460122 608912
rect 457621 608907 457687 608910
rect 58801 608426 58867 608429
rect 148409 608426 148475 608429
rect 237373 608426 237439 608429
rect 58801 608424 60076 608426
rect 58801 608368 58806 608424
rect 58862 608368 60076 608424
rect 58801 608366 60076 608368
rect 148409 608424 150052 608426
rect 148409 608368 148414 608424
rect 148470 608368 150052 608424
rect 148409 608366 150052 608368
rect 237373 608424 240032 608426
rect 237373 608368 237378 608424
rect 237434 608368 240032 608424
rect 237373 608366 240032 608368
rect 58801 608363 58867 608366
rect 148409 608363 148475 608366
rect 237373 608363 237439 608366
rect 123477 607746 123543 607749
rect 120796 607744 123543 607746
rect 120796 607688 123482 607744
rect 123538 607688 123543 607744
rect 120796 607686 123543 607688
rect 123477 607683 123543 607686
rect 210742 607338 210802 607716
rect 212993 607338 213059 607341
rect 210742 607336 213059 607338
rect 210742 607280 212998 607336
rect 213054 607280 213059 607336
rect 210742 607278 213059 607280
rect 300718 607338 300778 607716
rect 302693 607338 302759 607341
rect 300718 607336 302759 607338
rect 300718 607280 302698 607336
rect 302754 607280 302759 607336
rect 300718 607278 302759 607280
rect 212993 607275 213059 607278
rect 302693 607275 302759 607278
rect 436318 606658 436324 606660
rect 433780 606598 436324 606658
rect 436318 606596 436324 606598
rect 436388 606596 436394 606660
rect 509926 606386 509986 606832
rect 512177 606386 512243 606389
rect 509926 606384 512243 606386
rect 509926 606328 512182 606384
rect 512238 606328 512243 606384
rect 509926 606326 512243 606328
rect 512177 606323 512243 606326
rect -960 605964 480 606204
rect 321553 605978 321619 605981
rect 321553 605976 325036 605978
rect 321553 605920 321558 605976
rect 321614 605920 325036 605976
rect 321553 605918 325036 605920
rect 321553 605915 321619 605918
rect 57421 605026 57487 605029
rect 146293 605026 146359 605029
rect 237373 605026 237439 605029
rect 57421 605024 60076 605026
rect 57421 604968 57426 605024
rect 57482 604968 60076 605024
rect 57421 604966 60076 604968
rect 146293 605024 150052 605026
rect 146293 604968 146298 605024
rect 146354 604968 150052 605024
rect 146293 604966 150052 604968
rect 237373 605024 240032 605026
rect 237373 604968 237378 605024
rect 237434 604968 240032 605024
rect 237373 604966 240032 604968
rect 57421 604963 57487 604966
rect 146293 604963 146359 604966
rect 237373 604963 237439 604966
rect 124121 604346 124187 604349
rect 120796 604344 124187 604346
rect 120796 604288 124126 604344
rect 124182 604288 124187 604344
rect 120796 604286 124187 604288
rect 124121 604283 124187 604286
rect 210742 603802 210802 604316
rect 214005 603802 214071 603805
rect 210742 603800 214071 603802
rect 210742 603744 214010 603800
rect 214066 603744 214071 603800
rect 210742 603742 214071 603744
rect 300718 603802 300778 604316
rect 583520 604060 584960 604300
rect 302877 603802 302943 603805
rect 303153 603802 303219 603805
rect 300718 603800 303219 603802
rect 300718 603744 302882 603800
rect 302938 603744 303158 603800
rect 303214 603744 303219 603800
rect 300718 603742 303219 603744
rect 214005 603739 214071 603742
rect 302877 603739 302943 603742
rect 303153 603739 303219 603742
rect 457529 603122 457595 603125
rect 460062 603122 460122 603432
rect 457529 603120 460122 603122
rect 457529 603064 457534 603120
rect 457590 603064 460122 603120
rect 457529 603062 460122 603064
rect 457529 603059 457595 603062
rect 57697 602306 57763 602309
rect 147121 602306 147187 602309
rect 237373 602306 237439 602309
rect 57697 602304 60076 602306
rect 57697 602248 57702 602304
rect 57758 602248 60076 602304
rect 57697 602246 60076 602248
rect 147121 602304 150052 602306
rect 147121 602248 147126 602304
rect 147182 602248 150052 602304
rect 147121 602246 150052 602248
rect 237373 602304 240032 602306
rect 237373 602248 237378 602304
rect 237434 602248 240032 602304
rect 237373 602246 240032 602248
rect 57697 602243 57763 602246
rect 147121 602243 147187 602246
rect 237373 602243 237439 602246
rect 433382 601629 433442 601868
rect 122005 601626 122071 601629
rect 120796 601624 122071 601626
rect 120796 601568 122010 601624
rect 122066 601568 122071 601624
rect 433382 601624 433491 601629
rect 120796 601566 122071 601568
rect 122005 601563 122071 601566
rect 210742 601082 210802 601596
rect 211705 601082 211771 601085
rect 210742 601080 211771 601082
rect 210742 601024 211710 601080
rect 211766 601024 211771 601080
rect 210742 601022 211771 601024
rect 300718 601082 300778 601596
rect 433382 601568 433430 601624
rect 433486 601568 433491 601624
rect 433382 601566 433491 601568
rect 433425 601563 433491 601566
rect 324221 601218 324287 601221
rect 324221 601216 325036 601218
rect 324221 601160 324226 601216
rect 324282 601160 325036 601216
rect 324221 601158 325036 601160
rect 324221 601155 324287 601158
rect 301221 601082 301287 601085
rect 300718 601080 301287 601082
rect 300718 601024 301226 601080
rect 301282 601024 301287 601080
rect 300718 601022 301287 601024
rect 211705 601019 211771 601022
rect 301221 601019 301287 601022
rect 509926 600402 509986 600712
rect 512085 600402 512151 600405
rect 509926 600400 512151 600402
rect 509926 600344 512090 600400
rect 512146 600344 512151 600400
rect 509926 600342 512151 600344
rect 512085 600339 512151 600342
rect 57237 598906 57303 598909
rect 148501 598906 148567 598909
rect 237373 598906 237439 598909
rect 57237 598904 60076 598906
rect 57237 598848 57242 598904
rect 57298 598848 60076 598904
rect 57237 598846 60076 598848
rect 148501 598904 150052 598906
rect 148501 598848 148506 598904
rect 148562 598848 150052 598904
rect 148501 598846 150052 598848
rect 237373 598904 240032 598906
rect 237373 598848 237378 598904
rect 237434 598848 240032 598904
rect 237373 598846 240032 598848
rect 57237 598843 57303 598846
rect 148501 598843 148567 598846
rect 237373 598843 237439 598846
rect 121085 598226 121151 598229
rect 120796 598224 121151 598226
rect 120796 598168 121090 598224
rect 121146 598168 121151 598224
rect 120796 598166 121151 598168
rect 121085 598163 121151 598166
rect 210742 597682 210802 598196
rect 211613 597682 211679 597685
rect 210742 597680 211679 597682
rect 210742 597624 211618 597680
rect 211674 597624 211679 597680
rect 210742 597622 211679 597624
rect 300718 597682 300778 598196
rect 302601 597682 302667 597685
rect 300718 597680 302667 597682
rect 300718 597624 302606 597680
rect 302662 597624 302667 597680
rect 300718 597622 302667 597624
rect 211613 597619 211679 597622
rect 302601 597619 302667 597622
rect 457437 597546 457503 597549
rect 457437 597544 460122 597546
rect 457437 597488 457442 597544
rect 457498 597488 460122 597544
rect 457437 597486 460122 597488
rect 457437 597483 457503 597486
rect 460062 597312 460122 597486
rect 436093 597138 436159 597141
rect 433780 597136 436159 597138
rect 433780 597080 436098 597136
rect 436154 597080 436159 597136
rect 433780 597078 436159 597080
rect 436093 597075 436159 597078
rect 321553 596458 321619 596461
rect 321553 596456 325036 596458
rect 321553 596400 321558 596456
rect 321614 596400 325036 596456
rect 321553 596398 325036 596400
rect 321553 596395 321619 596398
rect 57145 596186 57211 596189
rect 147213 596186 147279 596189
rect 237373 596186 237439 596189
rect 57145 596184 60076 596186
rect 57145 596128 57150 596184
rect 57206 596128 60076 596184
rect 57145 596126 60076 596128
rect 147213 596184 150052 596186
rect 147213 596128 147218 596184
rect 147274 596128 150052 596184
rect 147213 596126 150052 596128
rect 237373 596184 240032 596186
rect 237373 596128 237378 596184
rect 237434 596128 240032 596184
rect 237373 596126 240032 596128
rect 57145 596123 57211 596126
rect 147213 596123 147279 596126
rect 237373 596123 237439 596126
rect 122097 595506 122163 595509
rect 120796 595504 122163 595506
rect 120796 595448 122102 595504
rect 122158 595448 122163 595504
rect 120796 595446 122163 595448
rect 122097 595443 122163 595446
rect 210742 594962 210802 595476
rect 211521 594962 211587 594965
rect 210742 594960 211587 594962
rect 210742 594904 211526 594960
rect 211582 594904 211587 594960
rect 210742 594902 211587 594904
rect 300718 594962 300778 595476
rect 302785 594962 302851 594965
rect 300718 594960 302851 594962
rect 300718 594904 302790 594960
rect 302846 594904 302851 594960
rect 300718 594902 302851 594904
rect 211521 594899 211587 594902
rect 302785 594899 302851 594902
rect 509926 594010 509986 594592
rect 512269 594010 512335 594013
rect 509926 594008 512335 594010
rect 509926 593952 512274 594008
rect 512330 593952 512335 594008
rect 509926 593950 512335 593952
rect 512269 593947 512335 593950
rect -960 592908 480 593148
rect 58709 592786 58775 592789
rect 146293 592786 146359 592789
rect 237373 592786 237439 592789
rect 58709 592784 60076 592786
rect 58709 592728 58714 592784
rect 58770 592728 60076 592784
rect 58709 592726 60076 592728
rect 146293 592784 150052 592786
rect 146293 592728 146298 592784
rect 146354 592728 150052 592784
rect 146293 592726 150052 592728
rect 237373 592784 240032 592786
rect 237373 592728 237378 592784
rect 237434 592728 240032 592784
rect 237373 592726 240032 592728
rect 58709 592723 58775 592726
rect 146293 592723 146359 592726
rect 237373 592723 237439 592726
rect 211797 592378 211863 592381
rect 301405 592378 301471 592381
rect 434805 592378 434871 592381
rect 210558 592376 211863 592378
rect 210558 592320 211802 592376
rect 211858 592320 211863 592376
rect 210558 592318 211863 592320
rect 122189 592106 122255 592109
rect 120796 592104 122255 592106
rect 120796 592048 122194 592104
rect 122250 592048 122255 592104
rect 210558 592076 210618 592318
rect 211797 592315 211863 592318
rect 300534 592376 301471 592378
rect 300534 592320 301410 592376
rect 301466 592320 301471 592376
rect 300534 592318 301471 592320
rect 433780 592376 434871 592378
rect 433780 592320 434810 592376
rect 434866 592320 434871 592376
rect 433780 592318 434871 592320
rect 300534 592076 300594 592318
rect 301405 592315 301471 592318
rect 434805 592315 434871 592318
rect 120796 592046 122255 592048
rect 122189 592043 122255 592046
rect 321553 591698 321619 591701
rect 321553 591696 325036 591698
rect 321553 591640 321558 591696
rect 321614 591640 325036 591696
rect 321553 591638 325036 591640
rect 321553 591635 321619 591638
rect 457437 590746 457503 590749
rect 460062 590746 460122 591192
rect 583520 590868 584960 591108
rect 457437 590744 460122 590746
rect 457437 590688 457442 590744
rect 457498 590688 460122 590744
rect 457437 590686 460122 590688
rect 457437 590683 457503 590686
rect 57053 590066 57119 590069
rect 146293 590066 146359 590069
rect 237373 590066 237439 590069
rect 57053 590064 60076 590066
rect 57053 590008 57058 590064
rect 57114 590008 60076 590064
rect 57053 590006 60076 590008
rect 146293 590064 150052 590066
rect 146293 590008 146298 590064
rect 146354 590008 150052 590064
rect 146293 590006 150052 590008
rect 237373 590064 240032 590066
rect 237373 590008 237378 590064
rect 237434 590008 240032 590064
rect 237373 590006 240032 590008
rect 57053 590003 57119 590006
rect 146293 590003 146359 590006
rect 237373 590003 237439 590006
rect 213177 589658 213243 589661
rect 301497 589658 301563 589661
rect 210558 589656 213243 589658
rect 210558 589600 213182 589656
rect 213238 589600 213243 589656
rect 210558 589598 213243 589600
rect 122281 589386 122347 589389
rect 120796 589384 122347 589386
rect 120796 589328 122286 589384
rect 122342 589328 122347 589384
rect 210558 589356 210618 589598
rect 213177 589595 213243 589598
rect 300534 589656 301563 589658
rect 300534 589600 301502 589656
rect 301558 589600 301563 589656
rect 300534 589598 301563 589600
rect 300534 589356 300594 589598
rect 301497 589595 301563 589598
rect 120796 589326 122347 589328
rect 122281 589323 122347 589326
rect 321553 586938 321619 586941
rect 433750 586938 433810 587588
rect 509926 587074 509986 587792
rect 509926 587014 512010 587074
rect 321553 586936 325036 586938
rect 321553 586880 321558 586936
rect 321614 586880 325036 586936
rect 321553 586878 325036 586880
rect 433750 586878 434730 586938
rect 321553 586875 321619 586878
rect 57329 586666 57395 586669
rect 146293 586666 146359 586669
rect 237373 586666 237439 586669
rect 57329 586664 60076 586666
rect 57329 586608 57334 586664
rect 57390 586608 60076 586664
rect 57329 586606 60076 586608
rect 146293 586664 150052 586666
rect 146293 586608 146298 586664
rect 146354 586608 150052 586664
rect 146293 586606 150052 586608
rect 237373 586664 240032 586666
rect 237373 586608 237378 586664
rect 237434 586608 240032 586664
rect 237373 586606 240032 586608
rect 57329 586603 57395 586606
rect 146293 586603 146359 586606
rect 237373 586603 237439 586606
rect 434670 586394 434730 586878
rect 436502 586468 436508 586532
rect 436572 586468 436578 586532
rect 436510 586394 436570 586468
rect 434670 586334 436570 586394
rect 511950 586394 512010 587014
rect 513281 586530 513347 586533
rect 513238 586528 513347 586530
rect 513238 586472 513286 586528
rect 513342 586472 513347 586528
rect 513238 586467 513347 586472
rect 513238 586394 513298 586467
rect 511950 586334 513298 586394
rect 123477 585986 123543 585989
rect 120796 585984 123543 585986
rect 120796 585928 123482 585984
rect 123538 585928 123543 585984
rect 120796 585926 123543 585928
rect 123477 585923 123543 585926
rect 210742 585445 210802 585956
rect 210742 585440 210851 585445
rect 210742 585384 210790 585440
rect 210846 585384 210851 585440
rect 210742 585382 210851 585384
rect 300718 585442 300778 585956
rect 302969 585442 303035 585445
rect 300718 585440 303035 585442
rect 300718 585384 302974 585440
rect 303030 585384 303035 585440
rect 300718 585382 303035 585384
rect 210785 585379 210851 585382
rect 302969 585379 303035 585382
rect 58525 583946 58591 583949
rect 147029 583946 147095 583949
rect 237373 583946 237439 583949
rect 58525 583944 60076 583946
rect 58525 583888 58530 583944
rect 58586 583888 60076 583944
rect 58525 583886 60076 583888
rect 147029 583944 150052 583946
rect 147029 583888 147034 583944
rect 147090 583888 150052 583944
rect 147029 583886 150052 583888
rect 237373 583944 240032 583946
rect 237373 583888 237378 583944
rect 237434 583888 240032 583944
rect 237373 583886 240032 583888
rect 58525 583883 58591 583886
rect 147029 583883 147095 583886
rect 237373 583883 237439 583886
rect 123569 583266 123635 583269
rect 120796 583264 123635 583266
rect 120796 583208 123574 583264
rect 123630 583208 123635 583264
rect 120796 583206 123635 583208
rect 123569 583203 123635 583206
rect 210742 582722 210802 583236
rect 213269 582722 213335 582725
rect 210742 582720 213335 582722
rect 210742 582664 213274 582720
rect 213330 582664 213335 582720
rect 210742 582662 213335 582664
rect 300718 582722 300778 583236
rect 301589 582722 301655 582725
rect 300718 582720 301655 582722
rect 300718 582664 301594 582720
rect 301650 582664 301655 582720
rect 300718 582662 301655 582664
rect 213269 582659 213335 582662
rect 301589 582659 301655 582662
rect 436185 582178 436251 582181
rect 433780 582176 436251 582178
rect 433780 582120 436190 582176
rect 436246 582120 436251 582176
rect 433780 582118 436251 582120
rect 436185 582115 436251 582118
rect 321553 581498 321619 581501
rect 321553 581496 325036 581498
rect 321553 581440 321558 581496
rect 321614 581440 325036 581496
rect 321553 581438 325036 581440
rect 321553 581435 321619 581438
rect 57697 580546 57763 580549
rect 237373 580546 237439 580549
rect 57697 580544 60076 580546
rect 57697 580488 57702 580544
rect 57758 580488 60076 580544
rect 237373 580544 240032 580546
rect 57697 580486 60076 580488
rect 149789 580510 149855 580513
rect 149789 580508 150052 580510
rect 57697 580483 57763 580486
rect 149789 580452 149794 580508
rect 149850 580452 150052 580508
rect 237373 580488 237378 580544
rect 237434 580488 240032 580544
rect 237373 580486 240032 580488
rect 237373 580483 237439 580486
rect 149789 580450 150052 580452
rect 149789 580447 149855 580450
rect 210877 580138 210943 580141
rect 303061 580138 303127 580141
rect 210742 580136 210943 580138
rect -960 580002 480 580092
rect 210742 580080 210882 580136
rect 210938 580080 210943 580136
rect 210742 580078 210943 580080
rect 3785 580002 3851 580005
rect -960 580000 3851 580002
rect -960 579944 3790 580000
rect 3846 579944 3851 580000
rect -960 579942 3851 579944
rect -960 579852 480 579942
rect 3785 579939 3851 579942
rect 121913 579866 121979 579869
rect 120796 579864 121979 579866
rect 120796 579808 121918 579864
rect 121974 579808 121979 579864
rect 210742 579836 210802 580078
rect 210877 580075 210943 580078
rect 300534 580136 303127 580138
rect 300534 580080 303066 580136
rect 303122 580080 303127 580136
rect 300534 580078 303127 580080
rect 300534 579836 300594 580078
rect 303061 580075 303127 580078
rect 120796 579806 121979 579808
rect 121913 579803 121979 579806
rect 237373 577826 237439 577829
rect 237373 577824 240032 577826
rect 59537 577790 59603 577793
rect 149605 577790 149671 577793
rect 59537 577788 60076 577790
rect 59537 577732 59542 577788
rect 59598 577732 60076 577788
rect 59537 577730 60076 577732
rect 149605 577788 150052 577790
rect 149605 577732 149610 577788
rect 149666 577732 150052 577788
rect 237373 577768 237378 577824
rect 237434 577768 240032 577824
rect 237373 577766 240032 577768
rect 237373 577763 237439 577766
rect 149605 577730 150052 577732
rect 59537 577727 59603 577730
rect 149605 577727 149671 577730
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect 436277 577418 436343 577421
rect 433780 577416 436343 577418
rect 433780 577360 436282 577416
rect 436338 577360 436343 577416
rect 433780 577358 436343 577360
rect 436277 577355 436343 577358
rect 120766 576877 120826 577116
rect 120717 576872 120826 576877
rect 120717 576816 120722 576872
rect 120778 576816 120826 576872
rect 120717 576814 120826 576816
rect 210742 576874 210802 577116
rect 300718 576877 300778 577116
rect 210969 576874 211035 576877
rect 210742 576872 211035 576874
rect 210742 576816 210974 576872
rect 211030 576816 211035 576872
rect 210742 576814 211035 576816
rect 120717 576811 120783 576814
rect 210969 576811 211035 576814
rect 300669 576872 300778 576877
rect 300669 576816 300674 576872
rect 300730 576816 300778 576872
rect 300669 576814 300778 576816
rect 300669 576811 300735 576814
rect 321001 576738 321067 576741
rect 321001 576736 325036 576738
rect 321001 576680 321006 576736
rect 321062 576680 325036 576736
rect 321001 576678 325036 576680
rect 321001 576675 321067 576678
rect 436369 572658 436435 572661
rect 433780 572656 436435 572658
rect 433780 572600 436374 572656
rect 436430 572600 436435 572656
rect 433780 572598 436435 572600
rect 436369 572595 436435 572598
rect 321553 571978 321619 571981
rect 321553 571976 325036 571978
rect 321553 571920 321558 571976
rect 321614 571920 325036 571976
rect 321553 571918 325036 571920
rect 321553 571915 321619 571918
rect 433566 567493 433626 567868
rect 433517 567488 433626 567493
rect 433517 567432 433522 567488
rect 433578 567432 433626 567488
rect 433517 567430 433626 567432
rect 433517 567427 433583 567430
rect 321553 567218 321619 567221
rect 321553 567216 325036 567218
rect 321553 567160 321558 567216
rect 321614 567160 325036 567216
rect 321553 567158 325036 567160
rect 321553 567155 321619 567158
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect 436461 563138 436527 563141
rect 433780 563136 436527 563138
rect 433780 563080 436466 563136
rect 436522 563080 436527 563136
rect 433780 563078 436527 563080
rect 436461 563075 436527 563078
rect 321553 562458 321619 562461
rect 321553 562456 325036 562458
rect 321553 562400 321558 562456
rect 321614 562400 325036 562456
rect 321553 562398 325036 562400
rect 321553 562395 321619 562398
rect 436553 558378 436619 558381
rect 433780 558376 436619 558378
rect 433780 558320 436558 558376
rect 436614 558320 436619 558376
rect 433780 558318 436619 558320
rect 436553 558315 436619 558318
rect 321553 557698 321619 557701
rect 321553 557696 325036 557698
rect 321553 557640 321558 557696
rect 321614 557640 325036 557696
rect 321553 557638 325036 557640
rect 321553 557635 321619 557638
rect -960 553740 480 553980
rect 436645 553618 436711 553621
rect 433780 553616 436711 553618
rect 433780 553560 436650 553616
rect 436706 553560 436711 553616
rect 433780 553558 436711 553560
rect 436645 553555 436711 553558
rect 321553 552938 321619 552941
rect 321553 552936 325036 552938
rect 321553 552880 321558 552936
rect 321614 552880 325036 552936
rect 321553 552878 325036 552880
rect 321553 552875 321619 552878
rect 583520 551020 584960 551260
rect 238661 550082 238727 550085
rect 301681 550082 301747 550085
rect 238661 550080 301747 550082
rect 238661 550024 238666 550080
rect 238722 550024 301686 550080
rect 301742 550024 301747 550080
rect 238661 550022 301747 550024
rect 238661 550019 238727 550022
rect 301681 550019 301747 550022
rect 298093 549946 298159 549949
rect 322197 549946 322263 549949
rect 298093 549944 322263 549946
rect 298093 549888 298098 549944
rect 298154 549888 322202 549944
rect 322258 549888 322263 549944
rect 298093 549886 322263 549888
rect 298093 549883 298159 549886
rect 322197 549883 322263 549886
rect 255129 549810 255195 549813
rect 323945 549810 324011 549813
rect 255129 549808 324011 549810
rect 255129 549752 255134 549808
rect 255190 549752 323950 549808
rect 324006 549752 324011 549808
rect 255129 549750 324011 549752
rect 255129 549747 255195 549750
rect 323945 549747 324011 549750
rect 248689 549674 248755 549677
rect 300393 549674 300459 549677
rect 248689 549672 300459 549674
rect 248689 549616 248694 549672
rect 248750 549616 300398 549672
rect 300454 549616 300459 549672
rect 248689 549614 300459 549616
rect 248689 549611 248755 549614
rect 300393 549611 300459 549614
rect 294505 549538 294571 549541
rect 324814 549538 324820 549540
rect 294505 549536 324820 549538
rect 294505 549480 294510 549536
rect 294566 549480 324820 549536
rect 294505 549478 324820 549480
rect 294505 549475 294571 549478
rect 324814 549476 324820 549478
rect 324884 549476 324890 549540
rect 293125 549402 293191 549405
rect 301497 549402 301563 549405
rect 293125 549400 301563 549402
rect 293125 549344 293130 549400
rect 293186 549344 301502 549400
rect 301558 549344 301563 549400
rect 293125 549342 301563 549344
rect 293125 549339 293191 549342
rect 301497 549339 301563 549342
rect 436737 548858 436803 548861
rect 433780 548856 436803 548858
rect 433780 548800 436742 548856
rect 436798 548800 436803 548856
rect 433780 548798 436803 548800
rect 436737 548795 436803 548798
rect 321553 548178 321619 548181
rect 321553 548176 325036 548178
rect 321553 548120 321558 548176
rect 321614 548120 325036 548176
rect 321553 548118 325036 548120
rect 321553 548115 321619 548118
rect 3509 548042 3575 548045
rect 322197 548042 322263 548045
rect 3509 548040 322263 548042
rect 3509 547984 3514 548040
rect 3570 547984 322202 548040
rect 322258 547984 322263 548040
rect 3509 547982 322263 547984
rect 3509 547979 3575 547982
rect 322197 547979 322263 547982
rect 436829 544098 436895 544101
rect 433780 544096 436895 544098
rect 433780 544040 436834 544096
rect 436890 544040 436895 544096
rect 433780 544038 436895 544040
rect 436829 544035 436895 544038
rect 321553 543418 321619 543421
rect 321553 543416 325036 543418
rect 321553 543360 321558 543416
rect 321614 543360 325036 543416
rect 321553 543358 325036 543360
rect 321553 543355 321619 543358
rect -960 540684 480 540924
rect 302785 540426 302851 540429
rect 299828 540424 302851 540426
rect 299828 540368 302790 540424
rect 302846 540368 302851 540424
rect 299828 540366 302851 540368
rect 302785 540363 302851 540366
rect 434897 539338 434963 539341
rect 433780 539336 434963 539338
rect 433780 539280 434902 539336
rect 434958 539280 434963 539336
rect 433780 539278 434963 539280
rect 434897 539275 434963 539278
rect 321553 538658 321619 538661
rect 321553 538656 325036 538658
rect 321553 538600 321558 538656
rect 321614 538600 325036 538656
rect 321553 538598 325036 538600
rect 321553 538595 321619 538598
rect 583520 537692 584960 537932
rect 436921 534578 436987 534581
rect 433780 534576 436987 534578
rect 433780 534520 436926 534576
rect 436982 534520 436987 534576
rect 433780 534518 436987 534520
rect 436921 534515 436987 534518
rect 322105 533898 322171 533901
rect 322105 533896 325036 533898
rect 322105 533840 322110 533896
rect 322166 533840 325036 533896
rect 322105 533838 325036 533840
rect 322105 533835 322171 533838
rect 434621 529818 434687 529821
rect 433780 529816 434687 529818
rect 433780 529760 434626 529816
rect 434682 529760 434687 529816
rect 433780 529758 434687 529760
rect 434621 529755 434687 529758
rect 324814 529484 324820 529548
rect 324884 529546 324890 529548
rect 500953 529546 501019 529549
rect 324884 529544 501019 529546
rect 324884 529488 500958 529544
rect 501014 529488 501019 529544
rect 324884 529486 501019 529488
rect 324884 529484 324890 529486
rect 500953 529483 501019 529486
rect 300393 528458 300459 528461
rect 436318 528458 436324 528460
rect 300393 528456 436324 528458
rect 300393 528400 300398 528456
rect 300454 528400 436324 528456
rect 300393 528398 436324 528400
rect 300393 528395 300459 528398
rect 436318 528396 436324 528398
rect 436388 528396 436394 528460
rect 301681 528322 301747 528325
rect 436502 528322 436508 528324
rect 301681 528320 436508 528322
rect 301681 528264 301686 528320
rect 301742 528264 436508 528320
rect 301681 528262 436508 528264
rect 301681 528259 301747 528262
rect 436502 528260 436508 528262
rect 436572 528260 436578 528324
rect 323945 528186 324011 528189
rect 436134 528186 436140 528188
rect 323945 528184 436140 528186
rect 323945 528128 323950 528184
rect 324006 528128 436140 528184
rect 323945 528126 436140 528128
rect 323945 528123 324011 528126
rect 436134 528124 436140 528126
rect 436204 528124 436210 528188
rect -960 527764 480 528004
rect 304257 527098 304323 527101
rect 424501 527098 424567 527101
rect 304257 527096 424567 527098
rect 304257 527040 304262 527096
rect 304318 527040 424506 527096
rect 424562 527040 424567 527096
rect 304257 527038 424567 527040
rect 304257 527035 304323 527038
rect 424501 527035 424567 527038
rect 321185 526962 321251 526965
rect 429193 526962 429259 526965
rect 321185 526960 429259 526962
rect 321185 526904 321190 526960
rect 321246 526904 429198 526960
rect 429254 526904 429259 526960
rect 321185 526902 429259 526904
rect 321185 526899 321251 526902
rect 429193 526899 429259 526902
rect 322197 526826 322263 526829
rect 360745 526826 360811 526829
rect 322197 526824 360811 526826
rect 322197 526768 322202 526824
rect 322258 526768 360750 526824
rect 360806 526768 360811 526824
rect 322197 526766 360811 526768
rect 322197 526763 322263 526766
rect 360745 526763 360811 526766
rect 324037 526690 324103 526693
rect 342713 526690 342779 526693
rect 324037 526688 342779 526690
rect 324037 526632 324042 526688
rect 324098 526632 342718 526688
rect 342774 526632 342779 526688
rect 324037 526630 342779 526632
rect 324037 526627 324103 526630
rect 342713 526627 342779 526630
rect 302877 525466 302943 525469
rect 299828 525464 302943 525466
rect 299828 525408 302882 525464
rect 302938 525408 302943 525464
rect 299828 525406 302943 525408
rect 302877 525403 302943 525406
rect 583520 524364 584960 524604
rect 363454 523636 363460 523700
rect 363524 523698 363530 523700
rect 397453 523698 397519 523701
rect 363524 523696 397519 523698
rect 363524 523640 397458 523696
rect 397514 523640 397519 523696
rect 363524 523638 397519 523640
rect 363524 523636 363530 523638
rect 397453 523635 397519 523638
rect 360694 518060 360700 518124
rect 360764 518122 360770 518124
rect 506473 518122 506539 518125
rect 360764 518120 506539 518122
rect 360764 518064 506478 518120
rect 506534 518064 506539 518120
rect 360764 518062 506539 518064
rect 360764 518060 360770 518062
rect 506473 518059 506539 518062
rect 57881 517986 57947 517989
rect 57881 517984 60076 517986
rect 57881 517928 57886 517984
rect 57942 517928 60076 517984
rect 57881 517926 60076 517928
rect 57881 517923 57947 517926
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 303337 510506 303403 510509
rect 299828 510504 303403 510506
rect 299828 510448 303342 510504
rect 303398 510448 303403 510504
rect 299828 510446 303403 510448
rect 303337 510443 303403 510446
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 302233 495546 302299 495549
rect 299828 495544 302299 495546
rect 299828 495488 302238 495544
rect 302294 495488 302299 495544
rect 299828 495486 302299 495488
rect 302233 495483 302299 495486
rect 367686 489092 367692 489156
rect 367756 489154 367762 489156
rect 476062 489154 476068 489156
rect 367756 489094 476068 489154
rect 367756 489092 367762 489094
rect 476062 489092 476068 489094
rect 476132 489092 476138 489156
rect -960 488596 480 488836
rect 364926 487732 364932 487796
rect 364996 487794 365002 487796
rect 511993 487794 512059 487797
rect 364996 487792 512059 487794
rect 364996 487736 511998 487792
rect 512054 487736 512059 487792
rect 364996 487734 512059 487736
rect 364996 487732 365002 487734
rect 511993 487731 512059 487734
rect 365110 486508 365116 486572
rect 365180 486570 365186 486572
rect 457529 486570 457595 486573
rect 365180 486568 457595 486570
rect 365180 486512 457534 486568
rect 457590 486512 457595 486568
rect 365180 486510 457595 486512
rect 365180 486508 365186 486510
rect 457529 486507 457595 486510
rect 206134 486372 206140 486436
rect 206204 486434 206210 486436
rect 488574 486434 488580 486436
rect 206204 486374 488580 486434
rect 206204 486372 206210 486374
rect 488574 486372 488580 486374
rect 488644 486372 488650 486436
rect 59302 485692 59308 485756
rect 59372 485754 59378 485756
rect 76005 485754 76071 485757
rect 59372 485694 70410 485754
rect 59372 485692 59378 485694
rect 55070 485556 55076 485620
rect 55140 485618 55146 485620
rect 65425 485618 65491 485621
rect 55140 485616 65491 485618
rect 55140 485560 65430 485616
rect 65486 485560 65491 485616
rect 55140 485558 65491 485560
rect 70350 485618 70410 485694
rect 72742 485752 76071 485754
rect 72742 485696 76010 485752
rect 76066 485696 76071 485752
rect 72742 485694 76071 485696
rect 72509 485618 72575 485621
rect 70350 485616 72575 485618
rect 70350 485560 72514 485616
rect 72570 485560 72575 485616
rect 70350 485558 72575 485560
rect 55140 485556 55146 485558
rect 65425 485555 65491 485558
rect 72509 485555 72575 485558
rect 55622 485420 55628 485484
rect 55692 485482 55698 485484
rect 72742 485482 72802 485694
rect 76005 485691 76071 485694
rect 187049 485754 187115 485757
rect 199326 485754 199332 485756
rect 187049 485752 199332 485754
rect 187049 485696 187054 485752
rect 187110 485696 199332 485752
rect 187049 485694 199332 485696
rect 187049 485691 187115 485694
rect 199326 485692 199332 485694
rect 199396 485692 199402 485756
rect 73337 485618 73403 485621
rect 78673 485618 78739 485621
rect 73337 485616 78739 485618
rect 73337 485560 73342 485616
rect 73398 485560 78678 485616
rect 78734 485560 78739 485616
rect 73337 485558 78739 485560
rect 73337 485555 73403 485558
rect 78673 485555 78739 485558
rect 171133 485618 171199 485621
rect 198038 485618 198044 485620
rect 171133 485616 198044 485618
rect 171133 485560 171138 485616
rect 171194 485560 198044 485616
rect 171133 485558 198044 485560
rect 171133 485555 171199 485558
rect 198038 485556 198044 485558
rect 198108 485556 198114 485620
rect 235809 485618 235875 485621
rect 357934 485618 357940 485620
rect 235809 485616 357940 485618
rect 235809 485560 235814 485616
rect 235870 485560 357940 485616
rect 235809 485558 357940 485560
rect 235809 485555 235875 485558
rect 357934 485556 357940 485558
rect 358004 485556 358010 485620
rect 55692 485422 72802 485482
rect 73245 485482 73311 485485
rect 77753 485482 77819 485485
rect 73245 485480 77819 485482
rect 73245 485424 73250 485480
rect 73306 485424 77758 485480
rect 77814 485424 77819 485480
rect 73245 485422 77819 485424
rect 55692 485420 55698 485422
rect 73245 485419 73311 485422
rect 77753 485419 77819 485422
rect 163681 485482 163747 485485
rect 196566 485482 196572 485484
rect 163681 485480 196572 485482
rect 163681 485424 163686 485480
rect 163742 485424 196572 485480
rect 163681 485422 196572 485424
rect 163681 485419 163747 485422
rect 196566 485420 196572 485422
rect 196636 485420 196642 485484
rect 212533 485482 212599 485485
rect 213678 485482 213684 485484
rect 212533 485480 213684 485482
rect 212533 485424 212538 485480
rect 212594 485424 213684 485480
rect 212533 485422 213684 485424
rect 212533 485419 212599 485422
rect 213678 485420 213684 485422
rect 213748 485420 213754 485484
rect 233233 485482 233299 485485
rect 367870 485482 367876 485484
rect 233233 485480 367876 485482
rect 233233 485424 233238 485480
rect 233294 485424 367876 485480
rect 233233 485422 367876 485424
rect 233233 485419 233299 485422
rect 367870 485420 367876 485422
rect 367940 485420 367946 485484
rect 51942 485284 51948 485348
rect 52012 485346 52018 485348
rect 63217 485346 63283 485349
rect 52012 485344 63283 485346
rect 52012 485288 63222 485344
rect 63278 485288 63283 485344
rect 52012 485286 63283 485288
rect 52012 485284 52018 485286
rect 63217 485283 63283 485286
rect 65425 485346 65491 485349
rect 73797 485346 73863 485349
rect 65425 485344 73863 485346
rect 65425 485288 65430 485344
rect 65486 485288 73802 485344
rect 73858 485288 73863 485344
rect 65425 485286 73863 485288
rect 65425 485283 65491 485286
rect 73797 485283 73863 485286
rect 145649 485346 145715 485349
rect 197854 485346 197860 485348
rect 145649 485344 197860 485346
rect 145649 485288 145654 485344
rect 145710 485288 197860 485344
rect 145649 485286 197860 485288
rect 145649 485283 145715 485286
rect 197854 485284 197860 485286
rect 197924 485284 197930 485348
rect 200481 485346 200547 485349
rect 201350 485346 201356 485348
rect 200481 485344 201356 485346
rect 200481 485288 200486 485344
rect 200542 485288 201356 485344
rect 200481 485286 201356 485288
rect 200481 485283 200547 485286
rect 201350 485284 201356 485286
rect 201420 485284 201426 485348
rect 208485 485346 208551 485349
rect 209630 485346 209636 485348
rect 208485 485344 209636 485346
rect 208485 485288 208490 485344
rect 208546 485288 209636 485344
rect 208485 485286 209636 485288
rect 208485 485283 208551 485286
rect 209630 485284 209636 485286
rect 209700 485284 209706 485348
rect 211153 485346 211219 485349
rect 211654 485346 211660 485348
rect 211153 485344 211660 485346
rect 211153 485288 211158 485344
rect 211214 485288 211660 485344
rect 211153 485286 211660 485288
rect 211153 485283 211219 485286
rect 211654 485284 211660 485286
rect 211724 485284 211730 485348
rect 235901 485346 235967 485349
rect 371734 485346 371740 485348
rect 235901 485344 371740 485346
rect 235901 485288 235906 485344
rect 235962 485288 371740 485344
rect 235901 485286 371740 485288
rect 235901 485283 235967 485286
rect 371734 485284 371740 485286
rect 371804 485284 371810 485348
rect 53230 485148 53236 485212
rect 53300 485210 53306 485212
rect 77293 485210 77359 485213
rect 53300 485208 77359 485210
rect 53300 485152 77298 485208
rect 77354 485152 77359 485208
rect 53300 485150 77359 485152
rect 53300 485148 53306 485150
rect 77293 485147 77359 485150
rect 147581 485210 147647 485213
rect 200798 485210 200804 485212
rect 147581 485208 200804 485210
rect 147581 485152 147586 485208
rect 147642 485152 200804 485208
rect 147581 485150 200804 485152
rect 147581 485147 147647 485150
rect 200798 485148 200804 485150
rect 200868 485148 200874 485212
rect 201493 485210 201559 485213
rect 202638 485210 202644 485212
rect 201493 485208 202644 485210
rect 201493 485152 201498 485208
rect 201554 485152 202644 485208
rect 201493 485150 202644 485152
rect 201493 485147 201559 485150
rect 202638 485148 202644 485150
rect 202708 485148 202714 485212
rect 204253 485210 204319 485213
rect 205214 485210 205220 485212
rect 204253 485208 205220 485210
rect 204253 485152 204258 485208
rect 204314 485152 205220 485208
rect 204253 485150 205220 485152
rect 204253 485147 204319 485150
rect 205214 485148 205220 485150
rect 205284 485148 205290 485212
rect 234337 485210 234403 485213
rect 375966 485210 375972 485212
rect 234337 485208 375972 485210
rect 234337 485152 234342 485208
rect 234398 485152 375972 485208
rect 234337 485150 375972 485152
rect 234337 485147 234403 485150
rect 375966 485148 375972 485150
rect 376036 485148 376042 485212
rect 57830 485012 57836 485076
rect 57900 485074 57906 485076
rect 91369 485074 91435 485077
rect 57900 485072 91435 485074
rect 57900 485016 91374 485072
rect 91430 485016 91435 485072
rect 57900 485014 91435 485016
rect 57900 485012 57906 485014
rect 91369 485011 91435 485014
rect 145465 485074 145531 485077
rect 200614 485074 200620 485076
rect 145465 485072 200620 485074
rect 145465 485016 145470 485072
rect 145526 485016 200620 485072
rect 145465 485014 200620 485016
rect 145465 485011 145531 485014
rect 200614 485012 200620 485014
rect 200684 485012 200690 485076
rect 202873 485074 202939 485077
rect 216990 485074 216996 485076
rect 202873 485072 216996 485074
rect 202873 485016 202878 485072
rect 202934 485016 216996 485072
rect 202873 485014 216996 485016
rect 202873 485011 202939 485014
rect 216990 485012 216996 485014
rect 217060 485012 217066 485076
rect 219198 485012 219204 485076
rect 219268 485074 219274 485076
rect 226149 485074 226215 485077
rect 219268 485072 226215 485074
rect 219268 485016 226154 485072
rect 226210 485016 226215 485072
rect 219268 485014 226215 485016
rect 219268 485012 219274 485014
rect 226149 485011 226215 485014
rect 232313 485074 232379 485077
rect 374678 485074 374684 485076
rect 232313 485072 374684 485074
rect 232313 485016 232318 485072
rect 232374 485016 374684 485072
rect 232313 485014 374684 485016
rect 232313 485011 232379 485014
rect 374678 485012 374684 485014
rect 374748 485012 374754 485076
rect 59118 484876 59124 484940
rect 59188 484938 59194 484940
rect 68921 484938 68987 484941
rect 59188 484936 68987 484938
rect 59188 484880 68926 484936
rect 68982 484880 68987 484936
rect 59188 484878 68987 484880
rect 59188 484876 59194 484878
rect 68921 484875 68987 484878
rect 185669 484938 185735 484941
rect 196750 484938 196756 484940
rect 185669 484936 196756 484938
rect 185669 484880 185674 484936
rect 185730 484880 196756 484936
rect 185669 484878 196756 484880
rect 185669 484875 185735 484878
rect 196750 484876 196756 484878
rect 196820 484876 196826 484940
rect 197353 484938 197419 484941
rect 198406 484938 198412 484940
rect 197353 484936 198412 484938
rect 197353 484880 197358 484936
rect 197414 484880 198412 484936
rect 197353 484878 198412 484880
rect 197353 484875 197419 484878
rect 198406 484876 198412 484878
rect 198476 484876 198482 484940
rect 204253 484938 204319 484941
rect 205398 484938 205404 484940
rect 204253 484936 205404 484938
rect 204253 484880 204258 484936
rect 204314 484880 205404 484936
rect 204253 484878 205404 484880
rect 204253 484875 204319 484878
rect 205398 484876 205404 484878
rect 205468 484876 205474 484940
rect 63217 484802 63283 484805
rect 74257 484802 74323 484805
rect 63217 484800 74323 484802
rect 63217 484744 63222 484800
rect 63278 484744 74262 484800
rect 74318 484744 74323 484800
rect 63217 484742 74323 484744
rect 63217 484739 63283 484742
rect 74257 484739 74323 484742
rect 197445 484802 197511 484805
rect 198590 484802 198596 484804
rect 197445 484800 198596 484802
rect 197445 484744 197450 484800
rect 197506 484744 198596 484800
rect 197445 484742 198596 484744
rect 197445 484739 197511 484742
rect 198590 484740 198596 484742
rect 198660 484740 198666 484804
rect 205633 484802 205699 484805
rect 206686 484802 206692 484804
rect 205633 484800 206692 484802
rect 205633 484744 205638 484800
rect 205694 484744 206692 484800
rect 205633 484742 206692 484744
rect 205633 484739 205699 484742
rect 206686 484740 206692 484742
rect 206756 484740 206762 484804
rect 211153 484802 211219 484805
rect 212390 484802 212396 484804
rect 211153 484800 212396 484802
rect 211153 484744 211158 484800
rect 211214 484744 212396 484800
rect 211153 484742 212396 484744
rect 211153 484739 211219 484742
rect 212390 484740 212396 484742
rect 212460 484740 212466 484804
rect 50286 484468 50292 484532
rect 50356 484530 50362 484532
rect 50613 484530 50679 484533
rect 50889 484532 50955 484533
rect 50838 484530 50844 484532
rect 50356 484528 50679 484530
rect 50356 484472 50618 484528
rect 50674 484472 50679 484528
rect 50356 484470 50679 484472
rect 50798 484470 50844 484530
rect 50908 484528 50955 484532
rect 50950 484472 50955 484528
rect 50356 484468 50362 484470
rect 50613 484467 50679 484470
rect 50838 484468 50844 484470
rect 50908 484468 50955 484472
rect 50889 484467 50955 484468
rect 214833 484530 214899 484533
rect 217542 484530 217548 484532
rect 214833 484528 217548 484530
rect 214833 484472 214838 484528
rect 214894 484472 217548 484528
rect 214833 484470 217548 484472
rect 214833 484467 214899 484470
rect 217542 484468 217548 484470
rect 217612 484468 217618 484532
rect 219934 484468 219940 484532
rect 220004 484530 220010 484532
rect 224861 484530 224927 484533
rect 220004 484528 224927 484530
rect 220004 484472 224866 484528
rect 224922 484472 224927 484528
rect 583520 484516 584960 484756
rect 220004 484470 224927 484472
rect 220004 484468 220010 484470
rect 224861 484467 224927 484470
rect 155861 483850 155927 483853
rect 213862 483850 213868 483852
rect 155861 483848 213868 483850
rect 155861 483792 155866 483848
rect 155922 483792 213868 483848
rect 155861 483790 213868 483792
rect 155861 483787 155927 483790
rect 213862 483788 213868 483790
rect 213932 483788 213938 483852
rect 228449 483850 228515 483853
rect 370446 483850 370452 483852
rect 228449 483848 370452 483850
rect 228449 483792 228454 483848
rect 228510 483792 370452 483848
rect 228449 483790 370452 483792
rect 228449 483787 228515 483790
rect 370446 483788 370452 483790
rect 370516 483788 370522 483852
rect 144361 483714 144427 483717
rect 214598 483714 214604 483716
rect 144361 483712 214604 483714
rect 144361 483656 144366 483712
rect 144422 483656 214604 483712
rect 144361 483654 214604 483656
rect 144361 483651 144427 483654
rect 214598 483652 214604 483654
rect 214668 483652 214674 483716
rect 231393 483714 231459 483717
rect 374494 483714 374500 483716
rect 231393 483712 374500 483714
rect 231393 483656 231398 483712
rect 231454 483656 374500 483712
rect 231393 483654 374500 483656
rect 231393 483651 231459 483654
rect 374494 483652 374500 483654
rect 374564 483652 374570 483716
rect 46790 482700 46796 482764
rect 46860 482762 46866 482764
rect 66345 482762 66411 482765
rect 46860 482760 66411 482762
rect 46860 482704 66350 482760
rect 66406 482704 66411 482760
rect 46860 482702 66411 482704
rect 46860 482700 46866 482702
rect 66345 482699 66411 482702
rect 57094 482564 57100 482628
rect 57164 482626 57170 482628
rect 121361 482626 121427 482629
rect 57164 482624 121427 482626
rect 57164 482568 121366 482624
rect 121422 482568 121427 482624
rect 57164 482566 121427 482568
rect 57164 482564 57170 482566
rect 121361 482563 121427 482566
rect 47945 482490 48011 482493
rect 120441 482490 120507 482493
rect 47945 482488 120507 482490
rect 47945 482432 47950 482488
rect 48006 482432 120446 482488
rect 120502 482432 120507 482488
rect 47945 482430 120507 482432
rect 47945 482427 48011 482430
rect 120441 482427 120507 482430
rect 256233 482490 256299 482493
rect 359406 482490 359412 482492
rect 256233 482488 359412 482490
rect 256233 482432 256238 482488
rect 256294 482432 359412 482488
rect 256233 482430 359412 482432
rect 256233 482427 256299 482430
rect 359406 482428 359412 482430
rect 359476 482428 359482 482492
rect 46841 482354 46907 482357
rect 127065 482354 127131 482357
rect 46841 482352 127131 482354
rect 46841 482296 46846 482352
rect 46902 482296 127070 482352
rect 127126 482296 127131 482352
rect 46841 482294 127131 482296
rect 46841 482291 46907 482294
rect 127065 482291 127131 482294
rect 155217 482354 155283 482357
rect 215334 482354 215340 482356
rect 155217 482352 215340 482354
rect 155217 482296 155222 482352
rect 155278 482296 215340 482352
rect 155217 482294 215340 482296
rect 155217 482291 155283 482294
rect 215334 482292 215340 482294
rect 215404 482292 215410 482356
rect 236545 482354 236611 482357
rect 375414 482354 375420 482356
rect 236545 482352 375420 482354
rect 236545 482296 236550 482352
rect 236606 482296 375420 482352
rect 236545 482294 375420 482296
rect 236545 482291 236611 482294
rect 375414 482292 375420 482294
rect 375484 482292 375490 482356
rect 3509 482218 3575 482221
rect 318057 482218 318123 482221
rect 3509 482216 318123 482218
rect 3509 482160 3514 482216
rect 3570 482160 318062 482216
rect 318118 482160 318123 482216
rect 3509 482158 318123 482160
rect 3509 482155 3575 482158
rect 318057 482155 318123 482158
rect 172421 480994 172487 480997
rect 202454 480994 202460 480996
rect 172421 480992 202460 480994
rect 172421 480936 172426 480992
rect 172482 480936 202460 480992
rect 172421 480934 202460 480936
rect 172421 480931 172487 480934
rect 202454 480932 202460 480934
rect 202524 480932 202530 480996
rect 154481 480858 154547 480861
rect 214046 480858 214052 480860
rect 154481 480856 214052 480858
rect 154481 480800 154486 480856
rect 154542 480800 214052 480856
rect 154481 480798 214052 480800
rect 154481 480795 154547 480798
rect 214046 480796 214052 480798
rect 214116 480796 214122 480860
rect 232129 480858 232195 480861
rect 370078 480858 370084 480860
rect 232129 480856 370084 480858
rect 232129 480800 232134 480856
rect 232190 480800 370084 480856
rect 232129 480798 370084 480800
rect 232129 480795 232195 480798
rect 370078 480796 370084 480798
rect 370148 480796 370154 480860
rect 42609 480042 42675 480045
rect 80513 480042 80579 480045
rect 42609 480040 80579 480042
rect 42609 479984 42614 480040
rect 42670 479984 80518 480040
rect 80574 479984 80579 480040
rect 42609 479982 80579 479984
rect 42609 479979 42675 479982
rect 80513 479979 80579 479982
rect 57646 479844 57652 479908
rect 57716 479906 57722 479908
rect 118693 479906 118759 479909
rect 57716 479904 118759 479906
rect 57716 479848 118698 479904
rect 118754 479848 118759 479904
rect 57716 479846 118759 479848
rect 57716 479844 57722 479846
rect 118693 479843 118759 479846
rect 50337 479770 50403 479773
rect 121913 479770 121979 479773
rect 50337 479768 121979 479770
rect 50337 479712 50342 479768
rect 50398 479712 121918 479768
rect 121974 479712 121979 479768
rect 50337 479710 121979 479712
rect 50337 479707 50403 479710
rect 121913 479707 121979 479710
rect 178677 479770 178743 479773
rect 217174 479770 217180 479772
rect 178677 479768 217180 479770
rect 178677 479712 178682 479768
rect 178738 479712 217180 479768
rect 178677 479710 217180 479712
rect 178677 479707 178743 479710
rect 217174 479708 217180 479710
rect 217244 479708 217250 479772
rect 286133 479770 286199 479773
rect 359590 479770 359596 479772
rect 286133 479768 359596 479770
rect 286133 479712 286138 479768
rect 286194 479712 359596 479768
rect 286133 479710 359596 479712
rect 286133 479707 286199 479710
rect 359590 479708 359596 479710
rect 359660 479708 359666 479772
rect 43805 479634 43871 479637
rect 118785 479634 118851 479637
rect 43805 479632 118851 479634
rect 43805 479576 43810 479632
rect 43866 479576 118790 479632
rect 118846 479576 118851 479632
rect 43805 479574 118851 479576
rect 43805 479571 43871 479574
rect 118785 479571 118851 479574
rect 146661 479634 146727 479637
rect 215886 479634 215892 479636
rect 146661 479632 215892 479634
rect 146661 479576 146666 479632
rect 146722 479576 215892 479632
rect 146661 479574 215892 479576
rect 146661 479571 146727 479574
rect 215886 479572 215892 479574
rect 215956 479572 215962 479636
rect 223665 479634 223731 479637
rect 378726 479634 378732 479636
rect 223665 479632 378732 479634
rect 223665 479576 223670 479632
rect 223726 479576 378732 479632
rect 223665 479574 378732 479576
rect 223665 479571 223731 479574
rect 378726 479572 378732 479574
rect 378796 479572 378802 479636
rect 42241 479498 42307 479501
rect 122373 479498 122439 479501
rect 42241 479496 122439 479498
rect 42241 479440 42246 479496
rect 42302 479440 122378 479496
rect 122434 479440 122439 479496
rect 42241 479438 122439 479440
rect 42241 479435 42307 479438
rect 122373 479435 122439 479438
rect 152733 479498 152799 479501
rect 208342 479498 208348 479500
rect 152733 479496 208348 479498
rect 152733 479440 152738 479496
rect 152794 479440 208348 479496
rect 152733 479438 208348 479440
rect 152733 479435 152799 479438
rect 208342 479436 208348 479438
rect 208412 479436 208418 479500
rect 210366 479436 210372 479500
rect 210436 479498 210442 479500
rect 512085 479498 512151 479501
rect 210436 479496 512151 479498
rect 210436 479440 512090 479496
rect 512146 479440 512151 479496
rect 210436 479438 512151 479440
rect 210436 479436 210442 479438
rect 512085 479435 512151 479438
rect 170305 478410 170371 478413
rect 213310 478410 213316 478412
rect 170305 478408 213316 478410
rect 170305 478352 170310 478408
rect 170366 478352 213316 478408
rect 170305 478350 213316 478352
rect 170305 478347 170371 478350
rect 213310 478348 213316 478350
rect 213380 478348 213386 478412
rect 151813 478274 151879 478277
rect 210550 478274 210556 478276
rect 151813 478272 210556 478274
rect 151813 478216 151818 478272
rect 151874 478216 210556 478272
rect 151813 478214 210556 478216
rect 151813 478211 151879 478214
rect 210550 478212 210556 478214
rect 210620 478212 210626 478276
rect 228541 478274 228607 478277
rect 358118 478274 358124 478276
rect 228541 478272 358124 478274
rect 228541 478216 228546 478272
rect 228602 478216 358124 478272
rect 228541 478214 358124 478216
rect 228541 478211 228607 478214
rect 358118 478212 358124 478214
rect 358188 478212 358194 478276
rect 147765 478138 147831 478141
rect 213126 478138 213132 478140
rect 147765 478136 213132 478138
rect 147765 478080 147770 478136
rect 147826 478080 213132 478136
rect 147765 478078 213132 478080
rect 147765 478075 147831 478078
rect 213126 478076 213132 478078
rect 213196 478076 213202 478140
rect 240317 478138 240383 478141
rect 379462 478138 379468 478140
rect 240317 478136 379468 478138
rect 240317 478080 240322 478136
rect 240378 478080 379468 478136
rect 240317 478078 379468 478080
rect 240317 478075 240383 478078
rect 379462 478076 379468 478078
rect 379532 478076 379538 478140
rect 57462 477260 57468 477324
rect 57532 477322 57538 477324
rect 128353 477322 128419 477325
rect 57532 477320 128419 477322
rect 57532 477264 128358 477320
rect 128414 477264 128419 477320
rect 57532 477262 128419 477264
rect 57532 477260 57538 477262
rect 128353 477259 128419 477262
rect 44766 477124 44772 477188
rect 44836 477186 44842 477188
rect 124213 477186 124279 477189
rect 44836 477184 124279 477186
rect 44836 477128 124218 477184
rect 124274 477128 124279 477184
rect 44836 477126 124279 477128
rect 44836 477124 44842 477126
rect 124213 477123 124279 477126
rect 44950 476988 44956 477052
rect 45020 477050 45026 477052
rect 125777 477050 125843 477053
rect 45020 477048 125843 477050
rect 45020 476992 125782 477048
rect 125838 476992 125843 477048
rect 45020 476990 125843 476992
rect 45020 476988 45026 476990
rect 125777 476987 125843 476990
rect 43529 476914 43595 476917
rect 124949 476914 125015 476917
rect 43529 476912 125015 476914
rect 43529 476856 43534 476912
rect 43590 476856 124954 476912
rect 125010 476856 125015 476912
rect 43529 476854 125015 476856
rect 43529 476851 43595 476854
rect 124949 476851 125015 476854
rect 157517 476914 157583 476917
rect 209814 476914 209820 476916
rect 157517 476912 209820 476914
rect 157517 476856 157522 476912
rect 157578 476856 209820 476912
rect 157517 476854 209820 476856
rect 157517 476851 157583 476854
rect 209814 476852 209820 476854
rect 209884 476852 209890 476916
rect 42333 476778 42399 476781
rect 124489 476778 124555 476781
rect 42333 476776 124555 476778
rect 42333 476720 42338 476776
rect 42394 476720 124494 476776
rect 124550 476720 124555 476776
rect 42333 476718 124555 476720
rect 42333 476715 42399 476718
rect 124489 476715 124555 476718
rect 151353 476778 151419 476781
rect 214414 476778 214420 476780
rect 151353 476776 214420 476778
rect 151353 476720 151358 476776
rect 151414 476720 214420 476776
rect 151353 476718 214420 476720
rect 151353 476715 151419 476718
rect 214414 476716 214420 476718
rect 214484 476716 214490 476780
rect 234613 476778 234679 476781
rect 378174 476778 378180 476780
rect 234613 476776 378180 476778
rect 234613 476720 234618 476776
rect 234674 476720 378180 476776
rect 234613 476718 378180 476720
rect 234613 476715 234679 476718
rect 378174 476716 378180 476718
rect 378244 476716 378250 476780
rect -960 475540 480 475780
rect 270493 475690 270559 475693
rect 359774 475690 359780 475692
rect 270493 475688 359780 475690
rect 270493 475632 270498 475688
rect 270554 475632 359780 475688
rect 270493 475630 359780 475632
rect 270493 475627 270559 475630
rect 359774 475628 359780 475630
rect 359844 475628 359850 475692
rect 156781 475554 156847 475557
rect 218646 475554 218652 475556
rect 156781 475552 218652 475554
rect 156781 475496 156786 475552
rect 156842 475496 218652 475552
rect 156781 475494 218652 475496
rect 156781 475491 156847 475494
rect 218646 475492 218652 475494
rect 218716 475492 218722 475556
rect 232405 475554 232471 475557
rect 360142 475554 360148 475556
rect 232405 475552 360148 475554
rect 232405 475496 232410 475552
rect 232466 475496 360148 475552
rect 232405 475494 360148 475496
rect 232405 475491 232471 475494
rect 360142 475492 360148 475494
rect 360212 475492 360218 475556
rect 202086 475356 202092 475420
rect 202156 475418 202162 475420
rect 483013 475418 483079 475421
rect 202156 475416 483079 475418
rect 202156 475360 483018 475416
rect 483074 475360 483079 475416
rect 202156 475358 483079 475360
rect 202156 475356 202162 475358
rect 483013 475355 483079 475358
rect 155953 474194 156019 474197
rect 207054 474194 207060 474196
rect 155953 474192 207060 474194
rect 155953 474136 155958 474192
rect 156014 474136 207060 474192
rect 155953 474134 207060 474136
rect 155953 474131 156019 474134
rect 207054 474132 207060 474134
rect 207124 474132 207130 474196
rect 150433 474058 150499 474061
rect 216070 474058 216076 474060
rect 150433 474056 216076 474058
rect 150433 474000 150438 474056
rect 150494 474000 216076 474056
rect 150433 473998 216076 474000
rect 150433 473995 150499 473998
rect 216070 473996 216076 473998
rect 216140 473996 216146 474060
rect 223573 474058 223639 474061
rect 378910 474058 378916 474060
rect 223573 474056 378916 474058
rect 223573 474000 223578 474056
rect 223634 474000 378916 474056
rect 223573 473998 378916 474000
rect 223573 473995 223639 473998
rect 378910 473996 378916 473998
rect 378980 473996 378986 474060
rect 252645 472970 252711 472973
rect 377254 472970 377260 472972
rect 252645 472968 377260 472970
rect 252645 472912 252650 472968
rect 252706 472912 377260 472968
rect 252645 472910 377260 472912
rect 252645 472907 252711 472910
rect 377254 472908 377260 472910
rect 377324 472908 377330 472972
rect 169845 472834 169911 472837
rect 216254 472834 216260 472836
rect 169845 472832 216260 472834
rect 169845 472776 169850 472832
rect 169906 472776 216260 472832
rect 169845 472774 216260 472776
rect 169845 472771 169911 472774
rect 216254 472772 216260 472774
rect 216324 472772 216330 472836
rect 366950 472772 366956 472836
rect 367020 472834 367026 472836
rect 506606 472834 506612 472836
rect 367020 472774 506612 472834
rect 367020 472772 367026 472774
rect 506606 472772 506612 472774
rect 506676 472772 506682 472836
rect 147673 472698 147739 472701
rect 202270 472698 202276 472700
rect 147673 472696 202276 472698
rect 147673 472640 147678 472696
rect 147734 472640 202276 472696
rect 147673 472638 202276 472640
rect 147673 472635 147739 472638
rect 202270 472636 202276 472638
rect 202340 472636 202346 472700
rect 226333 472698 226399 472701
rect 371918 472698 371924 472700
rect 226333 472696 371924 472698
rect 226333 472640 226338 472696
rect 226394 472640 371924 472696
rect 226333 472638 371924 472640
rect 226333 472635 226399 472638
rect 371918 472636 371924 472638
rect 371988 472636 371994 472700
rect 145741 472562 145807 472565
rect 203190 472562 203196 472564
rect 145741 472560 203196 472562
rect 145741 472504 145746 472560
rect 145802 472504 203196 472560
rect 145741 472502 203196 472504
rect 145741 472499 145807 472502
rect 203190 472500 203196 472502
rect 203260 472500 203266 472564
rect 229093 472562 229159 472565
rect 379094 472562 379100 472564
rect 229093 472560 379100 472562
rect 229093 472504 229098 472560
rect 229154 472504 379100 472560
rect 229093 472502 379100 472504
rect 229093 472499 229159 472502
rect 379094 472500 379100 472502
rect 379164 472500 379170 472564
rect 174813 471746 174879 471749
rect 199510 471746 199516 471748
rect 174813 471744 199516 471746
rect 174813 471688 174818 471744
rect 174874 471688 199516 471744
rect 174813 471686 199516 471688
rect 174813 471683 174879 471686
rect 199510 471684 199516 471686
rect 199580 471684 199586 471748
rect 53557 471610 53623 471613
rect 84285 471610 84351 471613
rect 53557 471608 84351 471610
rect 53557 471552 53562 471608
rect 53618 471552 84290 471608
rect 84346 471552 84351 471608
rect 53557 471550 84351 471552
rect 53557 471547 53623 471550
rect 84285 471547 84351 471550
rect 171225 471610 171291 471613
rect 204846 471610 204852 471612
rect 171225 471608 204852 471610
rect 171225 471552 171230 471608
rect 171286 471552 204852 471608
rect 171225 471550 204852 471552
rect 171225 471547 171291 471550
rect 204846 471548 204852 471550
rect 204916 471548 204922 471612
rect 56317 471474 56383 471477
rect 88517 471474 88583 471477
rect 56317 471472 88583 471474
rect 56317 471416 56322 471472
rect 56378 471416 88522 471472
rect 88578 471416 88583 471472
rect 56317 471414 88583 471416
rect 56317 471411 56383 471414
rect 88517 471411 88583 471414
rect 182265 471474 182331 471477
rect 217358 471474 217364 471476
rect 182265 471472 217364 471474
rect 182265 471416 182270 471472
rect 182326 471416 217364 471472
rect 182265 471414 217364 471416
rect 182265 471411 182331 471414
rect 217358 471412 217364 471414
rect 217428 471412 217434 471476
rect 53649 471338 53715 471341
rect 85757 471338 85823 471341
rect 53649 471336 85823 471338
rect 53649 471280 53654 471336
rect 53710 471280 85762 471336
rect 85818 471280 85823 471336
rect 53649 471278 85823 471280
rect 53649 471275 53715 471278
rect 85757 471275 85823 471278
rect 172697 471338 172763 471341
rect 211981 471338 212047 471341
rect 172697 471336 212047 471338
rect 172697 471280 172702 471336
rect 172758 471280 211986 471336
rect 212042 471280 212047 471336
rect 172697 471278 212047 471280
rect 172697 471275 172763 471278
rect 211981 471275 212047 471278
rect 296805 471338 296871 471341
rect 377438 471338 377444 471340
rect 296805 471336 377444 471338
rect 296805 471280 296810 471336
rect 296866 471280 377444 471336
rect 296805 471278 377444 471280
rect 296805 471275 296871 471278
rect 377438 471276 377444 471278
rect 377508 471276 377514 471340
rect 583520 471324 584960 471564
rect 55029 471202 55095 471205
rect 88425 471202 88491 471205
rect 55029 471200 88491 471202
rect 55029 471144 55034 471200
rect 55090 471144 88430 471200
rect 88486 471144 88491 471200
rect 55029 471142 88491 471144
rect 55029 471139 55095 471142
rect 88425 471139 88491 471142
rect 162485 471202 162551 471205
rect 203609 471202 203675 471205
rect 162485 471200 203675 471202
rect 162485 471144 162490 471200
rect 162546 471144 203614 471200
rect 203670 471144 203675 471200
rect 162485 471142 203675 471144
rect 162485 471139 162551 471142
rect 203609 471139 203675 471142
rect 295517 471202 295583 471205
rect 377622 471202 377628 471204
rect 295517 471200 377628 471202
rect 295517 471144 295522 471200
rect 295578 471144 377628 471200
rect 295517 471142 377628 471144
rect 295517 471139 295583 471142
rect 377622 471140 377628 471142
rect 377692 471140 377698 471204
rect 47894 469780 47900 469844
rect 47964 469842 47970 469844
rect 81525 469842 81591 469845
rect 47964 469840 81591 469842
rect 47964 469784 81530 469840
rect 81586 469784 81591 469840
rect 47964 469782 81591 469784
rect 47964 469780 47970 469782
rect 81525 469779 81591 469782
rect 60222 469100 60228 469164
rect 60292 469162 60298 469164
rect 73153 469162 73219 469165
rect 60292 469160 73219 469162
rect 60292 469104 73158 469160
rect 73214 469104 73219 469160
rect 60292 469102 73219 469104
rect 60292 469100 60298 469102
rect 73153 469099 73219 469102
rect 48078 468964 48084 469028
rect 48148 469026 48154 469028
rect 69105 469026 69171 469029
rect 48148 469024 69171 469026
rect 48148 468968 69110 469024
rect 69166 468968 69171 469024
rect 48148 468966 69171 468968
rect 48148 468964 48154 468966
rect 69105 468963 69171 468966
rect 171133 469026 171199 469029
rect 206318 469026 206324 469028
rect 171133 469024 206324 469026
rect 171133 468968 171138 469024
rect 171194 468968 206324 469024
rect 171133 468966 206324 468968
rect 171133 468963 171199 468966
rect 206318 468964 206324 468966
rect 206388 468964 206394 469028
rect 46606 468828 46612 468892
rect 46676 468890 46682 468892
rect 69197 468890 69263 468893
rect 46676 468888 69263 468890
rect 46676 468832 69202 468888
rect 69258 468832 69263 468888
rect 46676 468830 69263 468832
rect 46676 468828 46682 468830
rect 69197 468827 69263 468830
rect 169753 468890 169819 468893
rect 205030 468890 205036 468892
rect 169753 468888 205036 468890
rect 169753 468832 169758 468888
rect 169814 468832 205036 468888
rect 169753 468830 205036 468832
rect 169753 468827 169819 468830
rect 205030 468828 205036 468830
rect 205100 468828 205106 468892
rect 55438 468692 55444 468756
rect 55508 468754 55514 468756
rect 78673 468754 78739 468757
rect 55508 468752 78739 468754
rect 55508 468696 78678 468752
rect 78734 468696 78739 468752
rect 55508 468694 78739 468696
rect 55508 468692 55514 468694
rect 78673 468691 78739 468694
rect 160093 468754 160159 468757
rect 200982 468754 200988 468756
rect 160093 468752 200988 468754
rect 160093 468696 160098 468752
rect 160154 468696 200988 468752
rect 160093 468694 200988 468696
rect 160093 468691 160159 468694
rect 200982 468692 200988 468694
rect 201052 468692 201058 468756
rect 53598 468556 53604 468620
rect 53668 468618 53674 468620
rect 78857 468618 78923 468621
rect 53668 468616 78923 468618
rect 53668 468560 78862 468616
rect 78918 468560 78923 468616
rect 53668 468558 78923 468560
rect 53668 468556 53674 468558
rect 78857 468555 78923 468558
rect 161473 468618 161539 468621
rect 206502 468618 206508 468620
rect 161473 468616 206508 468618
rect 161473 468560 161478 468616
rect 161534 468560 206508 468616
rect 161473 468558 206508 468560
rect 161473 468555 161539 468558
rect 206502 468556 206508 468558
rect 206572 468556 206578 468620
rect 50470 468420 50476 468484
rect 50540 468482 50546 468484
rect 94037 468482 94103 468485
rect 50540 468480 94103 468482
rect 50540 468424 94042 468480
rect 94098 468424 94103 468480
rect 50540 468422 94103 468424
rect 50540 468420 50546 468422
rect 94037 468419 94103 468422
rect 168373 468482 168439 468485
rect 213494 468482 213500 468484
rect 168373 468480 213500 468482
rect 168373 468424 168378 468480
rect 168434 468424 213500 468480
rect 168373 468422 213500 468424
rect 168373 468419 168439 468422
rect 213494 468420 213500 468422
rect 213564 468420 213570 468484
rect 296713 468482 296779 468485
rect 377806 468482 377812 468484
rect 296713 468480 377812 468482
rect 296713 468424 296718 468480
rect 296774 468424 377812 468480
rect 296713 468422 377812 468424
rect 296713 468419 296779 468422
rect 377806 468420 377812 468422
rect 377876 468420 377882 468484
rect 58934 468284 58940 468348
rect 59004 468346 59010 468348
rect 67817 468346 67883 468349
rect 59004 468344 67883 468346
rect 59004 468288 67822 468344
rect 67878 468288 67883 468344
rect 59004 468286 67883 468288
rect 59004 468284 59010 468286
rect 67817 468283 67883 468286
rect 48630 467876 48636 467940
rect 48700 467938 48706 467940
rect 49509 467938 49575 467941
rect 50705 467940 50771 467941
rect 50654 467938 50660 467940
rect 48700 467936 49575 467938
rect 48700 467880 49514 467936
rect 49570 467880 49575 467936
rect 48700 467878 49575 467880
rect 50614 467878 50660 467938
rect 50724 467936 50771 467940
rect 50766 467880 50771 467936
rect 48700 467876 48706 467878
rect 49509 467875 49575 467878
rect 50654 467876 50660 467878
rect 50724 467876 50771 467880
rect 50705 467875 50771 467876
rect 44081 467258 44147 467261
rect 71865 467258 71931 467261
rect 44081 467256 71931 467258
rect 44081 467200 44086 467256
rect 44142 467200 71870 467256
rect 71926 467200 71931 467256
rect 44081 467198 71931 467200
rect 44081 467195 44147 467198
rect 71865 467195 71931 467198
rect 172605 467258 172671 467261
rect 208894 467258 208900 467260
rect 172605 467256 208900 467258
rect 172605 467200 172610 467256
rect 172666 467200 208900 467256
rect 172605 467198 208900 467200
rect 172605 467195 172671 467198
rect 208894 467196 208900 467198
rect 208964 467196 208970 467260
rect 42701 467122 42767 467125
rect 70485 467122 70551 467125
rect 42701 467120 70551 467122
rect 42701 467064 42706 467120
rect 42762 467064 70490 467120
rect 70546 467064 70551 467120
rect 42701 467062 70551 467064
rect 42701 467059 42767 467062
rect 70485 467059 70551 467062
rect 153193 467122 153259 467125
rect 218830 467122 218836 467124
rect 153193 467120 218836 467122
rect 153193 467064 153198 467120
rect 153254 467064 218836 467120
rect 153193 467062 218836 467064
rect 153193 467059 153259 467062
rect 218830 467060 218836 467062
rect 218900 467060 218906 467124
rect 179638 466924 179644 466988
rect 179708 466986 179714 466988
rect 180149 466986 180215 466989
rect 179708 466984 180215 466986
rect 179708 466928 180154 466984
rect 180210 466928 180215 466984
rect 179708 466926 180215 466928
rect 179708 466924 179714 466926
rect 180149 466923 180215 466926
rect 178033 466578 178099 466581
rect 190913 466580 190979 466581
rect 338481 466580 338547 466581
rect 339769 466580 339835 466581
rect 350993 466580 351059 466581
rect 178350 466578 178356 466580
rect 178033 466576 178356 466578
rect 178033 466520 178038 466576
rect 178094 466520 178356 466576
rect 178033 466518 178356 466520
rect 178033 466515 178099 466518
rect 178350 466516 178356 466518
rect 178420 466516 178426 466580
rect 190862 466578 190868 466580
rect 190822 466518 190868 466578
rect 190932 466576 190979 466580
rect 338430 466578 338436 466580
rect 190974 466520 190979 466576
rect 190862 466516 190868 466518
rect 190932 466516 190979 466520
rect 338390 466518 338436 466578
rect 338500 466576 338547 466580
rect 339718 466578 339724 466580
rect 338542 466520 338547 466576
rect 338430 466516 338436 466518
rect 338500 466516 338547 466520
rect 339678 466518 339724 466578
rect 339788 466576 339835 466580
rect 350942 466578 350948 466580
rect 339830 466520 339835 466576
rect 339718 466516 339724 466518
rect 339788 466516 339835 466520
rect 350902 466518 350948 466578
rect 351012 466576 351059 466580
rect 351054 466520 351059 466576
rect 350942 466516 350948 466518
rect 351012 466516 351059 466520
rect 190913 466515 190979 466516
rect 338481 466515 338547 466516
rect 339769 466515 339835 466516
rect 350993 466515 351059 466516
rect 498469 466580 498535 466581
rect 499757 466580 499823 466581
rect 510889 466580 510955 466581
rect 498469 466576 498516 466580
rect 498580 466578 498586 466580
rect 498469 466520 498474 466576
rect 498469 466516 498516 466520
rect 498580 466518 498626 466578
rect 499757 466576 499804 466580
rect 499868 466578 499874 466580
rect 510838 466578 510844 466580
rect 499757 466520 499762 466576
rect 498580 466516 498586 466518
rect 499757 466516 499804 466520
rect 499868 466518 499914 466578
rect 510798 466518 510844 466578
rect 510908 466576 510955 466580
rect 510950 466520 510955 466576
rect 499868 466516 499874 466518
rect 510838 466516 510844 466518
rect 510908 466516 510955 466520
rect 498469 466515 498535 466516
rect 499757 466515 499823 466516
rect 510889 466515 510955 466516
rect 58566 466380 58572 466444
rect 58636 466442 58642 466444
rect 69013 466442 69079 466445
rect 58636 466440 69079 466442
rect 58636 466384 69018 466440
rect 69074 466384 69079 466440
rect 58636 466382 69079 466384
rect 58636 466380 58642 466382
rect 69013 466379 69079 466382
rect 54886 466244 54892 466308
rect 54956 466306 54962 466308
rect 71773 466306 71839 466309
rect 54956 466304 71839 466306
rect 54956 466248 71778 466304
rect 71834 466248 71839 466304
rect 54956 466246 71839 466248
rect 54956 466244 54962 466246
rect 71773 466243 71839 466246
rect 53414 466108 53420 466172
rect 53484 466170 53490 466172
rect 74625 466170 74691 466173
rect 53484 466168 74691 466170
rect 53484 466112 74630 466168
rect 74686 466112 74691 466168
rect 53484 466110 74691 466112
rect 53484 466108 53490 466110
rect 74625 466107 74691 466110
rect 170397 466170 170463 466173
rect 198774 466170 198780 466172
rect 170397 466168 198780 466170
rect 170397 466112 170402 466168
rect 170458 466112 198780 466168
rect 170397 466110 198780 466112
rect 170397 466107 170463 466110
rect 198774 466108 198780 466110
rect 198844 466108 198850 466172
rect 54702 465972 54708 466036
rect 54772 466034 54778 466036
rect 76005 466034 76071 466037
rect 54772 466032 76071 466034
rect 54772 465976 76010 466032
rect 76066 465976 76071 466032
rect 54772 465974 76071 465976
rect 54772 465972 54778 465974
rect 76005 465971 76071 465974
rect 165613 466034 165679 466037
rect 203701 466034 203767 466037
rect 165613 466032 203767 466034
rect 165613 465976 165618 466032
rect 165674 465976 203706 466032
rect 203762 465976 203767 466032
rect 165613 465974 203767 465976
rect 165613 465971 165679 465974
rect 203701 465971 203767 465974
rect 51574 465836 51580 465900
rect 51644 465898 51650 465900
rect 51993 465898 52059 465901
rect 51644 465896 52059 465898
rect 51644 465840 51998 465896
rect 52054 465840 52059 465896
rect 51644 465838 52059 465840
rect 51644 465836 51650 465838
rect 51993 465835 52059 465838
rect 53046 465836 53052 465900
rect 53116 465898 53122 465900
rect 74533 465898 74599 465901
rect 53116 465896 74599 465898
rect 53116 465840 74538 465896
rect 74594 465840 74599 465896
rect 53116 465838 74599 465840
rect 53116 465836 53122 465838
rect 74533 465835 74599 465838
rect 166993 465898 167059 465901
rect 207974 465898 207980 465900
rect 166993 465896 207980 465898
rect 166993 465840 166998 465896
rect 167054 465840 207980 465896
rect 166993 465838 207980 465840
rect 166993 465835 167059 465838
rect 207974 465836 207980 465838
rect 208044 465836 208050 465900
rect 277393 465898 277459 465901
rect 359958 465898 359964 465900
rect 277393 465896 359964 465898
rect 277393 465840 277398 465896
rect 277454 465840 359964 465896
rect 277393 465838 359964 465840
rect 277393 465835 277459 465838
rect 359958 465836 359964 465838
rect 360028 465836 360034 465900
rect 52126 465700 52132 465764
rect 52196 465762 52202 465764
rect 74717 465762 74783 465765
rect 52196 465760 74783 465762
rect 52196 465704 74722 465760
rect 74778 465704 74783 465760
rect 52196 465702 74783 465704
rect 52196 465700 52202 465702
rect 74717 465699 74783 465702
rect 162853 465762 162919 465765
rect 216029 465762 216095 465765
rect 162853 465760 216095 465762
rect 162853 465704 162858 465760
rect 162914 465704 216034 465760
rect 216090 465704 216095 465760
rect 162853 465702 216095 465704
rect 162853 465699 162919 465702
rect 216029 465699 216095 465702
rect 248413 465762 248479 465765
rect 370630 465762 370636 465764
rect 248413 465760 370636 465762
rect 248413 465704 248418 465760
rect 248474 465704 370636 465760
rect 248413 465702 370636 465704
rect 248413 465699 248479 465702
rect 370630 465700 370636 465702
rect 370700 465700 370706 465764
rect 58750 465564 58756 465628
rect 58820 465626 58826 465628
rect 67633 465626 67699 465629
rect 58820 465624 67699 465626
rect 58820 465568 67638 465624
rect 67694 465568 67699 465624
rect 58820 465566 67699 465568
rect 58820 465564 58826 465566
rect 67633 465563 67699 465566
rect 51758 465156 51764 465220
rect 51828 465218 51834 465220
rect 52269 465218 52335 465221
rect 51828 465216 52335 465218
rect 51828 465160 52274 465216
rect 52330 465160 52335 465216
rect 51828 465158 52335 465160
rect 51828 465156 51834 465158
rect 52269 465155 52335 465158
rect 187693 464402 187759 464405
rect 199142 464402 199148 464404
rect 187693 464400 199148 464402
rect 187693 464344 187698 464400
rect 187754 464344 199148 464400
rect 187693 464342 199148 464344
rect 187693 464339 187759 464342
rect 199142 464340 199148 464342
rect 199212 464340 199218 464404
rect -960 462634 480 462724
rect 3785 462634 3851 462637
rect -960 462632 3851 462634
rect -960 462576 3790 462632
rect 3846 462576 3851 462632
rect -960 462574 3851 462576
rect -960 462484 480 462574
rect 3785 462571 3851 462574
rect 196558 460186 196618 460190
rect 199009 460186 199075 460189
rect 196558 460184 199075 460186
rect 196558 460128 199014 460184
rect 199070 460128 199075 460184
rect 196558 460126 199075 460128
rect 356562 460186 356622 460190
rect 358905 460186 358971 460189
rect 356562 460184 358971 460186
rect 356562 460128 358910 460184
rect 358966 460128 358971 460184
rect 356562 460126 358971 460128
rect 199009 460123 199075 460126
rect 358905 460123 358971 460126
rect 516558 459642 516618 460190
rect 518893 459642 518959 459645
rect 519445 459642 519511 459645
rect 516558 459640 519511 459642
rect 516558 459584 518898 459640
rect 518954 459584 519450 459640
rect 519506 459584 519511 459640
rect 516558 459582 519511 459584
rect 518893 459579 518959 459582
rect 519445 459579 519511 459582
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 57053 417890 57119 417893
rect 60002 417890 60062 417894
rect 57053 417888 60062 417890
rect 57053 417832 57058 417888
rect 57114 417832 60062 417888
rect 57053 417830 60062 417832
rect 216673 417890 216739 417893
rect 217869 417890 217935 417893
rect 219390 417890 220064 417924
rect 216673 417888 220064 417890
rect 216673 417832 216678 417888
rect 216734 417832 217874 417888
rect 217930 417864 220064 417888
rect 377765 417890 377831 417893
rect 379470 417890 380052 417924
rect 377765 417888 380052 417890
rect 217930 417832 219450 417864
rect 216673 417830 219450 417832
rect 377765 417832 377770 417888
rect 377826 417864 380052 417888
rect 377826 417832 379530 417864
rect 377765 417830 379530 417832
rect 57053 417827 57119 417830
rect 216673 417827 216739 417830
rect 217869 417827 217935 417830
rect 377765 417827 377831 417830
rect 57237 416938 57303 416941
rect 60002 416938 60062 416942
rect 57237 416936 60062 416938
rect 57237 416880 57242 416936
rect 57298 416880 60062 416936
rect 57237 416878 60062 416880
rect 217225 416938 217291 416941
rect 219390 416938 220064 416972
rect 217225 416936 220064 416938
rect 217225 416880 217230 416936
rect 217286 416912 220064 416936
rect 377213 416938 377279 416941
rect 377949 416938 378015 416941
rect 379470 416938 380052 416972
rect 377213 416936 380052 416938
rect 217286 416880 219450 416912
rect 217225 416878 219450 416880
rect 377213 416880 377218 416936
rect 377274 416880 377954 416936
rect 378010 416912 380052 416936
rect 378010 416880 379530 416912
rect 377213 416878 379530 416880
rect 57237 416875 57303 416878
rect 217225 416875 217291 416878
rect 377213 416875 377279 416878
rect 377949 416875 378015 416878
rect 206686 415244 206692 415308
rect 206756 415306 206762 415308
rect 206921 415306 206987 415309
rect 206756 415304 206987 415306
rect 206756 415248 206926 415304
rect 206982 415248 206987 415304
rect 206756 415246 206987 415248
rect 206756 415244 206762 415246
rect 206921 415243 206987 415246
rect 376937 415306 377003 415309
rect 377397 415306 377463 415309
rect 376937 415304 377463 415306
rect 376937 415248 376942 415304
rect 376998 415248 377402 415304
rect 377458 415248 377463 415304
rect 376937 415246 377463 415248
rect 376937 415243 377003 415246
rect 377397 415243 377463 415246
rect 57053 414218 57119 414221
rect 60002 414218 60062 414766
rect 217133 414762 217199 414765
rect 219390 414762 220064 414796
rect 217133 414760 220064 414762
rect 217133 414704 217138 414760
rect 217194 414736 220064 414760
rect 376937 414762 377003 414765
rect 379470 414762 380052 414796
rect 376937 414760 380052 414762
rect 217194 414704 219450 414736
rect 217133 414702 219450 414704
rect 376937 414704 376942 414760
rect 376998 414736 380052 414760
rect 376998 414704 379530 414736
rect 376937 414702 379530 414704
rect 217133 414699 217199 414702
rect 376937 414699 377003 414702
rect 57053 414216 60062 414218
rect 57053 414160 57058 414216
rect 57114 414160 60062 414216
rect 57053 414158 60062 414160
rect 57053 414155 57119 414158
rect 377581 413946 377647 413949
rect 377857 413946 377923 413949
rect 377581 413944 379530 413946
rect 377581 413888 377586 413944
rect 377642 413888 377862 413944
rect 377918 413888 379530 413944
rect 377581 413886 379530 413888
rect 377581 413883 377647 413886
rect 377857 413883 377923 413886
rect 379470 413844 379530 413886
rect 57237 413266 57303 413269
rect 60002 413266 60062 413814
rect 216857 413810 216923 413813
rect 219390 413810 220064 413844
rect 216857 413808 220064 413810
rect 216857 413752 216862 413808
rect 216918 413784 220064 413808
rect 379470 413784 380052 413844
rect 216918 413752 219450 413784
rect 216857 413750 219450 413752
rect 216857 413747 216923 413750
rect 57237 413264 60062 413266
rect 57237 413208 57242 413264
rect 57298 413208 60062 413264
rect 57237 413206 60062 413208
rect 57237 413203 57303 413206
rect 57237 411498 57303 411501
rect 60002 411498 60062 412046
rect 217317 412042 217383 412045
rect 219390 412042 220064 412076
rect 217317 412040 220064 412042
rect 217317 411984 217322 412040
rect 217378 412016 220064 412040
rect 377213 412042 377279 412045
rect 377581 412042 377647 412045
rect 379470 412042 380052 412076
rect 377213 412040 380052 412042
rect 217378 411984 219450 412016
rect 217317 411982 219450 411984
rect 377213 411984 377218 412040
rect 377274 411984 377586 412040
rect 377642 412016 380052 412040
rect 377642 411984 379530 412016
rect 377213 411982 379530 411984
rect 217317 411979 217383 411982
rect 377213 411979 377279 411982
rect 377581 411979 377647 411982
rect 57237 411496 60062 411498
rect 57237 411440 57242 411496
rect 57298 411440 60062 411496
rect 57237 411438 60062 411440
rect 57237 411435 57303 411438
rect 217317 411362 217383 411365
rect 217777 411362 217843 411365
rect 217317 411360 217843 411362
rect 217317 411304 217322 411360
rect 217378 411304 217782 411360
rect 217838 411304 217843 411360
rect 217317 411302 217843 411304
rect 217317 411299 217383 411302
rect 217777 411299 217843 411302
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 56685 410410 56751 410413
rect 60002 410410 60062 410958
rect 216673 410954 216739 410957
rect 219390 410954 220064 410988
rect 216673 410952 220064 410954
rect 216673 410896 216678 410952
rect 216734 410928 220064 410952
rect 377213 410954 377279 410957
rect 379470 410954 380052 410988
rect 377213 410952 380052 410954
rect 216734 410896 219450 410928
rect 216673 410894 219450 410896
rect 377213 410896 377218 410952
rect 377274 410928 380052 410952
rect 377274 410896 379530 410928
rect 377213 410894 379530 410896
rect 216673 410891 216739 410894
rect 377213 410891 377279 410894
rect 56685 410408 60062 410410
rect 56685 410352 56690 410408
rect 56746 410352 60062 410408
rect 56685 410350 60062 410352
rect 56685 410347 56751 410350
rect 57237 408642 57303 408645
rect 60002 408642 60062 409190
rect 216673 409186 216739 409189
rect 216949 409186 217015 409189
rect 219390 409186 220064 409220
rect 216673 409184 220064 409186
rect 216673 409128 216678 409184
rect 216734 409128 216954 409184
rect 217010 409160 220064 409184
rect 377397 409186 377463 409189
rect 378041 409186 378107 409189
rect 379470 409186 380052 409220
rect 377397 409184 380052 409186
rect 217010 409128 219450 409160
rect 216673 409126 219450 409128
rect 377397 409128 377402 409184
rect 377458 409128 378046 409184
rect 378102 409160 380052 409184
rect 378102 409128 379530 409160
rect 377397 409126 379530 409128
rect 216673 409123 216739 409126
rect 216949 409123 217015 409126
rect 377397 409123 377463 409126
rect 378041 409123 378107 409126
rect 57237 408640 60062 408642
rect 57237 408584 57242 408640
rect 57298 408584 60062 408640
rect 57237 408582 60062 408584
rect 57237 408579 57303 408582
rect 580349 404970 580415 404973
rect 583520 404970 584960 405060
rect 580349 404968 584960 404970
rect 580349 404912 580354 404968
rect 580410 404912 584960 404968
rect 580349 404910 584960 404912
rect 580349 404907 580415 404910
rect 583520 404820 584960 404910
rect 198825 400890 198891 400893
rect 196558 400888 198891 400890
rect 196558 400832 198830 400888
rect 198886 400832 198891 400888
rect 196558 400830 198891 400832
rect 196558 400350 196618 400830
rect 198825 400827 198891 400830
rect 356562 400346 356622 400350
rect 358997 400346 359063 400349
rect 356562 400344 359063 400346
rect 356562 400288 359002 400344
rect 359058 400288 359063 400344
rect 356562 400286 359063 400288
rect 516558 400346 516618 400350
rect 519077 400346 519143 400349
rect 516558 400344 519143 400346
rect 516558 400288 519082 400344
rect 519138 400288 519143 400344
rect 516558 400286 519143 400288
rect 358997 400283 359063 400286
rect 519077 400283 519143 400286
rect 196558 398170 196618 398718
rect 199469 398170 199535 398173
rect 196558 398168 199535 398170
rect 196558 398112 199474 398168
rect 199530 398112 199535 398168
rect 196558 398110 199535 398112
rect 356562 398170 356622 398718
rect 359089 398170 359155 398173
rect 356562 398168 359155 398170
rect 356562 398112 359094 398168
rect 359150 398112 359155 398168
rect 356562 398110 359155 398112
rect 516558 398170 516618 398718
rect 518985 398170 519051 398173
rect 516558 398168 519051 398170
rect 516558 398112 518990 398168
rect 519046 398112 519051 398168
rect 516558 398110 519051 398112
rect 199469 398107 199535 398110
rect 359089 398107 359155 398110
rect 518985 398107 519051 398110
rect -960 397340 480 397580
rect 196558 397354 196618 397358
rect 199377 397354 199443 397357
rect 199837 397354 199903 397357
rect 196558 397352 199903 397354
rect 196558 397296 199382 397352
rect 199438 397296 199842 397352
rect 199898 397296 199903 397352
rect 196558 397294 199903 397296
rect 199377 397291 199443 397294
rect 199837 397291 199903 397294
rect 356562 396810 356622 397358
rect 359733 396810 359799 396813
rect 356562 396808 359799 396810
rect 356562 396752 359738 396808
rect 359794 396752 359799 396808
rect 356562 396750 359799 396752
rect 516558 396810 516618 397358
rect 519353 396810 519419 396813
rect 516558 396808 519419 396810
rect 516558 396752 519358 396808
rect 519414 396752 519419 396808
rect 516558 396750 519419 396752
rect 359733 396747 359799 396750
rect 519353 396747 519419 396750
rect 196558 395314 196618 395862
rect 199561 395314 199627 395317
rect 196558 395312 199627 395314
rect 196558 395256 199566 395312
rect 199622 395256 199627 395312
rect 196558 395254 199627 395256
rect 356562 395314 356622 395862
rect 359181 395314 359247 395317
rect 356562 395312 359247 395314
rect 356562 395256 359186 395312
rect 359242 395256 359247 395312
rect 356562 395254 359247 395256
rect 516558 395314 516618 395862
rect 519169 395314 519235 395317
rect 516558 395312 519235 395314
rect 516558 395256 519174 395312
rect 519230 395256 519235 395312
rect 516558 395254 519235 395256
rect 199561 395251 199627 395254
rect 359181 395251 359247 395254
rect 519169 395251 519235 395254
rect 196558 394634 196618 394638
rect 199285 394634 199351 394637
rect 196558 394632 199351 394634
rect 196558 394576 199290 394632
rect 199346 394576 199351 394632
rect 196558 394574 199351 394576
rect 199285 394571 199351 394574
rect 356562 394090 356622 394638
rect 359273 394090 359339 394093
rect 356562 394088 359339 394090
rect 356562 394032 359278 394088
rect 359334 394032 359339 394088
rect 356562 394030 359339 394032
rect 516558 394090 516618 394638
rect 519261 394090 519327 394093
rect 516558 394088 519327 394090
rect 516558 394032 519266 394088
rect 519322 394032 519327 394088
rect 516558 394030 519327 394032
rect 359273 394027 359339 394030
rect 519261 394027 519327 394030
rect 57237 391642 57303 391645
rect 57237 391640 60062 391642
rect 57237 391584 57242 391640
rect 57298 391584 60062 391640
rect 583520 391628 584960 391868
rect 57237 391582 60062 391584
rect 57237 391579 57303 391582
rect 60002 390966 60062 391582
rect 216673 390962 216739 390965
rect 219390 390962 220064 390996
rect 216673 390960 220064 390962
rect 216673 390904 216678 390960
rect 216734 390936 220064 390960
rect 376937 390962 377003 390965
rect 379470 390962 380052 390996
rect 376937 390960 380052 390962
rect 216734 390904 219450 390936
rect 216673 390902 219450 390904
rect 376937 390904 376942 390960
rect 376998 390936 380052 390960
rect 376998 390904 379530 390936
rect 376937 390902 379530 390904
rect 216673 390899 216739 390902
rect 376937 390899 377003 390902
rect 57513 389330 57579 389333
rect 59494 389330 60032 389364
rect 57513 389328 60032 389330
rect 57513 389272 57518 389328
rect 57574 389304 60032 389328
rect 216673 389330 216739 389333
rect 219390 389330 220064 389364
rect 216673 389328 220064 389330
rect 57574 389272 59554 389304
rect 57513 389270 59554 389272
rect 216673 389272 216678 389328
rect 216734 389304 220064 389328
rect 376937 389330 377003 389333
rect 379470 389330 380052 389364
rect 376937 389328 380052 389330
rect 216734 389272 219450 389304
rect 216673 389270 219450 389272
rect 376937 389272 376942 389328
rect 376998 389304 380052 389328
rect 376998 389272 379530 389304
rect 376937 389270 379530 389272
rect 57513 389267 57579 389270
rect 216673 389267 216739 389270
rect 376937 389267 377003 389270
rect 57145 389058 57211 389061
rect 60002 389058 60062 389062
rect 57145 389056 60062 389058
rect 57145 389000 57150 389056
rect 57206 389000 60062 389056
rect 57145 388998 60062 389000
rect 217685 389058 217751 389061
rect 219390 389058 220064 389092
rect 217685 389056 220064 389058
rect 217685 389000 217690 389056
rect 217746 389032 220064 389056
rect 376937 389058 377003 389061
rect 379470 389058 380052 389092
rect 376937 389056 380052 389058
rect 217746 389000 219450 389032
rect 217685 388998 219450 389000
rect 376937 389000 376942 389056
rect 376998 389032 380052 389056
rect 376998 389000 379530 389032
rect 376937 388998 379530 389000
rect 57145 388995 57211 388998
rect 217685 388995 217751 388998
rect 376937 388995 377003 388998
rect 53046 388452 53052 388516
rect 53116 388514 53122 388516
rect 53741 388514 53807 388517
rect 53116 388512 53807 388514
rect 53116 388456 53746 388512
rect 53802 388456 53807 388512
rect 53116 388454 53807 388456
rect 53116 388452 53122 388454
rect 53741 388451 53807 388454
rect 57462 388452 57468 388516
rect 57532 388514 57538 388516
rect 59537 388514 59603 388517
rect 57532 388512 59603 388514
rect 57532 388456 59542 388512
rect 59598 388456 59603 388512
rect 57532 388454 59603 388456
rect 57532 388452 57538 388454
rect 59537 388451 59603 388454
rect -960 384284 480 384524
rect 377438 382332 377444 382396
rect 377508 382394 377514 382396
rect 379697 382394 379763 382397
rect 377508 382392 379763 382394
rect 377508 382336 379702 382392
rect 379758 382336 379763 382392
rect 377508 382334 379763 382336
rect 377508 382332 377514 382334
rect 379697 382331 379763 382334
rect 199142 381516 199148 381580
rect 199212 381578 199218 381580
rect 209405 381578 209471 381581
rect 199212 381576 209471 381578
rect 199212 381520 209410 381576
rect 209466 381520 209471 381576
rect 199212 381518 209471 381520
rect 199212 381516 199218 381518
rect 209405 381515 209471 381518
rect 49601 380898 49667 380901
rect 216673 380898 216739 380901
rect 49601 380896 216739 380898
rect 49601 380840 49606 380896
rect 49662 380840 216678 380896
rect 216734 380840 216739 380896
rect 49601 380838 216739 380840
rect 49601 380835 49667 380838
rect 216673 380835 216739 380838
rect 216949 380898 217015 380901
rect 217317 380898 217383 380901
rect 216949 380896 217383 380898
rect 216949 380840 216954 380896
rect 217010 380840 217322 380896
rect 217378 380840 217383 380896
rect 216949 380838 217383 380840
rect 216949 380835 217015 380838
rect 217317 380835 217383 380838
rect 248229 380900 248295 380901
rect 431125 380900 431191 380901
rect 433609 380900 433675 380901
rect 438485 380900 438551 380901
rect 248229 380896 248294 380900
rect 248229 380840 248234 380896
rect 248290 380840 248294 380896
rect 248229 380836 248294 380840
rect 248358 380898 248364 380900
rect 248358 380838 248386 380898
rect 248358 380836 248364 380838
rect 359774 380836 359780 380900
rect 359844 380898 359850 380900
rect 428280 380898 428286 380900
rect 359844 380838 428286 380898
rect 359844 380836 359850 380838
rect 428280 380836 428286 380838
rect 428350 380836 428356 380900
rect 431125 380896 431142 380900
rect 431206 380898 431212 380900
rect 433584 380898 433590 380900
rect 431125 380840 431130 380896
rect 431125 380836 431142 380840
rect 431206 380838 431282 380898
rect 433518 380838 433590 380898
rect 433654 380896 433675 380900
rect 438480 380898 438486 380900
rect 433670 380840 433675 380896
rect 431206 380836 431212 380838
rect 433584 380836 433590 380838
rect 433654 380836 433675 380840
rect 438394 380838 438486 380898
rect 438480 380836 438486 380838
rect 438550 380836 438556 380900
rect 248229 380835 248295 380836
rect 431125 380835 431191 380836
rect 433609 380835 433675 380836
rect 438485 380835 438551 380836
rect 110965 380764 111031 380765
rect 113541 380764 113607 380765
rect 116025 380764 116091 380765
rect 118417 380764 118483 380765
rect 120993 380764 121059 380765
rect 110965 380760 111006 380764
rect 111070 380762 111076 380764
rect 110965 380704 110970 380760
rect 110965 380700 111006 380704
rect 111070 380702 111122 380762
rect 113541 380760 113590 380764
rect 113654 380762 113660 380764
rect 113541 380704 113546 380760
rect 111070 380700 111076 380702
rect 113541 380700 113590 380704
rect 113654 380702 113698 380762
rect 116025 380760 116038 380764
rect 116102 380762 116108 380764
rect 116025 380704 116030 380760
rect 113654 380700 113660 380702
rect 116025 380700 116038 380704
rect 116102 380702 116182 380762
rect 118417 380760 118486 380764
rect 118417 380704 118422 380760
rect 118478 380704 118486 380760
rect 116102 380700 116108 380702
rect 118417 380700 118486 380704
rect 118550 380762 118556 380764
rect 120928 380762 120934 380764
rect 118550 380702 118574 380762
rect 120902 380702 120934 380762
rect 118550 380700 118556 380702
rect 120928 380700 120934 380702
rect 120998 380760 121059 380764
rect 121054 380704 121059 380760
rect 120998 380700 121059 380704
rect 110965 380699 111031 380700
rect 113541 380699 113607 380700
rect 116025 380699 116091 380700
rect 118417 380699 118483 380700
rect 120993 380699 121059 380700
rect 123477 380764 123543 380765
rect 125961 380764 126027 380765
rect 131021 380764 131087 380765
rect 133505 380764 133571 380765
rect 140957 380764 141023 380765
rect 143533 380764 143599 380765
rect 146017 380764 146083 380765
rect 155953 380764 156019 380765
rect 158529 380764 158595 380765
rect 160921 380764 160987 380765
rect 163405 380764 163471 380765
rect 165981 380764 166047 380765
rect 123477 380760 123518 380764
rect 123582 380762 123588 380764
rect 123477 380704 123482 380760
rect 123477 380700 123518 380704
rect 123582 380702 123634 380762
rect 123582 380700 123588 380702
rect 125960 380700 125966 380764
rect 126030 380762 126036 380764
rect 130992 380762 130998 380764
rect 126030 380702 126118 380762
rect 130930 380702 130998 380762
rect 131062 380760 131087 380764
rect 133440 380762 133446 380764
rect 131082 380704 131087 380760
rect 126030 380700 126036 380702
rect 130992 380700 130998 380702
rect 131062 380700 131087 380704
rect 133414 380702 133446 380762
rect 133440 380700 133446 380702
rect 133510 380760 133571 380764
rect 140920 380762 140926 380764
rect 133566 380704 133571 380760
rect 133510 380700 133571 380704
rect 140866 380702 140926 380762
rect 140990 380760 141023 380764
rect 143504 380762 143510 380764
rect 141018 380704 141023 380760
rect 140920 380700 140926 380702
rect 140990 380700 141023 380704
rect 143442 380702 143510 380762
rect 143574 380760 143599 380764
rect 145952 380762 145958 380764
rect 143594 380704 143599 380760
rect 143504 380700 143510 380702
rect 143574 380700 143599 380704
rect 145926 380702 145958 380762
rect 145952 380700 145958 380702
rect 146022 380760 146083 380764
rect 155880 380762 155886 380764
rect 146078 380704 146083 380760
rect 146022 380700 146083 380704
rect 155862 380702 155886 380762
rect 155880 380700 155886 380702
rect 155950 380760 156019 380764
rect 158464 380762 158470 380764
rect 155950 380704 155958 380760
rect 156014 380704 156019 380760
rect 155950 380700 156019 380704
rect 158438 380702 158470 380762
rect 158464 380700 158470 380702
rect 158534 380760 158595 380764
rect 160912 380762 160918 380764
rect 158590 380704 158595 380760
rect 158534 380700 158595 380704
rect 160830 380702 160918 380762
rect 160912 380700 160918 380702
rect 160982 380700 160988 380764
rect 163360 380762 163366 380764
rect 163314 380702 163366 380762
rect 163430 380760 163471 380764
rect 165944 380762 165950 380764
rect 163466 380704 163471 380760
rect 163360 380700 163366 380702
rect 163430 380700 163471 380704
rect 165890 380702 165950 380762
rect 166014 380760 166047 380764
rect 166042 380704 166047 380760
rect 165944 380700 165950 380702
rect 166014 380700 166047 380704
rect 202638 380700 202644 380764
rect 202708 380762 202714 380764
rect 202781 380762 202847 380765
rect 205173 380764 205239 380765
rect 205173 380762 205220 380764
rect 202708 380760 202847 380762
rect 202708 380704 202786 380760
rect 202842 380704 202847 380760
rect 202708 380702 202847 380704
rect 205128 380760 205220 380762
rect 205128 380704 205178 380760
rect 205128 380702 205220 380704
rect 202708 380700 202714 380702
rect 123477 380699 123543 380700
rect 125961 380699 126027 380700
rect 131021 380699 131087 380700
rect 133505 380699 133571 380700
rect 140957 380699 141023 380700
rect 143533 380699 143599 380700
rect 146017 380699 146083 380700
rect 155953 380699 156019 380700
rect 158529 380699 158595 380700
rect 160921 380699 160987 380700
rect 163405 380699 163471 380700
rect 165981 380699 166047 380700
rect 202781 380699 202847 380702
rect 205173 380700 205220 380702
rect 205284 380700 205290 380764
rect 208393 380762 208459 380765
rect 209681 380762 209747 380765
rect 410701 380764 410767 380765
rect 421097 380764 421163 380765
rect 279160 380762 279166 380764
rect 208393 380760 279166 380762
rect 208393 380704 208398 380760
rect 208454 380704 209686 380760
rect 209742 380704 279166 380760
rect 208393 380702 279166 380704
rect 205173 380699 205239 380700
rect 208393 380699 208459 380702
rect 209681 380699 209747 380702
rect 279160 380700 279166 380702
rect 279230 380700 279236 380764
rect 410701 380760 410742 380764
rect 410806 380762 410812 380764
rect 421072 380762 421078 380764
rect 410701 380704 410706 380760
rect 410701 380700 410742 380704
rect 410806 380702 410858 380762
rect 421006 380702 421078 380762
rect 421142 380760 421163 380764
rect 421158 380704 421163 380760
rect 410806 380700 410812 380702
rect 421072 380700 421078 380702
rect 421142 380700 421163 380704
rect 410701 380699 410767 380700
rect 421097 380699 421163 380700
rect 436001 380764 436067 380765
rect 440877 380764 440943 380765
rect 443453 380764 443519 380765
rect 436001 380760 436038 380764
rect 436102 380762 436108 380764
rect 436001 380704 436006 380760
rect 436001 380700 436038 380704
rect 436102 380702 436158 380762
rect 440877 380760 440934 380764
rect 440998 380762 441004 380764
rect 440877 380704 440882 380760
rect 436102 380700 436108 380702
rect 440877 380700 440934 380704
rect 440998 380702 441034 380762
rect 443453 380760 443518 380764
rect 443453 380704 443458 380760
rect 443514 380704 443518 380760
rect 440998 380700 441004 380702
rect 443453 380700 443518 380704
rect 443582 380762 443588 380764
rect 443582 380702 443610 380762
rect 443582 380700 443588 380702
rect 436001 380699 436067 380700
rect 440877 380699 440943 380700
rect 443453 380699 443519 380700
rect 52361 380626 52427 380629
rect 216949 380626 217015 380629
rect 52361 380624 217015 380626
rect 52361 380568 52366 380624
rect 52422 380568 216954 380624
rect 217010 380568 217015 380624
rect 52361 380566 217015 380568
rect 52361 380563 52427 380566
rect 216949 380563 217015 380566
rect 217133 380626 217199 380629
rect 217593 380626 217659 380629
rect 217133 380624 217659 380626
rect 217133 380568 217138 380624
rect 217194 380568 217598 380624
rect 217654 380568 217659 380624
rect 217133 380566 217659 380568
rect 217133 380563 217199 380566
rect 217593 380563 217659 380566
rect 235993 380628 236059 380629
rect 237097 380628 237163 380629
rect 243077 380628 243143 380629
rect 245377 380628 245443 380629
rect 247585 380628 247651 380629
rect 254485 380628 254551 380629
rect 255865 380628 255931 380629
rect 256969 380628 257035 380629
rect 258073 380628 258139 380629
rect 259453 380628 259519 380629
rect 265249 380628 265315 380629
rect 235993 380624 236054 380628
rect 235993 380568 235998 380624
rect 235993 380564 236054 380568
rect 236118 380626 236124 380628
rect 236118 380566 236150 380626
rect 237097 380624 237142 380628
rect 237206 380626 237212 380628
rect 237097 380568 237102 380624
rect 236118 380564 236124 380566
rect 237097 380564 237142 380568
rect 237206 380566 237254 380626
rect 243077 380624 243126 380628
rect 243190 380626 243196 380628
rect 243077 380568 243082 380624
rect 237206 380564 237212 380566
rect 243077 380564 243126 380568
rect 243190 380566 243234 380626
rect 245377 380624 245438 380628
rect 245377 380568 245382 380624
rect 243190 380564 243196 380566
rect 245377 380564 245438 380568
rect 245502 380626 245508 380628
rect 245502 380566 245534 380626
rect 247585 380624 247614 380628
rect 247678 380626 247684 380628
rect 247585 380568 247590 380624
rect 245502 380564 245508 380566
rect 247585 380564 247614 380568
rect 247678 380566 247742 380626
rect 254485 380624 254550 380628
rect 254485 380568 254490 380624
rect 254546 380568 254550 380624
rect 247678 380564 247684 380566
rect 254485 380564 254550 380568
rect 254614 380626 254620 380628
rect 254614 380566 254642 380626
rect 255865 380624 255910 380628
rect 255974 380626 255980 380628
rect 255865 380568 255870 380624
rect 254614 380564 254620 380566
rect 255865 380564 255910 380568
rect 255974 380566 256022 380626
rect 256969 380624 256998 380628
rect 257062 380626 257068 380628
rect 256969 380568 256974 380624
rect 255974 380564 255980 380566
rect 256969 380564 256998 380568
rect 257062 380566 257126 380626
rect 258073 380624 258086 380628
rect 258150 380626 258156 380628
rect 259440 380626 259446 380628
rect 258073 380568 258078 380624
rect 257062 380564 257068 380566
rect 258073 380564 258086 380568
rect 258150 380566 258230 380626
rect 259362 380566 259446 380626
rect 259510 380624 259519 380628
rect 259514 380568 259519 380624
rect 258150 380564 258156 380566
rect 259440 380564 259446 380566
rect 259510 380564 259519 380568
rect 260664 380564 260670 380628
rect 260734 380564 260740 380628
rect 265249 380624 265294 380628
rect 265358 380626 265364 380628
rect 265525 380626 265591 380629
rect 270953 380628 271019 380629
rect 405457 380628 405523 380629
rect 413461 380628 413527 380629
rect 419441 380628 419507 380629
rect 434345 380628 434411 380629
rect 485957 380628 486023 380629
rect 269776 380626 269782 380628
rect 265249 380568 265254 380624
rect 265249 380564 265294 380568
rect 265358 380566 265406 380626
rect 265525 380624 269782 380626
rect 265525 380568 265530 380624
rect 265586 380568 269782 380624
rect 265525 380566 269782 380568
rect 265358 380564 265364 380566
rect 235993 380563 236059 380564
rect 237097 380563 237163 380564
rect 243077 380563 243143 380564
rect 245377 380563 245443 380564
rect 247585 380563 247651 380564
rect 254485 380563 254551 380564
rect 255865 380563 255931 380564
rect 256969 380563 257035 380564
rect 258073 380563 258139 380564
rect 259453 380563 259519 380564
rect 76046 380428 76052 380492
rect 76116 380490 76122 380492
rect 202965 380490 203031 380493
rect 213821 380490 213887 380493
rect 76116 380488 213887 380490
rect 76116 380432 202970 380488
rect 203026 380432 213826 380488
rect 213882 380432 213887 380488
rect 76116 380430 213887 380432
rect 76116 380428 76122 380430
rect 202965 380427 203031 380430
rect 213821 380427 213887 380430
rect 216673 380490 216739 380493
rect 217777 380490 217843 380493
rect 216673 380488 217843 380490
rect 216673 380432 216678 380488
rect 216734 380432 217782 380488
rect 217838 380432 217843 380488
rect 216673 380430 217843 380432
rect 216673 380427 216739 380430
rect 217777 380427 217843 380430
rect 217910 380428 217916 380492
rect 217980 380490 217986 380492
rect 260672 380490 260732 380564
rect 265249 380563 265315 380564
rect 265525 380563 265591 380566
rect 269776 380564 269782 380566
rect 269846 380564 269852 380628
rect 270953 380624 271006 380628
rect 271070 380626 271076 380628
rect 405432 380626 405438 380628
rect 270953 380568 270958 380624
rect 270953 380564 271006 380568
rect 271070 380566 271110 380626
rect 405366 380566 405438 380626
rect 405502 380624 405523 380628
rect 413456 380626 413462 380628
rect 405518 380568 405523 380624
rect 271070 380564 271076 380566
rect 405432 380564 405438 380566
rect 405502 380564 405523 380568
rect 413370 380566 413462 380626
rect 413456 380564 413462 380566
rect 413526 380564 413532 380628
rect 419440 380564 419446 380628
rect 419510 380626 419516 380628
rect 419510 380566 419598 380626
rect 434345 380624 434406 380628
rect 434345 380568 434350 380624
rect 419510 380564 419516 380566
rect 434345 380564 434406 380568
rect 434470 380626 434476 380628
rect 485944 380626 485950 380628
rect 434470 380566 434502 380626
rect 485866 380566 485950 380626
rect 486014 380624 486023 380628
rect 486018 380568 486023 380624
rect 434470 380564 434476 380566
rect 485944 380564 485950 380566
rect 486014 380564 486023 380568
rect 270953 380563 271019 380564
rect 405457 380563 405523 380564
rect 413461 380563 413527 380564
rect 419441 380563 419507 380564
rect 434345 380563 434411 380564
rect 485957 380563 486023 380564
rect 426433 380492 426499 380493
rect 426382 380490 426388 380492
rect 217980 380430 260732 380490
rect 426342 380430 426388 380490
rect 426452 380488 426499 380492
rect 426494 380432 426499 380488
rect 217980 380428 217986 380430
rect 426382 380428 426388 380430
rect 426452 380428 426499 380432
rect 426433 380427 426499 380428
rect 119102 380292 119108 380356
rect 119172 380354 119178 380356
rect 208393 380354 208459 380357
rect 119172 380352 208459 380354
rect 119172 380296 208398 380352
rect 208454 380296 208459 380352
rect 119172 380294 208459 380296
rect 119172 380292 119178 380294
rect 208393 380291 208459 380294
rect 216990 380292 216996 380356
rect 217060 380354 217066 380356
rect 323342 380354 323348 380356
rect 217060 380294 323348 380354
rect 217060 380292 217066 380294
rect 323342 380292 323348 380294
rect 323412 380292 323418 380356
rect 128353 380220 128419 380221
rect 128302 380218 128308 380220
rect 128262 380158 128308 380218
rect 128372 380216 128419 380220
rect 128414 380160 128419 380216
rect 128302 380156 128308 380158
rect 128372 380156 128419 380160
rect 216622 380156 216628 380220
rect 216692 380218 216698 380220
rect 217542 380218 217548 380220
rect 216692 380158 217548 380218
rect 216692 380156 216698 380158
rect 217542 380156 217548 380158
rect 217612 380156 217618 380220
rect 279182 380156 279188 380220
rect 279252 380218 279258 380220
rect 357433 380218 357499 380221
rect 279252 380216 357499 380218
rect 279252 380160 357438 380216
rect 357494 380160 357499 380216
rect 279252 380158 357499 380160
rect 279252 380156 279258 380158
rect 128353 380155 128419 380156
rect 357433 380155 357499 380158
rect 359590 380156 359596 380220
rect 359660 380218 359666 380220
rect 371785 380218 371851 380221
rect 404118 380218 404124 380220
rect 359660 380216 404124 380218
rect 359660 380160 371790 380216
rect 371846 380160 404124 380216
rect 359660 380158 404124 380160
rect 359660 380156 359666 380158
rect 371785 380155 371851 380158
rect 404118 380156 404124 380158
rect 404188 380156 404194 380220
rect 51533 380082 51599 380085
rect 217593 380082 217659 380085
rect 51533 380080 217659 380082
rect 51533 380024 51538 380080
rect 51594 380024 217598 380080
rect 217654 380024 217659 380080
rect 51533 380022 217659 380024
rect 51533 380019 51599 380022
rect 217593 380019 217659 380022
rect 50286 379476 50292 379540
rect 50356 379538 50362 379540
rect 50981 379538 51047 379541
rect 50356 379536 51047 379538
rect 50356 379480 50986 379536
rect 51042 379480 51047 379536
rect 50356 379478 51047 379480
rect 50356 379476 50362 379478
rect 50981 379475 51047 379478
rect 51942 379476 51948 379540
rect 52012 379538 52018 379540
rect 52269 379538 52335 379541
rect 52012 379536 52335 379538
rect 52012 379480 52274 379536
rect 52330 379480 52335 379536
rect 52012 379478 52335 379480
rect 52012 379476 52018 379478
rect 52269 379475 52335 379478
rect 208342 379476 208348 379540
rect 208412 379538 208418 379540
rect 208853 379538 208919 379541
rect 208412 379536 208919 379538
rect 208412 379480 208858 379536
rect 208914 379480 208919 379536
rect 208412 379478 208919 379480
rect 208412 379476 208418 379478
rect 208853 379475 208919 379478
rect 47393 379402 47459 379405
rect 85481 379404 85547 379405
rect 86585 379404 86651 379405
rect 81750 379402 81756 379404
rect 47393 379400 81756 379402
rect 47393 379344 47398 379400
rect 47454 379344 81756 379400
rect 47393 379342 81756 379344
rect 47393 379339 47459 379342
rect 81750 379340 81756 379342
rect 81820 379402 81826 379404
rect 81934 379402 81940 379404
rect 81820 379342 81940 379402
rect 81820 379340 81826 379342
rect 81934 379340 81940 379342
rect 82004 379340 82010 379404
rect 85430 379402 85436 379404
rect 85390 379342 85436 379402
rect 85500 379400 85547 379404
rect 86534 379402 86540 379404
rect 85542 379344 85547 379400
rect 85430 379340 85436 379342
rect 85500 379340 85547 379344
rect 86494 379342 86540 379402
rect 86604 379400 86651 379404
rect 86646 379344 86651 379400
rect 86534 379340 86540 379342
rect 86604 379340 86651 379344
rect 87638 379340 87644 379404
rect 87708 379402 87714 379404
rect 87873 379402 87939 379405
rect 87708 379400 87939 379402
rect 87708 379344 87878 379400
rect 87934 379344 87939 379400
rect 87708 379342 87939 379344
rect 87708 379340 87714 379342
rect 85481 379339 85547 379340
rect 86585 379339 86651 379340
rect 87873 379339 87939 379342
rect 88333 379404 88399 379405
rect 88793 379404 88859 379405
rect 90081 379404 90147 379405
rect 88333 379400 88380 379404
rect 88444 379402 88450 379404
rect 88742 379402 88748 379404
rect 88333 379344 88338 379400
rect 88333 379340 88380 379344
rect 88444 379342 88490 379402
rect 88702 379342 88748 379402
rect 88812 379400 88859 379404
rect 90030 379402 90036 379404
rect 88854 379344 88859 379400
rect 88444 379340 88450 379342
rect 88742 379340 88748 379342
rect 88812 379340 88859 379344
rect 89990 379342 90036 379402
rect 90100 379400 90147 379404
rect 90142 379344 90147 379400
rect 90030 379340 90036 379342
rect 90100 379340 90147 379344
rect 88333 379339 88399 379340
rect 88793 379339 88859 379340
rect 90081 379339 90147 379340
rect 90633 379402 90699 379405
rect 91369 379404 91435 379405
rect 90766 379402 90772 379404
rect 90633 379400 90772 379402
rect 90633 379344 90638 379400
rect 90694 379344 90772 379400
rect 90633 379342 90772 379344
rect 90633 379339 90699 379342
rect 90766 379340 90772 379342
rect 90836 379340 90842 379404
rect 91318 379402 91324 379404
rect 91278 379342 91324 379402
rect 91388 379400 91435 379404
rect 91430 379344 91435 379400
rect 91318 379340 91324 379342
rect 91388 379340 91435 379344
rect 91369 379339 91435 379340
rect 92381 379404 92447 379405
rect 92381 379400 92428 379404
rect 92492 379402 92498 379404
rect 92381 379344 92386 379400
rect 92381 379340 92428 379344
rect 92492 379342 92538 379402
rect 92492 379340 92498 379342
rect 93342 379340 93348 379404
rect 93412 379402 93418 379404
rect 93577 379402 93643 379405
rect 93412 379400 93643 379402
rect 93412 379344 93582 379400
rect 93638 379344 93643 379400
rect 93412 379342 93643 379344
rect 93412 379340 93418 379342
rect 92381 379339 92447 379340
rect 93577 379339 93643 379342
rect 96061 379404 96127 379405
rect 96061 379400 96108 379404
rect 96172 379402 96178 379404
rect 96061 379344 96066 379400
rect 96061 379340 96108 379344
rect 96172 379342 96218 379402
rect 96172 379340 96178 379342
rect 98126 379340 98132 379404
rect 98196 379402 98202 379404
rect 98269 379402 98335 379405
rect 98196 379400 98335 379402
rect 98196 379344 98274 379400
rect 98330 379344 98335 379400
rect 98196 379342 98335 379344
rect 98196 379340 98202 379342
rect 96061 379339 96127 379340
rect 98269 379339 98335 379342
rect 98453 379404 98519 379405
rect 101029 379404 101095 379405
rect 98453 379400 98500 379404
rect 98564 379402 98570 379404
rect 98453 379344 98458 379400
rect 98453 379340 98500 379344
rect 98564 379342 98610 379402
rect 101029 379400 101076 379404
rect 101140 379402 101146 379404
rect 101029 379344 101034 379400
rect 98564 379340 98570 379342
rect 101029 379340 101076 379344
rect 101140 379342 101186 379402
rect 101140 379340 101146 379342
rect 103278 379340 103284 379404
rect 103348 379402 103354 379404
rect 103513 379402 103579 379405
rect 103348 379400 103579 379402
rect 103348 379344 103518 379400
rect 103574 379344 103579 379400
rect 103348 379342 103579 379344
rect 103348 379340 103354 379342
rect 98453 379339 98519 379340
rect 101029 379339 101095 379340
rect 103513 379339 103579 379342
rect 104893 379402 104959 379405
rect 108205 379404 108271 379405
rect 108849 379404 108915 379405
rect 105854 379402 105860 379404
rect 104893 379400 105860 379402
rect 104893 379344 104898 379400
rect 104954 379344 105860 379400
rect 104893 379342 105860 379344
rect 104893 379339 104959 379342
rect 105854 379340 105860 379342
rect 105924 379340 105930 379404
rect 108205 379400 108252 379404
rect 108316 379402 108322 379404
rect 108798 379402 108804 379404
rect 108205 379344 108210 379400
rect 108205 379340 108252 379344
rect 108316 379342 108362 379402
rect 108758 379342 108804 379402
rect 108868 379400 108915 379404
rect 108910 379344 108915 379400
rect 108316 379340 108322 379342
rect 108798 379340 108804 379342
rect 108868 379340 108915 379344
rect 111190 379340 111196 379404
rect 111260 379402 111266 379404
rect 111333 379402 111399 379405
rect 112345 379404 112411 379405
rect 113449 379404 113515 379405
rect 112294 379402 112300 379404
rect 111260 379400 111399 379402
rect 111260 379344 111338 379400
rect 111394 379344 111399 379400
rect 111260 379342 111399 379344
rect 112254 379342 112300 379402
rect 112364 379400 112411 379404
rect 113398 379402 113404 379404
rect 112406 379344 112411 379400
rect 111260 379340 111266 379342
rect 108205 379339 108271 379340
rect 108849 379339 108915 379340
rect 111333 379339 111399 379342
rect 112294 379340 112300 379342
rect 112364 379340 112411 379344
rect 113358 379342 113404 379402
rect 113468 379400 113515 379404
rect 113510 379344 113515 379400
rect 113398 379340 113404 379342
rect 113468 379340 113515 379344
rect 112345 379339 112411 379340
rect 113449 379339 113515 379340
rect 114461 379404 114527 379405
rect 115841 379404 115907 379405
rect 135897 379404 135963 379405
rect 138473 379404 138539 379405
rect 150985 379404 151051 379405
rect 114461 379400 114508 379404
rect 114572 379402 114578 379404
rect 115790 379402 115796 379404
rect 114461 379344 114466 379400
rect 114461 379340 114508 379344
rect 114572 379342 114618 379402
rect 115750 379342 115796 379402
rect 115860 379400 115907 379404
rect 135846 379402 135852 379404
rect 115902 379344 115907 379400
rect 114572 379340 114578 379342
rect 115790 379340 115796 379342
rect 115860 379340 115907 379344
rect 135806 379342 135852 379402
rect 135916 379400 135963 379404
rect 138422 379402 138428 379404
rect 135958 379344 135963 379400
rect 135846 379340 135852 379342
rect 135916 379340 135963 379344
rect 138382 379342 138428 379402
rect 138492 379400 138539 379404
rect 150934 379402 150940 379404
rect 138534 379344 138539 379400
rect 138422 379340 138428 379342
rect 138492 379340 138539 379344
rect 150894 379342 150940 379402
rect 151004 379400 151051 379404
rect 151046 379344 151051 379400
rect 150934 379340 150940 379342
rect 151004 379340 151051 379344
rect 153510 379340 153516 379404
rect 153580 379402 153586 379404
rect 154021 379402 154087 379405
rect 207013 379402 207079 379405
rect 153580 379400 154087 379402
rect 153580 379344 154026 379400
rect 154082 379344 154087 379400
rect 153580 379342 154087 379344
rect 153580 379340 153586 379342
rect 114461 379339 114527 379340
rect 115841 379339 115907 379340
rect 135897 379339 135963 379340
rect 138473 379339 138539 379340
rect 150985 379339 151051 379340
rect 154021 379339 154087 379342
rect 195930 379400 207079 379402
rect 195930 379344 207018 379400
rect 207074 379344 207079 379400
rect 195930 379342 207079 379344
rect 46105 379266 46171 379269
rect 80421 379268 80487 379269
rect 46105 379264 64890 379266
rect 46105 379208 46110 379264
rect 46166 379208 64890 379264
rect 46105 379206 64890 379208
rect 46105 379203 46171 379206
rect 51533 379130 51599 379133
rect 57094 379130 57100 379132
rect 51533 379128 57100 379130
rect 51533 379072 51538 379128
rect 51594 379072 57100 379128
rect 51533 379070 57100 379072
rect 51533 379067 51599 379070
rect 57094 379068 57100 379070
rect 57164 379068 57170 379132
rect 64830 379130 64890 379206
rect 80421 379264 80468 379268
rect 80532 379266 80538 379268
rect 93485 379266 93551 379269
rect 95969 379268 96035 379269
rect 99465 379268 99531 379269
rect 102961 379268 103027 379269
rect 93710 379266 93716 379268
rect 80421 379208 80426 379264
rect 80421 379204 80468 379208
rect 80532 379206 80578 379266
rect 93485 379264 93716 379266
rect 93485 379208 93490 379264
rect 93546 379208 93716 379264
rect 93485 379206 93716 379208
rect 80532 379204 80538 379206
rect 80421 379203 80487 379204
rect 93485 379203 93551 379206
rect 93710 379204 93716 379206
rect 93780 379204 93786 379268
rect 95918 379266 95924 379268
rect 95878 379206 95924 379266
rect 95988 379264 96035 379268
rect 99414 379266 99420 379268
rect 96030 379208 96035 379264
rect 95918 379204 95924 379206
rect 95988 379204 96035 379208
rect 99374 379206 99420 379266
rect 99484 379264 99531 379268
rect 102910 379266 102916 379268
rect 99526 379208 99531 379264
rect 99414 379204 99420 379206
rect 99484 379204 99531 379208
rect 102870 379206 102916 379266
rect 102980 379264 103027 379268
rect 103022 379208 103027 379264
rect 102910 379204 102916 379206
rect 102980 379204 103027 379208
rect 109718 379204 109724 379268
rect 109788 379266 109794 379268
rect 195930 379266 195990 379342
rect 207013 379339 207079 379342
rect 246205 379402 246271 379405
rect 248597 379404 248663 379405
rect 250069 379404 250135 379405
rect 251173 379404 251239 379405
rect 252277 379404 252343 379405
rect 253381 379404 253447 379405
rect 261661 379404 261727 379405
rect 263869 379404 263935 379405
rect 268653 379404 268719 379405
rect 271045 379404 271111 379405
rect 272149 379404 272215 379405
rect 273253 379404 273319 379405
rect 274357 379404 274423 379405
rect 275645 379404 275711 379405
rect 276105 379404 276171 379405
rect 277025 379404 277091 379405
rect 246430 379402 246436 379404
rect 246205 379400 246436 379402
rect 246205 379344 246210 379400
rect 246266 379344 246436 379400
rect 246205 379342 246436 379344
rect 246205 379339 246271 379342
rect 246430 379340 246436 379342
rect 246500 379340 246506 379404
rect 248597 379400 248644 379404
rect 248708 379402 248714 379404
rect 248597 379344 248602 379400
rect 248597 379340 248644 379344
rect 248708 379342 248754 379402
rect 250069 379400 250116 379404
rect 250180 379402 250186 379404
rect 250069 379344 250074 379400
rect 248708 379340 248714 379342
rect 250069 379340 250116 379344
rect 250180 379342 250226 379402
rect 251173 379400 251220 379404
rect 251284 379402 251290 379404
rect 251173 379344 251178 379400
rect 250180 379340 250186 379342
rect 251173 379340 251220 379344
rect 251284 379342 251330 379402
rect 252277 379400 252324 379404
rect 252388 379402 252394 379404
rect 252277 379344 252282 379400
rect 251284 379340 251290 379342
rect 252277 379340 252324 379344
rect 252388 379342 252434 379402
rect 253381 379400 253428 379404
rect 253492 379402 253498 379404
rect 253381 379344 253386 379400
rect 252388 379340 252394 379342
rect 253381 379340 253428 379344
rect 253492 379342 253538 379402
rect 261661 379400 261708 379404
rect 261772 379402 261778 379404
rect 261661 379344 261666 379400
rect 253492 379340 253498 379342
rect 261661 379340 261708 379344
rect 261772 379342 261818 379402
rect 263869 379400 263916 379404
rect 263980 379402 263986 379404
rect 263869 379344 263874 379400
rect 261772 379340 261778 379342
rect 263869 379340 263916 379344
rect 263980 379342 264026 379402
rect 268653 379400 268700 379404
rect 268764 379402 268770 379404
rect 268653 379344 268658 379400
rect 263980 379340 263986 379342
rect 268653 379340 268700 379344
rect 268764 379342 268810 379402
rect 271045 379400 271092 379404
rect 271156 379402 271162 379404
rect 271045 379344 271050 379400
rect 268764 379340 268770 379342
rect 271045 379340 271092 379344
rect 271156 379342 271202 379402
rect 272149 379400 272196 379404
rect 272260 379402 272266 379404
rect 272149 379344 272154 379400
rect 271156 379340 271162 379342
rect 272149 379340 272196 379344
rect 272260 379342 272306 379402
rect 273253 379400 273300 379404
rect 273364 379402 273370 379404
rect 273253 379344 273258 379400
rect 272260 379340 272266 379342
rect 273253 379340 273300 379344
rect 273364 379342 273410 379402
rect 274357 379400 274404 379404
rect 274468 379402 274474 379404
rect 274357 379344 274362 379400
rect 273364 379340 273370 379342
rect 274357 379340 274404 379344
rect 274468 379342 274514 379402
rect 275645 379400 275692 379404
rect 275756 379402 275762 379404
rect 276054 379402 276060 379404
rect 275645 379344 275650 379400
rect 274468 379340 274474 379342
rect 275645 379340 275692 379344
rect 275756 379342 275802 379402
rect 276014 379342 276060 379402
rect 276124 379400 276171 379404
rect 276974 379402 276980 379404
rect 276166 379344 276171 379400
rect 275756 379340 275762 379342
rect 276054 379340 276060 379342
rect 276124 379340 276171 379344
rect 276934 379342 276980 379402
rect 277044 379400 277091 379404
rect 277086 379344 277091 379400
rect 276974 379340 276980 379342
rect 277044 379340 277091 379344
rect 248597 379339 248663 379340
rect 250069 379339 250135 379340
rect 251173 379339 251239 379340
rect 252277 379339 252343 379340
rect 253381 379339 253447 379340
rect 261661 379339 261727 379340
rect 263869 379339 263935 379340
rect 268653 379339 268719 379340
rect 271045 379339 271111 379340
rect 272149 379339 272215 379340
rect 273253 379339 273319 379340
rect 274357 379339 274423 379340
rect 275645 379339 275711 379340
rect 276105 379339 276171 379340
rect 277025 379339 277091 379340
rect 278221 379402 278287 379405
rect 285949 379404 286015 379405
rect 278446 379402 278452 379404
rect 278221 379400 278452 379402
rect 278221 379344 278226 379400
rect 278282 379344 278452 379400
rect 278221 379342 278452 379344
rect 278221 379339 278287 379342
rect 278446 379340 278452 379342
rect 278516 379340 278522 379404
rect 285949 379400 285996 379404
rect 286060 379402 286066 379404
rect 287605 379402 287671 379405
rect 290917 379404 290983 379405
rect 288198 379402 288204 379404
rect 285949 379344 285954 379400
rect 285949 379340 285996 379344
rect 286060 379342 286106 379402
rect 287605 379400 288204 379402
rect 287605 379344 287610 379400
rect 287666 379344 288204 379400
rect 287605 379342 288204 379344
rect 286060 379340 286066 379342
rect 285949 379339 286015 379340
rect 287605 379339 287671 379342
rect 288198 379340 288204 379342
rect 288268 379340 288274 379404
rect 290917 379400 290964 379404
rect 291028 379402 291034 379404
rect 292665 379402 292731 379405
rect 293350 379402 293356 379404
rect 290917 379344 290922 379400
rect 290917 379340 290964 379344
rect 291028 379342 291074 379402
rect 292665 379400 293356 379402
rect 292665 379344 292670 379400
rect 292726 379344 293356 379400
rect 292665 379342 293356 379344
rect 291028 379340 291034 379342
rect 290917 379339 290983 379340
rect 292665 379339 292731 379342
rect 293350 379340 293356 379342
rect 293420 379340 293426 379404
rect 295425 379402 295491 379405
rect 298461 379404 298527 379405
rect 300853 379404 300919 379405
rect 295926 379402 295932 379404
rect 295425 379400 295932 379402
rect 295425 379344 295430 379400
rect 295486 379344 295932 379400
rect 295425 379342 295932 379344
rect 295425 379339 295491 379342
rect 295926 379340 295932 379342
rect 295996 379340 296002 379404
rect 298461 379400 298508 379404
rect 298572 379402 298578 379404
rect 298461 379344 298466 379400
rect 298461 379340 298508 379344
rect 298572 379342 298618 379402
rect 300853 379400 300900 379404
rect 300964 379402 300970 379404
rect 303245 379402 303311 379405
rect 305821 379404 305887 379405
rect 303470 379402 303476 379404
rect 300853 379344 300858 379400
rect 298572 379340 298578 379342
rect 300853 379340 300900 379344
rect 300964 379342 301010 379402
rect 303245 379400 303476 379402
rect 303245 379344 303250 379400
rect 303306 379344 303476 379400
rect 303245 379342 303476 379344
rect 300964 379340 300970 379342
rect 298461 379339 298527 379340
rect 300853 379339 300919 379340
rect 303245 379339 303311 379342
rect 303470 379340 303476 379342
rect 303540 379340 303546 379404
rect 305821 379400 305868 379404
rect 305932 379402 305938 379404
rect 307845 379402 307911 379405
rect 310973 379404 311039 379405
rect 313365 379404 313431 379405
rect 315757 379404 315823 379405
rect 308438 379402 308444 379404
rect 305821 379344 305826 379400
rect 305821 379340 305868 379344
rect 305932 379342 305978 379402
rect 307845 379400 308444 379402
rect 307845 379344 307850 379400
rect 307906 379344 308444 379400
rect 307845 379342 308444 379344
rect 305932 379340 305938 379342
rect 305821 379339 305887 379340
rect 307845 379339 307911 379342
rect 308438 379340 308444 379342
rect 308508 379340 308514 379404
rect 310973 379400 311020 379404
rect 311084 379402 311090 379404
rect 310973 379344 310978 379400
rect 310973 379340 311020 379344
rect 311084 379342 311130 379402
rect 313365 379400 313412 379404
rect 313476 379402 313482 379404
rect 313365 379344 313370 379400
rect 311084 379340 311090 379342
rect 313365 379340 313412 379344
rect 313476 379342 313522 379402
rect 315757 379400 315804 379404
rect 315868 379402 315874 379404
rect 317413 379402 317479 379405
rect 396073 379404 396139 379405
rect 318374 379402 318380 379404
rect 315757 379344 315762 379400
rect 313476 379340 313482 379342
rect 315757 379340 315804 379344
rect 315868 379342 315914 379402
rect 317413 379400 318380 379402
rect 317413 379344 317418 379400
rect 317474 379344 318380 379400
rect 317413 379342 318380 379344
rect 315868 379340 315874 379342
rect 310973 379339 311039 379340
rect 313365 379339 313431 379340
rect 315757 379339 315823 379340
rect 317413 379339 317479 379342
rect 318374 379340 318380 379342
rect 318444 379340 318450 379404
rect 396022 379402 396028 379404
rect 395982 379342 396028 379402
rect 396092 379400 396139 379404
rect 396134 379344 396139 379400
rect 396022 379340 396028 379342
rect 396092 379340 396139 379344
rect 396073 379339 396139 379340
rect 397085 379404 397151 379405
rect 397085 379400 397132 379404
rect 397196 379402 397202 379404
rect 401726 379402 401732 379404
rect 397085 379344 397090 379400
rect 397085 379340 397132 379344
rect 397196 379342 397242 379402
rect 398054 379342 401732 379402
rect 397196 379340 397202 379342
rect 397085 379339 397151 379340
rect 109788 379206 195990 379266
rect 202965 379266 203031 379269
rect 205265 379266 205331 379269
rect 216305 379266 216371 379269
rect 278078 379266 278084 379268
rect 202965 379264 278084 379266
rect 202965 379208 202970 379264
rect 203026 379208 205270 379264
rect 205326 379208 216310 379264
rect 216366 379208 278084 379264
rect 202965 379206 278084 379208
rect 109788 379204 109794 379206
rect 95969 379203 96035 379204
rect 99465 379203 99531 379204
rect 102961 379203 103027 379204
rect 202965 379203 203031 379206
rect 205265 379203 205331 379206
rect 216305 379203 216371 379206
rect 278078 379204 278084 379206
rect 278148 379204 278154 379268
rect 280245 379266 280311 379269
rect 283373 379268 283439 379269
rect 325877 379268 325943 379269
rect 280838 379266 280844 379268
rect 280245 379264 280844 379266
rect 280245 379208 280250 379264
rect 280306 379208 280844 379264
rect 280245 379206 280844 379208
rect 280245 379203 280311 379206
rect 280838 379204 280844 379206
rect 280908 379204 280914 379268
rect 283373 379264 283420 379268
rect 283484 379266 283490 379268
rect 283373 379208 283378 379264
rect 283373 379204 283420 379208
rect 283484 379206 283530 379266
rect 325877 379264 325924 379268
rect 325988 379266 325994 379268
rect 398054 379266 398114 379342
rect 401726 379340 401732 379342
rect 401796 379340 401802 379404
rect 405825 379402 405891 379405
rect 407573 379404 407639 379405
rect 408309 379404 408375 379405
rect 411253 379404 411319 379405
rect 412357 379404 412423 379405
rect 406510 379402 406516 379404
rect 405825 379400 406516 379402
rect 405825 379344 405830 379400
rect 405886 379344 406516 379400
rect 405825 379342 406516 379344
rect 405825 379339 405891 379342
rect 406510 379340 406516 379342
rect 406580 379340 406586 379404
rect 407573 379400 407620 379404
rect 407684 379402 407690 379404
rect 407573 379344 407578 379400
rect 407573 379340 407620 379344
rect 407684 379342 407730 379402
rect 408309 379400 408356 379404
rect 408420 379402 408426 379404
rect 408309 379344 408314 379400
rect 407684 379340 407690 379342
rect 408309 379340 408356 379344
rect 408420 379342 408466 379402
rect 411253 379400 411300 379404
rect 411364 379402 411370 379404
rect 411253 379344 411258 379400
rect 408420 379340 408426 379342
rect 411253 379340 411300 379344
rect 411364 379342 411410 379402
rect 412357 379400 412404 379404
rect 412468 379402 412474 379404
rect 415669 379402 415735 379405
rect 425973 379404 426039 379405
rect 416078 379402 416084 379404
rect 412357 379344 412362 379400
rect 411364 379340 411370 379342
rect 412357 379340 412404 379344
rect 412468 379342 412514 379402
rect 415669 379400 416084 379402
rect 415669 379344 415674 379400
rect 415730 379344 416084 379400
rect 415669 379342 416084 379344
rect 412468 379340 412474 379342
rect 407573 379339 407639 379340
rect 408309 379339 408375 379340
rect 411253 379339 411319 379340
rect 412357 379339 412423 379340
rect 415669 379339 415735 379342
rect 416078 379340 416084 379342
rect 416148 379340 416154 379404
rect 425973 379400 426020 379404
rect 426084 379402 426090 379404
rect 435173 379402 435239 379405
rect 435766 379402 435772 379404
rect 425973 379344 425978 379400
rect 425973 379340 426020 379344
rect 426084 379342 426130 379402
rect 435173 379400 435772 379402
rect 435173 379344 435178 379400
rect 435234 379344 435772 379400
rect 435173 379342 435772 379344
rect 426084 379340 426090 379342
rect 425973 379339 426039 379340
rect 435173 379339 435239 379342
rect 435766 379340 435772 379342
rect 435836 379340 435842 379404
rect 437841 379402 437907 379405
rect 445845 379404 445911 379405
rect 437974 379402 437980 379404
rect 437841 379400 437980 379402
rect 437841 379344 437846 379400
rect 437902 379344 437980 379400
rect 437841 379342 437980 379344
rect 437841 379339 437907 379342
rect 437974 379340 437980 379342
rect 438044 379340 438050 379404
rect 445845 379400 445892 379404
rect 445956 379402 445962 379404
rect 447501 379402 447567 379405
rect 450997 379404 451063 379405
rect 448278 379402 448284 379404
rect 445845 379344 445850 379400
rect 445845 379340 445892 379344
rect 445956 379342 446002 379402
rect 447501 379400 448284 379402
rect 447501 379344 447506 379400
rect 447562 379344 448284 379400
rect 447501 379342 448284 379344
rect 445956 379340 445962 379342
rect 445845 379339 445911 379340
rect 447501 379339 447567 379342
rect 448278 379340 448284 379342
rect 448348 379340 448354 379404
rect 450997 379400 451044 379404
rect 451108 379402 451114 379404
rect 453021 379402 453087 379405
rect 453430 379402 453436 379404
rect 450997 379344 451002 379400
rect 450997 379340 451044 379344
rect 451108 379342 451154 379402
rect 453021 379400 453436 379402
rect 453021 379344 453026 379400
rect 453082 379344 453436 379400
rect 453021 379342 453436 379344
rect 451108 379340 451114 379342
rect 450997 379339 451063 379340
rect 453021 379339 453087 379342
rect 453430 379340 453436 379342
rect 453500 379340 453506 379404
rect 455505 379402 455571 379405
rect 458357 379404 458423 379405
rect 460933 379404 460999 379405
rect 455822 379402 455828 379404
rect 455505 379400 455828 379402
rect 455505 379344 455510 379400
rect 455566 379344 455828 379400
rect 455505 379342 455828 379344
rect 455505 379339 455571 379342
rect 455822 379340 455828 379342
rect 455892 379340 455898 379404
rect 458357 379400 458404 379404
rect 458468 379402 458474 379404
rect 458357 379344 458362 379400
rect 458357 379340 458404 379344
rect 458468 379342 458514 379402
rect 460933 379400 460980 379404
rect 461044 379402 461050 379404
rect 474825 379402 474891 379405
rect 475878 379402 475884 379404
rect 460933 379344 460938 379400
rect 458468 379340 458474 379342
rect 460933 379340 460980 379344
rect 461044 379342 461090 379402
rect 474825 379400 475884 379402
rect 474825 379344 474830 379400
rect 474886 379344 475884 379400
rect 474825 379342 475884 379344
rect 461044 379340 461050 379342
rect 458357 379339 458423 379340
rect 460933 379339 460999 379340
rect 474825 379339 474891 379342
rect 475878 379340 475884 379342
rect 475948 379340 475954 379404
rect 399477 379268 399543 379269
rect 400397 379268 400463 379269
rect 402973 379268 403039 379269
rect 409965 379268 410031 379269
rect 415853 379268 415919 379269
rect 325877 379208 325882 379264
rect 283484 379204 283490 379206
rect 325877 379204 325924 379208
rect 325988 379206 326034 379266
rect 393270 379206 398114 379266
rect 325988 379204 325994 379206
rect 283373 379203 283439 379204
rect 325877 379203 325943 379204
rect 78254 379130 78260 379132
rect 64830 379070 78260 379130
rect 78254 379068 78260 379070
rect 78324 379130 78330 379132
rect 205357 379130 205423 379133
rect 208393 379130 208459 379133
rect 209497 379130 209563 379133
rect 241830 379130 241836 379132
rect 78324 379128 205834 379130
rect 78324 379072 205362 379128
rect 205418 379072 205834 379128
rect 78324 379070 205834 379072
rect 78324 379068 78330 379070
rect 205357 379067 205423 379070
rect 47761 378994 47827 378997
rect 77201 378996 77267 378997
rect 94681 378996 94747 378997
rect 77150 378994 77156 378996
rect 47761 378992 64890 378994
rect 47761 378936 47766 378992
rect 47822 378936 64890 378992
rect 47761 378934 64890 378936
rect 77110 378934 77156 378994
rect 77220 378992 77267 378996
rect 94630 378994 94636 378996
rect 77262 378936 77267 378992
rect 47761 378931 47827 378934
rect 64830 378858 64890 378934
rect 77150 378932 77156 378934
rect 77220 378932 77267 378936
rect 77201 378931 77267 378932
rect 79550 378934 84210 378994
rect 94590 378934 94636 378994
rect 94700 378992 94747 378996
rect 94742 378936 94747 378992
rect 79550 378860 79610 378934
rect 83273 378860 83339 378861
rect 79542 378858 79548 378860
rect 64830 378798 79548 378858
rect 79542 378796 79548 378798
rect 79612 378796 79618 378860
rect 83222 378858 83228 378860
rect 83182 378798 83228 378858
rect 83292 378856 83339 378860
rect 83334 378800 83339 378856
rect 83222 378796 83228 378798
rect 83292 378796 83339 378800
rect 84150 378858 84210 378934
rect 94630 378932 94636 378934
rect 94700 378932 94747 378936
rect 148542 378932 148548 378996
rect 148612 378994 148618 378996
rect 148685 378994 148751 378997
rect 148612 378992 148751 378994
rect 148612 378936 148690 378992
rect 148746 378936 148751 378992
rect 148612 378934 148751 378936
rect 148612 378932 148618 378934
rect 94681 378931 94747 378932
rect 148685 378931 148751 378934
rect 183134 378932 183140 378996
rect 183204 378994 183210 378996
rect 183461 378994 183527 378997
rect 183204 378992 183527 378994
rect 183204 378936 183466 378992
rect 183522 378936 183527 378992
rect 183204 378934 183527 378936
rect 205774 378994 205834 379070
rect 208393 379128 241836 379130
rect 208393 379072 208398 379128
rect 208454 379072 209502 379128
rect 209558 379072 241836 379128
rect 208393 379070 241836 379072
rect 208393 379067 208459 379070
rect 209497 379067 209563 379070
rect 241830 379068 241836 379070
rect 241900 379068 241906 379132
rect 253105 379130 253171 379133
rect 370957 379130 371023 379133
rect 393270 379130 393330 379206
rect 398230 379204 398236 379268
rect 398300 379204 398306 379268
rect 399477 379264 399524 379268
rect 399588 379266 399594 379268
rect 399477 379208 399482 379264
rect 399477 379204 399524 379208
rect 399588 379206 399634 379266
rect 400397 379264 400444 379268
rect 400508 379266 400514 379268
rect 400397 379208 400402 379264
rect 399588 379204 399594 379206
rect 400397 379204 400444 379208
rect 400508 379206 400554 379266
rect 402973 379264 403020 379268
rect 403084 379266 403090 379268
rect 402973 379208 402978 379264
rect 400508 379204 400514 379206
rect 402973 379204 403020 379208
rect 403084 379206 403130 379266
rect 409965 379264 410012 379268
rect 410076 379266 410082 379268
rect 409965 379208 409970 379264
rect 403084 379204 403090 379206
rect 409965 379204 410012 379208
rect 410076 379206 410122 379266
rect 415853 379264 415900 379268
rect 415964 379266 415970 379268
rect 416865 379266 416931 379269
rect 416998 379266 417004 379268
rect 415853 379208 415858 379264
rect 410076 379204 410082 379206
rect 415853 379204 415900 379208
rect 415964 379206 416010 379266
rect 416865 379264 417004 379266
rect 416865 379208 416870 379264
rect 416926 379208 417004 379264
rect 416865 379206 417004 379208
rect 415964 379204 415970 379206
rect 253105 379128 393330 379130
rect 253105 379072 253110 379128
rect 253166 379072 370962 379128
rect 371018 379072 393330 379128
rect 253105 379070 393330 379072
rect 253105 379067 253171 379070
rect 370957 379067 371023 379070
rect 238150 378994 238156 378996
rect 205774 378934 238156 378994
rect 183204 378932 183210 378934
rect 183461 378931 183527 378934
rect 238150 378932 238156 378934
rect 238220 378994 238226 378996
rect 370865 378994 370931 378997
rect 398238 378994 398298 379204
rect 399477 379203 399543 379204
rect 400397 379203 400463 379204
rect 402973 379203 403039 379204
rect 409965 379203 410031 379204
rect 415853 379203 415919 379204
rect 416865 379203 416931 379206
rect 416998 379204 417004 379206
rect 417068 379204 417074 379268
rect 422845 379266 422911 379269
rect 463509 379268 463575 379269
rect 473445 379268 473511 379269
rect 503069 379268 503135 379269
rect 503529 379268 503595 379269
rect 423438 379266 423444 379268
rect 422845 379264 423444 379266
rect 422845 379208 422850 379264
rect 422906 379208 423444 379264
rect 422845 379206 423444 379208
rect 422845 379203 422911 379206
rect 423438 379204 423444 379206
rect 423508 379204 423514 379268
rect 463509 379264 463556 379268
rect 463620 379266 463626 379268
rect 463509 379208 463514 379264
rect 463509 379204 463556 379208
rect 463620 379206 463666 379266
rect 473445 379264 473492 379268
rect 473556 379266 473562 379268
rect 473445 379208 473450 379264
rect 463620 379204 463626 379206
rect 473445 379204 473492 379208
rect 473556 379206 473602 379266
rect 503069 379264 503116 379268
rect 503180 379266 503186 379268
rect 503069 379208 503074 379264
rect 473556 379204 473562 379206
rect 503069 379204 503116 379208
rect 503180 379206 503226 379266
rect 503180 379204 503186 379206
rect 503478 379204 503484 379268
rect 503548 379266 503595 379268
rect 503548 379264 503640 379266
rect 503590 379208 503640 379264
rect 503548 379206 503640 379208
rect 503548 379204 503595 379206
rect 463509 379203 463575 379204
rect 473445 379203 473511 379204
rect 503069 379203 503135 379204
rect 503529 379203 503595 379204
rect 238220 378992 398298 378994
rect 238220 378936 370870 378992
rect 370926 378936 398298 378992
rect 238220 378934 398298 378936
rect 465165 378994 465231 378997
rect 465942 378994 465948 378996
rect 465165 378992 465948 378994
rect 465165 378936 465170 378992
rect 465226 378936 465948 378992
rect 465165 378934 465948 378936
rect 238220 378932 238226 378934
rect 370865 378931 370931 378934
rect 465165 378931 465231 378934
rect 465942 378932 465948 378934
rect 466012 378932 466018 378996
rect 477585 378994 477651 378997
rect 478454 378994 478460 378996
rect 477585 378992 478460 378994
rect 477585 378936 477590 378992
rect 477646 378936 478460 378992
rect 477585 378934 478460 378936
rect 477585 378931 477651 378934
rect 478454 378932 478460 378934
rect 478524 378932 478530 378996
rect 206185 378858 206251 378861
rect 239254 378858 239260 378860
rect 84150 378856 239260 378858
rect 84150 378800 206190 378856
rect 206246 378800 239260 378856
rect 84150 378798 239260 378800
rect 83273 378795 83339 378796
rect 206185 378795 206251 378798
rect 239254 378796 239260 378798
rect 239324 378858 239330 378860
rect 372705 378858 372771 378861
rect 239324 378856 372771 378858
rect 239324 378800 372710 378856
rect 372766 378800 372771 378856
rect 239324 378798 372771 378800
rect 239324 378796 239330 378798
rect 372705 378795 372771 378798
rect 377622 378796 377628 378860
rect 377692 378858 377698 378860
rect 381261 378858 381327 378861
rect 427670 378858 427676 378860
rect 377692 378856 427676 378858
rect 377692 378800 381266 378856
rect 381322 378800 427676 378856
rect 377692 378798 427676 378800
rect 377692 378796 377698 378798
rect 381261 378795 381327 378798
rect 427670 378796 427676 378798
rect 427740 378796 427746 378860
rect 430665 378858 430731 378861
rect 430982 378858 430988 378860
rect 430665 378856 430988 378858
rect 430665 378800 430670 378856
rect 430726 378800 430988 378856
rect 430665 378798 430988 378800
rect 430665 378795 430731 378798
rect 430982 378796 430988 378798
rect 431052 378796 431058 378860
rect 470777 378858 470843 378861
rect 483381 378860 483447 378861
rect 470910 378858 470916 378860
rect 470777 378856 470916 378858
rect 470777 378800 470782 378856
rect 470838 378800 470916 378856
rect 470777 378798 470916 378800
rect 470777 378795 470843 378798
rect 470910 378796 470916 378798
rect 470980 378796 470986 378860
rect 483381 378856 483428 378860
rect 483492 378858 483498 378860
rect 483381 378800 483386 378856
rect 483381 378796 483428 378800
rect 483492 378798 483538 378858
rect 483492 378796 483498 378798
rect 483381 378795 483447 378796
rect 81934 378660 81940 378724
rect 82004 378722 82010 378724
rect 208393 378722 208459 378725
rect 82004 378720 208459 378722
rect 82004 378664 208398 378720
rect 208454 378664 208459 378720
rect 82004 378662 208459 378664
rect 82004 378660 82010 378662
rect 208393 378659 208459 378662
rect 209814 378660 209820 378724
rect 209884 378722 209890 378724
rect 210233 378722 210299 378725
rect 209884 378720 210299 378722
rect 209884 378664 210238 378720
rect 210294 378664 210299 378720
rect 209884 378662 210299 378664
rect 209884 378660 209890 378662
rect 210233 378659 210299 378662
rect 241462 378660 241468 378724
rect 241532 378722 241538 378724
rect 375097 378722 375163 378725
rect 375281 378722 375347 378725
rect 241532 378720 375347 378722
rect 241532 378664 375102 378720
rect 375158 378664 375286 378720
rect 375342 378664 375347 378720
rect 241532 378662 375347 378664
rect 241532 378660 241538 378662
rect 375097 378659 375163 378662
rect 375281 378659 375347 378662
rect 377806 378660 377812 378724
rect 377876 378722 377882 378724
rect 381077 378722 381143 378725
rect 433374 378722 433380 378724
rect 377876 378720 433380 378722
rect 377876 378664 381082 378720
rect 381138 378664 433380 378720
rect 377876 378662 433380 378664
rect 377876 378660 377882 378662
rect 381077 378659 381143 378662
rect 433374 378660 433380 378662
rect 433444 378660 433450 378724
rect 436185 378722 436251 378725
rect 436870 378722 436876 378724
rect 436185 378720 436876 378722
rect 436185 378664 436190 378720
rect 436246 378664 436876 378720
rect 436185 378662 436876 378664
rect 436185 378659 436251 378662
rect 436870 378660 436876 378662
rect 436940 378660 436946 378724
rect 467925 378722 467991 378725
rect 468518 378722 468524 378724
rect 467925 378720 468524 378722
rect 467925 378664 467930 378720
rect 467986 378664 468524 378720
rect 467925 378662 468524 378664
rect 467925 378659 467991 378662
rect 468518 378660 468524 378662
rect 468588 378660 468594 378724
rect 97022 378524 97028 378588
rect 97092 378586 97098 378588
rect 97809 378586 97875 378589
rect 97092 378584 97875 378586
rect 97092 378528 97814 378584
rect 97870 378528 97875 378584
rect 97092 378526 97875 378528
rect 97092 378524 97098 378526
rect 97809 378523 97875 378526
rect 100702 378524 100708 378588
rect 100772 378586 100778 378588
rect 100845 378586 100911 378589
rect 100772 378584 100911 378586
rect 100772 378528 100850 378584
rect 100906 378528 100911 378584
rect 100772 378526 100911 378528
rect 100772 378524 100778 378526
rect 100845 378523 100911 378526
rect 118182 378524 118188 378588
rect 118252 378586 118258 378588
rect 202965 378586 203031 378589
rect 118252 378584 203031 378586
rect 118252 378528 202970 378584
rect 203026 378528 203031 378584
rect 118252 378526 203031 378528
rect 118252 378524 118258 378526
rect 202965 378523 203031 378526
rect 207013 378586 207079 378589
rect 208209 378586 208275 378589
rect 218145 378586 218211 378589
rect 253565 378588 253631 378589
rect 255957 378588 256023 378589
rect 258349 378588 258415 378589
rect 260925 378588 260991 378589
rect 263593 378588 263659 378589
rect 207013 378584 253306 378586
rect 207013 378528 207018 378584
rect 207074 378528 208214 378584
rect 208270 378528 218150 378584
rect 218206 378528 253306 378584
rect 207013 378526 253306 378528
rect 207013 378523 207079 378526
rect 208209 378523 208275 378526
rect 218145 378523 218211 378526
rect 105302 378388 105308 378452
rect 105372 378450 105378 378452
rect 105721 378450 105787 378453
rect 105372 378448 105787 378450
rect 105372 378392 105726 378448
rect 105782 378392 105787 378448
rect 105372 378390 105787 378392
rect 105372 378388 105378 378390
rect 105721 378387 105787 378390
rect 182265 378450 182331 378453
rect 205357 378452 205423 378453
rect 183502 378450 183508 378452
rect 182265 378448 183508 378450
rect 182265 378392 182270 378448
rect 182326 378392 183508 378448
rect 182265 378390 183508 378392
rect 182265 378387 182331 378390
rect 183502 378388 183508 378390
rect 183572 378388 183578 378452
rect 205357 378450 205404 378452
rect 205312 378448 205404 378450
rect 205312 378392 205362 378448
rect 205312 378390 205404 378392
rect 205357 378388 205404 378390
rect 205468 378388 205474 378452
rect 241830 378388 241836 378452
rect 241900 378450 241906 378452
rect 253105 378450 253171 378453
rect 241900 378448 253171 378450
rect 241900 378392 253110 378448
rect 253166 378392 253171 378448
rect 241900 378390 253171 378392
rect 253246 378450 253306 378526
rect 253565 378584 253612 378588
rect 253676 378586 253682 378588
rect 253565 378528 253570 378584
rect 253565 378524 253612 378528
rect 253676 378526 253722 378586
rect 255957 378584 256004 378588
rect 256068 378586 256074 378588
rect 255957 378528 255962 378584
rect 253676 378524 253682 378526
rect 255957 378524 256004 378528
rect 256068 378526 256114 378586
rect 258349 378584 258396 378588
rect 258460 378586 258466 378588
rect 258349 378528 258354 378584
rect 256068 378524 256074 378526
rect 258349 378524 258396 378528
rect 258460 378526 258506 378586
rect 260925 378584 260972 378588
rect 261036 378586 261042 378588
rect 263542 378586 263548 378588
rect 260925 378528 260930 378584
rect 258460 378524 258466 378526
rect 260925 378524 260972 378528
rect 261036 378526 261082 378586
rect 263502 378526 263548 378586
rect 263612 378584 263659 378588
rect 263654 378528 263659 378584
rect 261036 378524 261042 378526
rect 263542 378524 263548 378526
rect 263612 378524 263659 378528
rect 253565 378523 253631 378524
rect 255957 378523 256023 378524
rect 258349 378523 258415 378524
rect 260925 378523 260991 378524
rect 263593 378523 263659 378524
rect 265893 378588 265959 378589
rect 265893 378584 265940 378588
rect 266004 378586 266010 378588
rect 268101 378586 268167 378589
rect 273437 378588 273503 378589
rect 320909 378588 320975 378589
rect 268326 378586 268332 378588
rect 265893 378528 265898 378584
rect 265893 378524 265940 378528
rect 266004 378526 266050 378586
rect 268101 378584 268332 378586
rect 268101 378528 268106 378584
rect 268162 378528 268332 378584
rect 268101 378526 268332 378528
rect 266004 378524 266010 378526
rect 265893 378523 265959 378524
rect 268101 378523 268167 378526
rect 268326 378524 268332 378526
rect 268396 378524 268402 378588
rect 273437 378584 273484 378588
rect 273548 378586 273554 378588
rect 273437 378528 273442 378584
rect 273437 378524 273484 378528
rect 273548 378526 273594 378586
rect 320909 378584 320956 378588
rect 321020 378586 321026 378588
rect 413277 378586 413343 378589
rect 414565 378588 414631 378589
rect 418429 378588 418495 378589
rect 413502 378586 413508 378588
rect 320909 378528 320914 378584
rect 273548 378524 273554 378526
rect 320909 378524 320956 378528
rect 321020 378526 321066 378586
rect 413277 378584 413508 378586
rect 413277 378528 413282 378584
rect 413338 378528 413508 378584
rect 413277 378526 413508 378528
rect 321020 378524 321026 378526
rect 273437 378523 273503 378524
rect 320909 378523 320975 378524
rect 413277 378523 413343 378526
rect 413502 378524 413508 378526
rect 413572 378524 413578 378588
rect 414565 378584 414612 378588
rect 414676 378586 414682 378588
rect 414565 378528 414570 378584
rect 414565 378524 414612 378528
rect 414676 378526 414722 378586
rect 418429 378584 418476 378588
rect 418540 378586 418546 378588
rect 418429 378528 418434 378584
rect 414676 378524 414682 378526
rect 418429 378524 418476 378528
rect 418540 378526 418586 378586
rect 418540 378524 418546 378526
rect 414565 378523 414631 378524
rect 418429 378523 418495 378524
rect 265525 378450 265591 378453
rect 253246 378448 265591 378450
rect 253246 378392 265530 378448
rect 265586 378392 265591 378448
rect 253246 378390 265591 378392
rect 241900 378388 241906 378390
rect 205357 378387 205423 378388
rect 253105 378387 253171 378390
rect 265525 378387 265591 378390
rect 343173 378452 343239 378453
rect 343173 378448 343220 378452
rect 343284 378450 343290 378452
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 343173 378392 343178 378448
rect 343173 378388 343220 378392
rect 343284 378390 343330 378450
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 343284 378388 343290 378390
rect 343173 378387 343239 378388
rect 580165 378387 580231 378390
rect 80421 378314 80487 378317
rect 208117 378314 208183 378317
rect 244273 378316 244339 378317
rect 240542 378314 240548 378316
rect 80421 378312 240548 378314
rect 80421 378256 80426 378312
rect 80482 378256 208122 378312
rect 208178 378256 240548 378312
rect 80421 378254 240548 378256
rect 80421 378251 80487 378254
rect 208117 378251 208183 378254
rect 240542 378252 240548 378254
rect 240612 378314 240618 378316
rect 241462 378314 241468 378316
rect 240612 378254 241468 378314
rect 240612 378252 240618 378254
rect 241462 378252 241468 378254
rect 241532 378252 241538 378316
rect 244222 378314 244228 378316
rect 244182 378254 244228 378314
rect 244292 378312 244339 378316
rect 244334 378256 244339 378312
rect 244222 378252 244228 378254
rect 244292 378252 244339 378256
rect 244273 378251 244339 378252
rect 250621 378316 250687 378317
rect 262765 378316 262831 378317
rect 266353 378316 266419 378317
rect 250621 378312 250668 378316
rect 250732 378314 250738 378316
rect 250621 378256 250626 378312
rect 250621 378252 250668 378256
rect 250732 378254 250778 378314
rect 262765 378312 262812 378316
rect 262876 378314 262882 378316
rect 266302 378314 266308 378316
rect 262765 378256 262770 378312
rect 250732 378252 250738 378254
rect 262765 378252 262812 378256
rect 262876 378254 262922 378314
rect 266262 378254 266308 378314
rect 266372 378312 266419 378316
rect 266414 378256 266419 378312
rect 262876 378252 262882 378254
rect 266302 378252 266308 378254
rect 266372 378252 266419 378256
rect 250621 378251 250687 378252
rect 262765 378251 262831 378252
rect 266353 378251 266419 378252
rect 267549 378316 267615 378317
rect 267549 378312 267596 378316
rect 267660 378314 267666 378316
rect 267549 378256 267554 378312
rect 267549 378252 267596 378256
rect 267660 378254 267706 378314
rect 267660 378252 267666 378254
rect 343398 378252 343404 378316
rect 343468 378314 343474 378316
rect 343541 378314 343607 378317
rect 343468 378312 343607 378314
rect 343468 378256 343546 378312
rect 343602 378256 343607 378312
rect 343468 378254 343607 378256
rect 343468 378252 343474 378254
rect 267549 378251 267615 378252
rect 343541 378251 343607 378254
rect 432229 378316 432295 378317
rect 432229 378312 432276 378316
rect 432340 378314 432346 378316
rect 432229 378256 432234 378312
rect 432229 378252 432276 378256
rect 432340 378254 432386 378314
rect 583520 378300 584960 378390
rect 432340 378252 432346 378254
rect 432229 378251 432295 378252
rect 84377 378180 84443 378181
rect 101857 378180 101923 378181
rect 106457 378180 106523 378181
rect 107561 378180 107627 378181
rect 84326 378178 84332 378180
rect 84286 378118 84332 378178
rect 84396 378176 84443 378180
rect 101806 378178 101812 378180
rect 84438 378120 84443 378176
rect 84326 378116 84332 378118
rect 84396 378116 84443 378120
rect 101766 378118 101812 378178
rect 101876 378176 101923 378180
rect 101918 378120 101923 378176
rect 101806 378116 101812 378118
rect 101876 378116 101923 378120
rect 104014 378116 104020 378180
rect 104084 378116 104090 378180
rect 106406 378178 106412 378180
rect 106366 378118 106412 378178
rect 106476 378176 106523 378180
rect 107510 378178 107516 378180
rect 106518 378120 106523 378176
rect 106406 378116 106412 378118
rect 106476 378116 106523 378120
rect 107470 378118 107516 378178
rect 107580 378176 107627 378180
rect 107622 378120 107627 378176
rect 107510 378116 107516 378118
rect 107580 378116 107627 378120
rect 117078 378116 117084 378180
rect 117148 378178 117154 378180
rect 208301 378178 208367 378181
rect 276013 378178 276079 378181
rect 117148 378176 276079 378178
rect 117148 378120 208306 378176
rect 208362 378120 276018 378176
rect 276074 378120 276079 378176
rect 117148 378118 276079 378120
rect 117148 378116 117154 378118
rect 84377 378115 84443 378116
rect 101857 378115 101923 378116
rect 57462 377980 57468 378044
rect 57532 378042 57538 378044
rect 59537 378042 59603 378045
rect 57532 378040 59603 378042
rect 57532 377984 59542 378040
rect 59598 377984 59603 378040
rect 57532 377982 59603 377984
rect 104022 378042 104082 378116
rect 106457 378115 106523 378116
rect 107561 378115 107627 378116
rect 208301 378115 208367 378118
rect 276013 378115 276079 378118
rect 377397 378180 377463 378181
rect 408677 378180 408743 378181
rect 418153 378180 418219 378181
rect 377397 378176 377444 378180
rect 377508 378178 377514 378180
rect 377397 378120 377402 378176
rect 377397 378116 377444 378120
rect 377508 378118 377554 378178
rect 408677 378176 408724 378180
rect 408788 378178 408794 378180
rect 418102 378178 418108 378180
rect 408677 378120 408682 378176
rect 377508 378116 377514 378118
rect 408677 378116 408724 378120
rect 408788 378118 408834 378178
rect 418062 378118 418108 378178
rect 418172 378176 418219 378180
rect 418214 378120 418219 378176
rect 408788 378116 408794 378118
rect 418102 378116 418108 378118
rect 418172 378116 418219 378120
rect 377397 378115 377463 378116
rect 408677 378115 408743 378116
rect 418153 378115 418219 378116
rect 420637 378180 420703 378181
rect 420637 378176 420684 378180
rect 420748 378178 420754 378180
rect 421189 378178 421255 378181
rect 421782 378178 421788 378180
rect 420637 378120 420642 378176
rect 420637 378116 420684 378120
rect 420748 378118 420794 378178
rect 421189 378176 421788 378178
rect 421189 378120 421194 378176
rect 421250 378120 421788 378176
rect 421189 378118 421788 378120
rect 420748 378116 420754 378118
rect 420637 378115 420703 378116
rect 421189 378115 421255 378118
rect 421782 378116 421788 378118
rect 421852 378116 421858 378180
rect 422661 378178 422727 378181
rect 423949 378180 424015 378181
rect 422886 378178 422892 378180
rect 422661 378176 422892 378178
rect 422661 378120 422666 378176
rect 422722 378120 422892 378176
rect 422661 378118 422892 378120
rect 422661 378115 422727 378118
rect 422886 378116 422892 378118
rect 422956 378116 422962 378180
rect 423949 378176 423996 378180
rect 424060 378178 424066 378180
rect 425145 378178 425211 378181
rect 428549 378180 428615 378181
rect 429653 378180 429719 378181
rect 439037 378180 439103 378181
rect 425278 378178 425284 378180
rect 423949 378120 423954 378176
rect 423949 378116 423996 378120
rect 424060 378118 424106 378178
rect 425145 378176 425284 378178
rect 425145 378120 425150 378176
rect 425206 378120 425284 378176
rect 425145 378118 425284 378120
rect 424060 378116 424066 378118
rect 423949 378115 424015 378116
rect 425145 378115 425211 378118
rect 425278 378116 425284 378118
rect 425348 378116 425354 378180
rect 428549 378176 428596 378180
rect 428660 378178 428666 378180
rect 428549 378120 428554 378176
rect 428549 378116 428596 378120
rect 428660 378118 428706 378178
rect 429653 378176 429700 378180
rect 429764 378178 429770 378180
rect 429653 378120 429658 378176
rect 428660 378116 428666 378118
rect 429653 378116 429700 378120
rect 429764 378118 429810 378178
rect 439037 378176 439084 378180
rect 439148 378178 439154 378180
rect 480662 378178 480668 378180
rect 439037 378120 439042 378176
rect 429764 378116 429770 378118
rect 439037 378116 439084 378120
rect 439148 378118 439194 378178
rect 480210 378118 480668 378178
rect 439148 378116 439154 378118
rect 428549 378115 428615 378116
rect 429653 378115 429719 378116
rect 439037 378115 439103 378116
rect 104022 377982 195990 378042
rect 57532 377980 57538 377982
rect 59537 377979 59603 377982
rect 195930 377906 195990 377982
rect 207054 377980 207060 378044
rect 207124 378042 207130 378044
rect 208301 378042 208367 378045
rect 207124 378040 208367 378042
rect 207124 377984 208306 378040
rect 208362 377984 208367 378040
rect 207124 377982 208367 377984
rect 207124 377980 207130 377982
rect 208301 377979 208367 377982
rect 211654 377980 211660 378044
rect 211724 378042 211730 378044
rect 212441 378042 212507 378045
rect 211724 378040 212507 378042
rect 211724 377984 212446 378040
rect 212502 377984 212507 378040
rect 211724 377982 212507 377984
rect 211724 377980 211730 377982
rect 212441 377979 212507 377982
rect 213678 377980 213684 378044
rect 213748 378042 213754 378044
rect 213821 378042 213887 378045
rect 213748 378040 213887 378042
rect 213748 377984 213826 378040
rect 213882 377984 213887 378040
rect 213748 377982 213887 377984
rect 213748 377980 213754 377982
rect 213821 377979 213887 377982
rect 214046 377980 214052 378044
rect 214116 378042 214122 378044
rect 215201 378042 215267 378045
rect 214116 378040 215267 378042
rect 214116 377984 215206 378040
rect 215262 377984 215267 378040
rect 214116 377982 215267 377984
rect 214116 377980 214122 377982
rect 215201 377979 215267 377982
rect 360142 377980 360148 378044
rect 360212 378042 360218 378044
rect 361481 378042 361547 378045
rect 360212 378040 361547 378042
rect 360212 377984 361486 378040
rect 361542 377984 361547 378040
rect 360212 377982 361547 377984
rect 360212 377980 360218 377982
rect 361481 377979 361547 377982
rect 363505 378042 363571 378045
rect 480210 378042 480270 378118
rect 480662 378116 480668 378118
rect 480732 378116 480738 378180
rect 363505 378040 480270 378042
rect 363505 377984 363510 378040
rect 363566 377984 480270 378040
rect 363505 377982 480270 377984
rect 363505 377979 363571 377982
rect 215477 377906 215543 377909
rect 217961 377906 218027 377909
rect 219893 377906 219959 377909
rect 195930 377904 219959 377906
rect 195930 377848 215482 377904
rect 215538 377848 217966 377904
rect 218022 377848 219898 377904
rect 219954 377848 219959 377904
rect 195930 377846 219959 377848
rect 215477 377843 215543 377846
rect 217961 377843 218027 377846
rect 219893 377843 219959 377846
rect 370078 377844 370084 377908
rect 370148 377906 370154 377908
rect 371141 377906 371207 377909
rect 370148 377904 371207 377906
rect 370148 377848 371146 377904
rect 371202 377848 371207 377904
rect 370148 377846 371207 377848
rect 370148 377844 370154 377846
rect 371141 377843 371207 377846
rect 213862 376620 213868 376684
rect 213932 376682 213938 376684
rect 215109 376682 215175 376685
rect 213932 376680 215175 376682
rect 213932 376624 215114 376680
rect 215170 376624 215175 376680
rect 213932 376622 215175 376624
rect 213932 376620 213938 376622
rect 215109 376619 215175 376622
rect 359958 376620 359964 376684
rect 360028 376682 360034 376684
rect 465165 376682 465231 376685
rect 360028 376680 465231 376682
rect 360028 376624 465170 376680
rect 465226 376624 465231 376680
rect 360028 376622 465231 376624
rect 360028 376620 360034 376622
rect 465165 376619 465231 376622
rect 214465 376546 214531 376549
rect 216622 376546 216628 376548
rect 214465 376544 216628 376546
rect 214465 376488 214470 376544
rect 214526 376488 216628 376544
rect 214465 376486 216628 376488
rect 214465 376483 214531 376486
rect 216622 376484 216628 376486
rect 216692 376484 216698 376548
rect 214005 376274 214071 376277
rect 214005 376272 215310 376274
rect 214005 376216 214010 376272
rect 214066 376216 215310 376272
rect 214005 376214 215310 376216
rect 214005 376211 214071 376214
rect 215250 376002 215310 376214
rect 216990 376002 216996 376004
rect 215250 375942 216996 376002
rect 216990 375940 216996 375942
rect 217060 376002 217066 376004
rect 239121 376002 239187 376005
rect 217060 376000 239187 376002
rect 217060 375944 239126 376000
rect 239182 375944 239187 376000
rect 217060 375942 239187 375944
rect 217060 375940 217066 375942
rect 239121 375939 239187 375942
rect 215334 375396 215340 375460
rect 215404 375458 215410 375460
rect 216581 375458 216647 375461
rect 215404 375456 216647 375458
rect 215404 375400 216586 375456
rect 216642 375400 216647 375456
rect 215404 375398 216647 375400
rect 215404 375396 215410 375398
rect 216581 375395 216647 375398
rect 376753 374916 376819 374917
rect 376702 374914 376708 374916
rect 376662 374854 376708 374914
rect 376772 374912 376819 374916
rect 376814 374856 376819 374912
rect 376702 374852 376708 374854
rect 376772 374852 376819 374856
rect 376753 374851 376819 374852
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect 178585 358868 178651 358869
rect 178534 358866 178540 358868
rect 178494 358806 178540 358866
rect 178604 358864 178651 358868
rect 178646 358808 178651 358864
rect 178534 358804 178540 358806
rect 178604 358804 178651 358808
rect 179638 358804 179644 358868
rect 179708 358866 179714 358868
rect 180149 358866 180215 358869
rect 190913 358868 190979 358869
rect 338481 358868 338547 358869
rect 190862 358866 190868 358868
rect 179708 358864 180215 358866
rect 179708 358808 180154 358864
rect 180210 358808 180215 358864
rect 179708 358806 180215 358808
rect 190822 358806 190868 358866
rect 190932 358864 190979 358868
rect 338430 358866 338436 358868
rect 190974 358808 190979 358864
rect 179708 358804 179714 358806
rect 178585 358803 178651 358804
rect 180149 358803 180215 358806
rect 190862 358804 190868 358806
rect 190932 358804 190979 358808
rect 338390 358806 338436 358866
rect 338500 358864 338547 358868
rect 338542 358808 338547 358864
rect 338430 358804 338436 358806
rect 338500 358804 338547 358808
rect 339718 358804 339724 358868
rect 339788 358866 339794 358868
rect 340045 358866 340111 358869
rect 339788 358864 340111 358866
rect 339788 358808 340050 358864
rect 340106 358808 340111 358864
rect 339788 358806 340111 358808
rect 339788 358804 339794 358806
rect 190913 358803 190979 358804
rect 338481 358803 338547 358804
rect 340045 358803 340111 358806
rect 350942 358804 350948 358868
rect 351012 358866 351018 358868
rect 351729 358866 351795 358869
rect 351012 358864 351795 358866
rect 351012 358808 351734 358864
rect 351790 358808 351795 358864
rect 351012 358806 351795 358808
rect 351012 358804 351018 358806
rect 351729 358803 351795 358806
rect 498510 358804 498516 358868
rect 498580 358866 498586 358868
rect 498929 358866 498995 358869
rect 498580 358864 498995 358866
rect 498580 358808 498934 358864
rect 498990 358808 498995 358864
rect 498580 358806 498995 358808
rect 498580 358804 498586 358806
rect 498929 358803 498995 358806
rect 499798 358804 499804 358868
rect 499868 358866 499874 358868
rect 500401 358866 500467 358869
rect 510889 358868 510955 358869
rect 510838 358866 510844 358868
rect 499868 358864 500467 358866
rect 499868 358808 500406 358864
rect 500462 358808 500467 358864
rect 499868 358806 500467 358808
rect 510798 358806 510844 358866
rect 510908 358864 510955 358868
rect 510950 358808 510955 358864
rect 499868 358804 499874 358806
rect 500401 358803 500467 358806
rect 510838 358804 510844 358806
rect 510908 358804 510955 358808
rect 510889 358803 510955 358804
rect -960 358458 480 358548
rect 3693 358458 3759 358461
rect -960 358456 3759 358458
rect -960 358400 3698 358456
rect 3754 358400 3759 358456
rect -960 358398 3759 358400
rect -960 358308 480 358398
rect 3693 358395 3759 358398
rect 377990 357308 377996 357372
rect 378060 357370 378066 357372
rect 379513 357370 379579 357373
rect 378060 357368 379579 357370
rect 378060 357312 379518 357368
rect 379574 357312 379579 357368
rect 378060 357310 379579 357312
rect 378060 357308 378066 357310
rect 379513 357307 379579 357310
rect 196558 353154 196618 353190
rect 199009 353154 199075 353157
rect 196558 353152 199075 353154
rect 196558 353096 199014 353152
rect 199070 353096 199075 353152
rect 196558 353094 199075 353096
rect 356562 353154 356622 353190
rect 358905 353154 358971 353157
rect 356562 353152 358971 353154
rect 356562 353096 358910 353152
rect 358966 353096 358971 353152
rect 356562 353094 358971 353096
rect 199009 353091 199075 353094
rect 358905 353091 358971 353094
rect 516558 352882 516618 353190
rect 519261 352882 519327 352885
rect 519445 352882 519511 352885
rect 516558 352880 519511 352882
rect 516558 352824 519266 352880
rect 519322 352824 519450 352880
rect 519506 352824 519511 352880
rect 516558 352822 519511 352824
rect 519261 352819 519327 352822
rect 519445 352819 519511 352822
rect 198825 351930 198891 351933
rect 199009 351930 199075 351933
rect 198825 351928 199075 351930
rect 198825 351872 198830 351928
rect 198886 351872 199014 351928
rect 199070 351872 199075 351928
rect 198825 351870 199075 351872
rect 198825 351867 198891 351870
rect 199009 351867 199075 351870
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 57605 311130 57671 311133
rect 57605 311128 60062 311130
rect 57605 311072 57610 311128
rect 57666 311072 60062 311128
rect 57605 311070 60062 311072
rect 57605 311067 57671 311070
rect 60002 310894 60062 311070
rect 217869 310994 217935 310997
rect 217869 310992 219450 310994
rect 217869 310936 217874 310992
rect 217930 310936 219450 310992
rect 217869 310934 219450 310936
rect 217869 310931 217935 310934
rect 219390 310924 219450 310934
rect 219390 310864 220064 310924
rect 379838 310864 380052 310924
rect 377397 310858 377463 310861
rect 377765 310858 377831 310861
rect 379838 310858 379898 310864
rect 377397 310856 379898 310858
rect 377397 310800 377402 310856
rect 377458 310800 377770 310856
rect 377826 310800 379898 310856
rect 377397 310798 379898 310800
rect 377397 310795 377463 310798
rect 377765 310795 377831 310798
rect 216857 310042 216923 310045
rect 217041 310042 217107 310045
rect 377213 310042 377279 310045
rect 377949 310042 378015 310045
rect 216857 310040 219450 310042
rect 216857 309984 216862 310040
rect 216918 309984 217046 310040
rect 217102 309984 219450 310040
rect 216857 309982 219450 309984
rect 216857 309979 216923 309982
rect 217041 309979 217107 309982
rect 219390 309972 219450 309982
rect 377213 310040 379898 310042
rect 377213 309984 377218 310040
rect 377274 309984 377954 310040
rect 378010 309984 379898 310040
rect 377213 309982 379898 309984
rect 377213 309979 377279 309982
rect 377949 309979 378015 309982
rect 379838 309972 379898 309982
rect 56869 309906 56935 309909
rect 57881 309906 57947 309909
rect 60002 309906 60062 309942
rect 219390 309912 220064 309972
rect 379838 309912 380052 309972
rect 56869 309904 60062 309906
rect 56869 309848 56874 309904
rect 56930 309848 57886 309904
rect 57942 309848 60062 309904
rect 56869 309846 60062 309848
rect 56869 309843 56935 309846
rect 57881 309843 57947 309846
rect 57421 309090 57487 309093
rect 57789 309090 57855 309093
rect 57421 309088 57855 309090
rect 57421 309032 57426 309088
rect 57482 309032 57794 309088
rect 57850 309032 57855 309088
rect 57421 309030 57855 309032
rect 57421 309027 57487 309030
rect 57789 309027 57855 309030
rect 57421 307866 57487 307869
rect 217593 307866 217659 307869
rect 376845 307866 376911 307869
rect 57421 307864 59922 307866
rect 57421 307808 57426 307864
rect 57482 307808 59922 307864
rect 57421 307806 59922 307808
rect 57421 307803 57487 307806
rect 59862 307796 59922 307806
rect 217593 307864 219450 307866
rect 217593 307808 217598 307864
rect 217654 307808 219450 307864
rect 217593 307806 219450 307808
rect 217593 307803 217659 307806
rect 219390 307796 219450 307806
rect 376845 307864 379898 307866
rect 376845 307808 376850 307864
rect 376906 307808 379898 307864
rect 376845 307806 379898 307808
rect 376845 307803 376911 307806
rect 379838 307796 379898 307806
rect 59862 307736 60032 307796
rect 219390 307736 220064 307796
rect 379838 307736 380052 307796
rect 376937 307730 377003 307733
rect 377857 307730 377923 307733
rect 376937 307728 377923 307730
rect 376937 307672 376942 307728
rect 376998 307672 377862 307728
rect 377918 307672 377923 307728
rect 376937 307670 377923 307672
rect 376937 307667 377003 307670
rect 377857 307667 377923 307670
rect 377857 306914 377923 306917
rect 377857 306912 379898 306914
rect 377857 306856 377862 306912
rect 377918 306856 379898 306912
rect 377857 306854 379898 306856
rect 377857 306851 377923 306854
rect 379838 306844 379898 306854
rect 57697 306778 57763 306781
rect 60002 306778 60062 306814
rect 219390 306784 220064 306844
rect 379838 306784 380052 306844
rect 57697 306776 60062 306778
rect 57697 306720 57702 306776
rect 57758 306720 60062 306776
rect 57697 306718 60062 306720
rect 217685 306778 217751 306781
rect 219390 306778 219450 306784
rect 217685 306776 219450 306778
rect 217685 306720 217690 306776
rect 217746 306720 219450 306776
rect 217685 306718 219450 306720
rect 57697 306715 57763 306718
rect 217685 306715 217751 306718
rect -960 306234 480 306324
rect 3601 306234 3667 306237
rect -960 306232 3667 306234
rect -960 306176 3606 306232
rect 3662 306176 3667 306232
rect -960 306174 3667 306176
rect -960 306084 480 306174
rect 3601 306171 3667 306174
rect 57513 305010 57579 305013
rect 57789 305010 57855 305013
rect 60002 305010 60062 305046
rect 219390 305016 220064 305076
rect 379838 305016 380052 305076
rect 57513 305008 60062 305010
rect 57513 304952 57518 305008
rect 57574 304952 57794 305008
rect 57850 304952 60062 305008
rect 57513 304950 60062 304952
rect 217777 305010 217843 305013
rect 219390 305010 219450 305016
rect 217777 305008 219450 305010
rect 217777 304952 217782 305008
rect 217838 304952 219450 305008
rect 217777 304950 219450 304952
rect 377581 305010 377647 305013
rect 379838 305010 379898 305016
rect 377581 305008 379898 305010
rect 377581 304952 377586 305008
rect 377642 304952 379898 305008
rect 377581 304950 379898 304952
rect 57513 304947 57579 304950
rect 57789 304947 57855 304950
rect 217777 304947 217843 304950
rect 377581 304947 377647 304950
rect 57513 303650 57579 303653
rect 60002 303650 60062 303958
rect 219390 303928 220064 303988
rect 379838 303928 380052 303988
rect 216949 303922 217015 303925
rect 217501 303922 217567 303925
rect 219390 303922 219450 303928
rect 216949 303920 219450 303922
rect 216949 303864 216954 303920
rect 217010 303864 217506 303920
rect 217562 303864 219450 303920
rect 216949 303862 219450 303864
rect 377857 303922 377923 303925
rect 379838 303922 379898 303928
rect 377857 303920 379898 303922
rect 377857 303864 377862 303920
rect 377918 303864 379898 303920
rect 377857 303862 379898 303864
rect 216949 303859 217015 303862
rect 217501 303859 217567 303862
rect 377857 303859 377923 303862
rect 57513 303648 60062 303650
rect 57513 303592 57518 303648
rect 57574 303592 60062 303648
rect 57513 303590 60062 303592
rect 57513 303587 57579 303590
rect 56777 301610 56843 301613
rect 60002 301610 60062 302190
rect 219390 302160 220064 302220
rect 379838 302160 380052 302220
rect 216949 302154 217015 302157
rect 217317 302154 217383 302157
rect 219390 302154 219450 302160
rect 216949 302152 219450 302154
rect 216949 302096 216954 302152
rect 217010 302096 217322 302152
rect 217378 302096 219450 302152
rect 216949 302094 219450 302096
rect 377305 302154 377371 302157
rect 378041 302154 378107 302157
rect 379838 302154 379898 302160
rect 377305 302152 379898 302154
rect 377305 302096 377310 302152
rect 377366 302096 378046 302152
rect 378102 302096 379898 302152
rect 377305 302094 379898 302096
rect 216949 302091 217015 302094
rect 217317 302091 217383 302094
rect 377305 302091 377371 302094
rect 378041 302091 378107 302094
rect 56777 301608 60062 301610
rect 56777 301552 56782 301608
rect 56838 301552 60062 301608
rect 56777 301550 60062 301552
rect 56777 301547 56843 301550
rect 583520 298604 584960 298844
rect 519353 293858 519419 293861
rect 516558 293856 519419 293858
rect 516558 293800 519358 293856
rect 519414 293800 519419 293856
rect 516558 293798 519419 293800
rect 516558 293350 516618 293798
rect 519353 293795 519419 293798
rect -960 293028 480 293268
rect 196558 292770 196618 293350
rect 199285 292770 199351 292773
rect 199561 292770 199627 292773
rect 196558 292768 199627 292770
rect 196558 292712 199290 292768
rect 199346 292712 199566 292768
rect 199622 292712 199627 292768
rect 196558 292710 199627 292712
rect 356562 292770 356622 293350
rect 359273 292770 359339 292773
rect 359549 292770 359615 292773
rect 356562 292768 359615 292770
rect 356562 292712 359278 292768
rect 359334 292712 359554 292768
rect 359610 292712 359615 292768
rect 356562 292710 359615 292712
rect 199285 292707 199351 292710
rect 199561 292707 199627 292710
rect 359273 292707 359339 292710
rect 359549 292707 359615 292710
rect 518893 292498 518959 292501
rect 519629 292498 519695 292501
rect 516558 292496 519695 292498
rect 516558 292440 518898 292496
rect 518954 292440 519634 292496
rect 519690 292440 519695 292496
rect 516558 292438 519695 292440
rect 359089 291818 359155 291821
rect 359641 291818 359707 291821
rect 356562 291816 359707 291818
rect 356562 291760 359094 291816
rect 359150 291760 359646 291816
rect 359702 291760 359707 291816
rect 356562 291758 359707 291760
rect 356562 291718 356622 291758
rect 359089 291755 359155 291758
rect 359641 291755 359707 291758
rect 516558 291718 516618 292438
rect 518893 292435 518959 292438
rect 519629 292435 519695 292438
rect 196558 291682 196618 291718
rect 199009 291682 199075 291685
rect 199469 291682 199535 291685
rect 196558 291680 199535 291682
rect 196558 291624 199014 291680
rect 199070 291624 199474 291680
rect 199530 291624 199535 291680
rect 196558 291622 199535 291624
rect 199009 291619 199075 291622
rect 199469 291619 199535 291622
rect 199193 291002 199259 291005
rect 199745 291002 199811 291005
rect 358997 291002 359063 291005
rect 359365 291002 359431 291005
rect 196558 291000 199811 291002
rect 196558 290944 199198 291000
rect 199254 290944 199750 291000
rect 199806 290944 199811 291000
rect 196558 290942 199811 290944
rect 196558 290358 196618 290942
rect 199193 290939 199259 290942
rect 199745 290939 199811 290942
rect 356562 291000 359431 291002
rect 356562 290944 359002 291000
rect 359058 290944 359370 291000
rect 359426 290944 359431 291000
rect 356562 290942 359431 290944
rect 356562 290358 356622 290942
rect 358997 290939 359063 290942
rect 359365 290939 359431 290942
rect 516558 290322 516618 290358
rect 519537 290322 519603 290325
rect 516558 290320 519603 290322
rect 516558 290264 519542 290320
rect 519598 290264 519603 290320
rect 516558 290262 519603 290264
rect 519537 290259 519603 290262
rect 198733 289778 198799 289781
rect 199377 289778 199443 289781
rect 198733 289776 199443 289778
rect 198733 289720 198738 289776
rect 198794 289720 199382 289776
rect 199438 289720 199443 289776
rect 198733 289718 199443 289720
rect 198733 289715 198799 289718
rect 199377 289715 199443 289718
rect 358997 289778 359063 289781
rect 359457 289778 359523 289781
rect 358997 289776 359523 289778
rect 358997 289720 359002 289776
rect 359058 289720 359462 289776
rect 359518 289720 359523 289776
rect 358997 289718 359523 289720
rect 358997 289715 359063 289718
rect 359457 289715 359523 289718
rect 196558 288826 196618 288862
rect 198733 288826 198799 288829
rect 196558 288824 198799 288826
rect 196558 288768 198738 288824
rect 198794 288768 198799 288824
rect 196558 288766 198799 288768
rect 356562 288826 356622 288862
rect 358997 288826 359063 288829
rect 356562 288824 359063 288826
rect 356562 288768 359002 288824
rect 359058 288768 359063 288824
rect 356562 288766 359063 288768
rect 516558 288826 516618 288862
rect 519169 288826 519235 288829
rect 520181 288826 520247 288829
rect 516558 288824 520247 288826
rect 516558 288768 519174 288824
rect 519230 288768 520186 288824
rect 520242 288768 520247 288824
rect 516558 288766 520247 288768
rect 198733 288763 198799 288766
rect 358997 288763 359063 288766
rect 519169 288763 519235 288766
rect 520181 288763 520247 288766
rect 199101 288418 199167 288421
rect 199653 288418 199719 288421
rect 199101 288416 199719 288418
rect 199101 288360 199106 288416
rect 199162 288360 199658 288416
rect 199714 288360 199719 288416
rect 199101 288358 199719 288360
rect 199101 288355 199167 288358
rect 199653 288355 199719 288358
rect 196558 287602 196618 287638
rect 199101 287602 199167 287605
rect 196558 287600 199167 287602
rect 196558 287544 199106 287600
rect 199162 287544 199167 287600
rect 196558 287542 199167 287544
rect 356562 287602 356622 287638
rect 359181 287602 359247 287605
rect 356562 287600 359247 287602
rect 356562 287544 359186 287600
rect 359242 287544 359247 287600
rect 356562 287542 359247 287544
rect 516558 287602 516618 287638
rect 518985 287602 519051 287605
rect 516558 287600 519051 287602
rect 516558 287544 518990 287600
rect 519046 287544 519051 287600
rect 516558 287542 519051 287544
rect 199101 287539 199167 287542
rect 359181 287539 359247 287542
rect 518985 287539 519051 287542
rect 583520 285276 584960 285516
rect 58617 284202 58683 284205
rect 58617 284200 60062 284202
rect 58617 284144 58622 284200
rect 58678 284144 60062 284200
rect 58617 284142 60062 284144
rect 58617 284139 58683 284142
rect 60002 283966 60062 284142
rect 216673 284066 216739 284069
rect 376845 284066 376911 284069
rect 216673 284064 219450 284066
rect 216673 284008 216678 284064
rect 216734 284008 219450 284064
rect 216673 284006 219450 284008
rect 216673 284003 216739 284006
rect 219390 283996 219450 284006
rect 376845 284064 379530 284066
rect 376845 284008 376850 284064
rect 376906 284008 379530 284064
rect 376845 284006 379530 284008
rect 376845 284003 376911 284006
rect 379470 283996 379530 284006
rect 219390 283936 220064 283996
rect 379470 283936 380052 283996
rect 57237 282570 57303 282573
rect 57881 282570 57947 282573
rect 57237 282568 60062 282570
rect 57237 282512 57242 282568
rect 57298 282512 57886 282568
rect 57942 282512 60062 282568
rect 57237 282510 60062 282512
rect 57237 282507 57303 282510
rect 57881 282507 57947 282510
rect 60002 282334 60062 282510
rect 219390 282304 220064 282364
rect 379470 282304 380052 282364
rect 51574 282236 51580 282300
rect 51644 282298 51650 282300
rect 52361 282298 52427 282301
rect 51644 282296 52427 282298
rect 51644 282240 52366 282296
rect 52422 282240 52427 282296
rect 51644 282238 52427 282240
rect 51644 282236 51650 282238
rect 52361 282235 52427 282238
rect 216673 282298 216739 282301
rect 219390 282298 219450 282304
rect 216673 282296 219450 282298
rect 216673 282240 216678 282296
rect 216734 282240 219450 282296
rect 216673 282238 219450 282240
rect 376937 282298 377003 282301
rect 379470 282298 379530 282304
rect 376937 282296 379530 282298
rect 376937 282240 376942 282296
rect 376998 282240 379530 282296
rect 376937 282238 379530 282240
rect 216673 282235 216739 282238
rect 376937 282235 377003 282238
rect 216765 282162 216831 282165
rect 377581 282162 377647 282165
rect 216765 282160 219450 282162
rect 216765 282104 216770 282160
rect 216826 282104 219450 282160
rect 216765 282102 219450 282104
rect 216765 282099 216831 282102
rect 219390 282092 219450 282102
rect 377581 282160 379530 282162
rect 377581 282104 377586 282160
rect 377642 282104 379530 282160
rect 377581 282102 379530 282104
rect 377581 282099 377647 282102
rect 379470 282092 379530 282102
rect 58709 282026 58775 282029
rect 60002 282026 60062 282062
rect 219390 282032 220064 282092
rect 379470 282032 380052 282092
rect 58709 282024 60062 282026
rect 58709 281968 58714 282024
rect 58770 281968 60062 282024
rect 58709 281966 60062 281968
rect 58709 281963 58775 281966
rect -960 279972 480 280212
rect 113357 273868 113423 273869
rect 426433 273868 426499 273869
rect 113312 273804 113318 273868
rect 113382 273866 113423 273868
rect 113382 273864 113474 273866
rect 113418 273808 113474 273864
rect 113382 273806 113474 273808
rect 113382 273804 113423 273806
rect 426376 273804 426382 273868
rect 426446 273866 426499 273868
rect 426446 273864 426538 273866
rect 426494 273808 426538 273864
rect 426446 273806 426538 273808
rect 426446 273804 426499 273806
rect 113357 273803 113423 273804
rect 426433 273803 426499 273804
rect 133413 273732 133479 273733
rect 133413 273730 133446 273732
rect 133354 273728 133446 273730
rect 133354 273672 133418 273728
rect 133354 273670 133446 273672
rect 133413 273668 133446 273670
rect 133510 273668 133516 273732
rect 133413 273667 133479 273668
rect 135897 273596 135963 273597
rect 138473 273596 138539 273597
rect 140865 273596 140931 273597
rect 143533 273596 143599 273597
rect 135888 273532 135894 273596
rect 135958 273594 135964 273596
rect 138472 273594 138478 273596
rect 135958 273534 136050 273594
rect 138386 273534 138478 273594
rect 135958 273532 135964 273534
rect 138472 273532 138478 273534
rect 138542 273532 138548 273596
rect 140865 273594 140926 273596
rect 140834 273592 140926 273594
rect 140834 273536 140870 273592
rect 140834 273534 140926 273536
rect 140865 273532 140926 273534
rect 140990 273532 140996 273596
rect 143504 273532 143510 273596
rect 143574 273594 143599 273596
rect 145925 273596 145991 273597
rect 266353 273596 266419 273597
rect 283465 273596 283531 273597
rect 421097 273596 421163 273597
rect 145925 273594 145958 273596
rect 143574 273592 143666 273594
rect 143594 273536 143666 273592
rect 143574 273534 143666 273536
rect 145866 273592 145958 273594
rect 145866 273536 145930 273592
rect 145866 273534 145958 273536
rect 143574 273532 143599 273534
rect 135897 273531 135963 273532
rect 138473 273531 138539 273532
rect 140865 273531 140931 273532
rect 143533 273531 143599 273532
rect 145925 273532 145958 273534
rect 146022 273532 146028 273596
rect 266353 273594 266382 273596
rect 266290 273592 266382 273594
rect 266290 273536 266358 273592
rect 266290 273534 266382 273536
rect 266353 273532 266382 273534
rect 266446 273532 266452 273596
rect 283465 273594 283518 273596
rect 283426 273592 283518 273594
rect 283426 273536 283470 273592
rect 283426 273534 283518 273536
rect 283465 273532 283518 273534
rect 283582 273532 283588 273596
rect 421072 273532 421078 273596
rect 421142 273594 421163 273596
rect 431125 273596 431191 273597
rect 433333 273596 433399 273597
rect 431125 273594 431142 273596
rect 421142 273592 421234 273594
rect 421158 273536 421234 273592
rect 421142 273534 421234 273536
rect 431050 273592 431142 273594
rect 431050 273536 431130 273592
rect 431050 273534 431142 273536
rect 421142 273532 421163 273534
rect 145925 273531 145991 273532
rect 266353 273531 266419 273532
rect 283465 273531 283531 273532
rect 421097 273531 421163 273532
rect 431125 273532 431142 273534
rect 431206 273532 431212 273596
rect 433312 273532 433318 273596
rect 433382 273594 433399 273596
rect 453389 273596 453455 273597
rect 453389 273594 453446 273596
rect 433382 273592 433474 273594
rect 433394 273536 433474 273592
rect 433382 273534 433474 273536
rect 453354 273592 453446 273594
rect 453354 273536 453394 273592
rect 453354 273534 453446 273536
rect 433382 273532 433399 273534
rect 431125 273531 431191 273532
rect 433333 273531 433399 273532
rect 453389 273532 453446 273534
rect 453510 273532 453516 273596
rect 453389 273531 453455 273532
rect 218421 273458 218487 273461
rect 273253 273460 273319 273461
rect 430941 273460 431007 273461
rect 218830 273458 218836 273460
rect 218421 273456 218836 273458
rect 218421 273400 218426 273456
rect 218482 273400 218836 273456
rect 218421 273398 218836 273400
rect 218421 273395 218487 273398
rect 218830 273396 218836 273398
rect 218900 273396 218906 273460
rect 273253 273458 273300 273460
rect 273208 273456 273300 273458
rect 273208 273400 273258 273456
rect 273208 273398 273300 273400
rect 273253 273396 273300 273398
rect 273364 273396 273370 273460
rect 430941 273458 430988 273460
rect 430896 273456 430988 273458
rect 430896 273400 430946 273456
rect 430896 273398 430988 273400
rect 430941 273396 430988 273398
rect 431052 273396 431058 273460
rect 273253 273395 273319 273396
rect 430941 273395 431007 273396
rect 57462 273260 57468 273324
rect 57532 273322 57538 273324
rect 61561 273322 61627 273325
rect 57532 273320 61627 273322
rect 57532 273264 61566 273320
rect 61622 273264 61627 273320
rect 57532 273262 61627 273264
rect 57532 273260 57538 273262
rect 61561 273259 61627 273262
rect 199510 273260 199516 273324
rect 199580 273322 199586 273324
rect 250662 273322 250668 273324
rect 199580 273262 250668 273322
rect 199580 273260 199586 273262
rect 250662 273260 250668 273262
rect 250732 273260 250738 273324
rect 371693 273322 371759 273325
rect 376886 273322 376892 273324
rect 371693 273320 376892 273322
rect 371693 273264 371698 273320
rect 371754 273264 376892 273320
rect 371693 273262 376892 273264
rect 371693 273259 371759 273262
rect 376886 273260 376892 273262
rect 376956 273322 376962 273324
rect 377806 273322 377812 273324
rect 376956 273262 377812 273322
rect 376956 273260 376962 273262
rect 377806 273260 377812 273262
rect 377876 273260 377882 273324
rect 378174 273260 378180 273324
rect 378244 273322 378250 273324
rect 378501 273322 378567 273325
rect 378244 273320 378567 273322
rect 378244 273264 378506 273320
rect 378562 273264 378567 273320
rect 378244 273262 378567 273264
rect 378244 273260 378250 273262
rect 378501 273259 378567 273262
rect 76005 273188 76071 273189
rect 77109 273188 77175 273189
rect 82997 273188 83063 273189
rect 90725 273188 90791 273189
rect 93669 273188 93735 273189
rect 95877 273188 95943 273189
rect 76005 273186 76052 273188
rect 75960 273184 76052 273186
rect 75960 273128 76010 273184
rect 75960 273126 76052 273128
rect 76005 273124 76052 273126
rect 76116 273124 76122 273188
rect 77109 273186 77156 273188
rect 77064 273184 77156 273186
rect 77064 273128 77114 273184
rect 77064 273126 77156 273128
rect 77109 273124 77156 273126
rect 77220 273124 77226 273188
rect 82997 273186 83044 273188
rect 82952 273184 83044 273186
rect 82952 273128 83002 273184
rect 82952 273126 83044 273128
rect 82997 273124 83044 273126
rect 83108 273124 83114 273188
rect 90725 273186 90772 273188
rect 90680 273184 90772 273186
rect 90680 273128 90730 273184
rect 90680 273126 90772 273128
rect 90725 273124 90772 273126
rect 90836 273124 90842 273188
rect 93669 273186 93716 273188
rect 93624 273184 93716 273186
rect 93624 273128 93674 273184
rect 93624 273126 93716 273128
rect 93669 273124 93716 273126
rect 93780 273124 93786 273188
rect 95877 273186 95924 273188
rect 95832 273184 95924 273186
rect 95832 273128 95882 273184
rect 95832 273126 95924 273128
rect 95877 273124 95924 273126
rect 95988 273124 95994 273188
rect 96061 273186 96127 273189
rect 101806 273186 101812 273188
rect 96061 273184 101812 273186
rect 96061 273128 96066 273184
rect 96122 273128 101812 273184
rect 96061 273126 101812 273128
rect 76005 273123 76071 273124
rect 77109 273123 77175 273124
rect 82997 273123 83063 273124
rect 90725 273123 90791 273124
rect 93669 273123 93735 273124
rect 95877 273123 95943 273124
rect 96061 273123 96127 273126
rect 101806 273124 101812 273126
rect 101876 273124 101882 273188
rect 199326 273124 199332 273188
rect 199396 273186 199402 273188
rect 318374 273186 318380 273188
rect 199396 273126 318380 273186
rect 199396 273124 199402 273126
rect 318374 273124 318380 273126
rect 318444 273124 318450 273188
rect 359406 273124 359412 273188
rect 359476 273186 359482 273188
rect 422661 273186 422727 273189
rect 422845 273188 422911 273189
rect 423397 273188 423463 273189
rect 425973 273188 426039 273189
rect 422845 273186 422892 273188
rect 359476 273184 422727 273186
rect 359476 273128 422666 273184
rect 422722 273128 422727 273184
rect 359476 273126 422727 273128
rect 422800 273184 422892 273186
rect 422800 273128 422850 273184
rect 422800 273126 422892 273128
rect 359476 273124 359482 273126
rect 422661 273123 422727 273126
rect 422845 273124 422892 273126
rect 422956 273124 422962 273188
rect 423397 273186 423444 273188
rect 423352 273184 423444 273186
rect 423352 273128 423402 273184
rect 423352 273126 423444 273128
rect 423397 273124 423444 273126
rect 423508 273124 423514 273188
rect 425973 273186 426020 273188
rect 425928 273184 426020 273186
rect 425928 273128 425978 273184
rect 425928 273126 426020 273128
rect 425973 273124 426020 273126
rect 426084 273124 426090 273188
rect 422845 273123 422911 273124
rect 423397 273123 423463 273124
rect 425973 273123 426039 273124
rect 61101 273050 61167 273053
rect 468477 273052 468543 273053
rect 470869 273052 470935 273053
rect 102726 273050 102732 273052
rect 61101 273048 102732 273050
rect 61101 272992 61106 273048
rect 61162 272992 102732 273048
rect 61101 272990 102732 272992
rect 61101 272987 61167 272990
rect 102726 272988 102732 272990
rect 102796 272988 102802 273052
rect 196750 272988 196756 273052
rect 196820 273050 196826 273052
rect 311014 273050 311020 273052
rect 196820 272990 311020 273050
rect 196820 272988 196826 272990
rect 311014 272988 311020 272990
rect 311084 272988 311090 273052
rect 377806 272988 377812 273052
rect 377876 273050 377882 273052
rect 425278 273050 425284 273052
rect 377876 272990 425284 273050
rect 377876 272988 377882 272990
rect 425278 272988 425284 272990
rect 425348 272988 425354 273052
rect 468477 273050 468524 273052
rect 468432 273048 468524 273050
rect 468432 272992 468482 273048
rect 468432 272990 468524 272992
rect 468477 272988 468524 272990
rect 468588 272988 468594 273052
rect 470869 273050 470916 273052
rect 470824 273048 470916 273050
rect 470824 272992 470874 273048
rect 470824 272990 470916 272992
rect 470869 272988 470916 272990
rect 470980 272988 470986 273052
rect 468477 272987 468543 272988
rect 470869 272987 470935 272988
rect 61469 272914 61535 272917
rect 285949 272916 286015 272917
rect 288157 272916 288223 272917
rect 290917 272916 290983 272917
rect 295885 272916 295951 272917
rect 303429 272916 303495 272917
rect 103830 272914 103836 272916
rect 61469 272912 103836 272914
rect 61469 272856 61474 272912
rect 61530 272856 103836 272912
rect 61469 272854 103836 272856
rect 61469 272851 61535 272854
rect 103830 272852 103836 272854
rect 103900 272852 103906 272916
rect 217358 272852 217364 272916
rect 217428 272914 217434 272916
rect 285949 272914 285996 272916
rect 217428 272854 277410 272914
rect 285904 272912 285996 272914
rect 285904 272856 285954 272912
rect 285904 272854 285996 272856
rect 217428 272852 217434 272854
rect 53833 272778 53899 272781
rect 54201 272778 54267 272781
rect 95877 272778 95943 272781
rect 96061 272780 96127 272781
rect 98453 272780 98519 272781
rect 96061 272778 96108 272780
rect 53833 272776 95943 272778
rect 53833 272720 53838 272776
rect 53894 272720 54206 272776
rect 54262 272720 95882 272776
rect 95938 272720 95943 272776
rect 53833 272718 95943 272720
rect 96016 272776 96108 272778
rect 96016 272720 96066 272776
rect 96016 272718 96108 272720
rect 53833 272715 53899 272718
rect 54201 272715 54267 272718
rect 95877 272715 95943 272718
rect 96061 272716 96108 272718
rect 96172 272716 96178 272780
rect 98453 272778 98500 272780
rect 98408 272776 98500 272778
rect 98408 272720 98458 272776
rect 98408 272718 98500 272720
rect 98453 272716 98500 272718
rect 98564 272716 98570 272780
rect 277350 272778 277410 272854
rect 285949 272852 285996 272854
rect 286060 272852 286066 272916
rect 288157 272914 288204 272916
rect 288112 272912 288204 272914
rect 288112 272856 288162 272912
rect 288112 272854 288204 272856
rect 288157 272852 288204 272854
rect 288268 272852 288274 272916
rect 290917 272914 290964 272916
rect 290872 272912 290964 272914
rect 290872 272856 290922 272912
rect 290872 272854 290964 272856
rect 290917 272852 290964 272854
rect 291028 272852 291034 272916
rect 295885 272914 295932 272916
rect 295840 272912 295932 272914
rect 295840 272856 295890 272912
rect 295840 272854 295932 272856
rect 295885 272852 295932 272854
rect 295996 272852 296002 272916
rect 303429 272914 303476 272916
rect 303384 272912 303476 272914
rect 303384 272856 303434 272912
rect 303384 272854 303476 272856
rect 303429 272852 303476 272854
rect 303540 272852 303546 272916
rect 422661 272914 422727 272917
rect 473445 272916 473511 272917
rect 475837 272916 475903 272917
rect 428222 272914 428228 272916
rect 422661 272912 428228 272914
rect 422661 272856 422666 272912
rect 422722 272856 428228 272912
rect 422661 272854 428228 272856
rect 285949 272851 286015 272852
rect 288157 272851 288223 272852
rect 290917 272851 290983 272852
rect 295885 272851 295951 272852
rect 303429 272851 303495 272852
rect 422661 272851 422727 272854
rect 428222 272852 428228 272854
rect 428292 272852 428298 272916
rect 473445 272914 473492 272916
rect 473400 272912 473492 272914
rect 473400 272856 473450 272912
rect 473400 272854 473492 272856
rect 473445 272852 473492 272854
rect 473556 272852 473562 272916
rect 475837 272914 475884 272916
rect 475792 272912 475884 272914
rect 475792 272856 475842 272912
rect 475792 272854 475884 272856
rect 475837 272852 475884 272854
rect 475948 272852 475954 272916
rect 473445 272851 473511 272852
rect 475837 272851 475903 272852
rect 298461 272780 298527 272781
rect 300853 272780 300919 272781
rect 478413 272780 478479 272781
rect 480805 272780 480871 272781
rect 293350 272778 293356 272780
rect 277350 272718 293356 272778
rect 293350 272716 293356 272718
rect 293420 272716 293426 272780
rect 298461 272778 298508 272780
rect 298416 272776 298508 272778
rect 298416 272720 298466 272776
rect 298416 272718 298508 272720
rect 298461 272716 298508 272718
rect 298572 272716 298578 272780
rect 300853 272778 300900 272780
rect 300808 272776 300900 272778
rect 300808 272720 300858 272776
rect 300808 272718 300900 272720
rect 300853 272716 300900 272718
rect 300964 272716 300970 272780
rect 478413 272778 478460 272780
rect 478368 272776 478460 272778
rect 478368 272720 478418 272776
rect 478368 272718 478460 272720
rect 478413 272716 478460 272718
rect 478524 272716 478530 272780
rect 480805 272778 480852 272780
rect 480760 272776 480852 272778
rect 480760 272720 480810 272776
rect 480760 272718 480852 272720
rect 480805 272716 480852 272718
rect 480916 272716 480922 272780
rect 96061 272715 96127 272716
rect 98453 272715 98519 272716
rect 298461 272715 298527 272716
rect 300853 272715 300919 272716
rect 478413 272715 478479 272716
rect 480805 272715 480871 272716
rect 59813 272642 59879 272645
rect 60917 272642 60983 272645
rect 305821 272644 305887 272645
rect 320909 272644 320975 272645
rect 116894 272642 116900 272644
rect 59813 272640 116900 272642
rect 59813 272584 59818 272640
rect 59874 272584 60922 272640
rect 60978 272584 116900 272640
rect 59813 272582 116900 272584
rect 59813 272579 59879 272582
rect 60917 272579 60983 272582
rect 116894 272580 116900 272582
rect 116964 272580 116970 272644
rect 305821 272642 305868 272644
rect 305776 272640 305868 272642
rect 305776 272584 305826 272640
rect 305776 272582 305868 272584
rect 305821 272580 305868 272582
rect 305932 272580 305938 272644
rect 320909 272642 320956 272644
rect 320864 272640 320956 272642
rect 320864 272584 320914 272640
rect 320864 272582 320956 272584
rect 320909 272580 320956 272582
rect 321020 272580 321026 272644
rect 377990 272580 377996 272644
rect 378060 272642 378066 272644
rect 380065 272642 380131 272645
rect 483197 272644 483263 272645
rect 485957 272644 486023 272645
rect 483197 272642 483244 272644
rect 378060 272640 380131 272642
rect 378060 272584 380070 272640
rect 380126 272584 380131 272640
rect 378060 272582 380131 272584
rect 483152 272640 483244 272642
rect 483152 272584 483202 272640
rect 483152 272582 483244 272584
rect 378060 272580 378066 272582
rect 305821 272579 305887 272580
rect 320909 272579 320975 272580
rect 380065 272579 380131 272582
rect 483197 272580 483244 272582
rect 483308 272580 483314 272644
rect 485957 272642 486004 272644
rect 485912 272640 486004 272642
rect 485912 272584 485962 272640
rect 485912 272582 486004 272584
rect 485957 272580 486004 272582
rect 486068 272580 486074 272644
rect 483197 272579 483263 272580
rect 485957 272579 486023 272580
rect 58525 272506 58591 272509
rect 60733 272506 60799 272509
rect 423765 272508 423831 272509
rect 117998 272506 118004 272508
rect 58525 272504 118004 272506
rect 58525 272448 58530 272504
rect 58586 272448 60738 272504
rect 60794 272448 118004 272504
rect 58525 272446 118004 272448
rect 58525 272443 58591 272446
rect 60733 272443 60799 272446
rect 117998 272444 118004 272446
rect 118068 272444 118074 272508
rect 423765 272506 423812 272508
rect 423720 272504 423812 272506
rect 423720 272448 423770 272504
rect 423720 272446 423812 272448
rect 423765 272444 423812 272446
rect 423876 272444 423882 272508
rect 423765 272443 423831 272444
rect 87597 272372 87663 272373
rect 94405 272372 94471 272373
rect 87597 272370 87644 272372
rect 87552 272368 87644 272370
rect 87552 272312 87602 272368
rect 87552 272310 87644 272312
rect 87597 272308 87644 272310
rect 87708 272308 87714 272372
rect 94405 272370 94452 272372
rect 94360 272368 94452 272370
rect 94360 272312 94410 272368
rect 94360 272310 94452 272312
rect 94405 272308 94452 272310
rect 94516 272308 94522 272372
rect 87597 272307 87663 272308
rect 94405 272307 94471 272308
rect 99373 272236 99439 272237
rect 265157 272236 265223 272237
rect 401685 272236 401751 272237
rect 415853 272236 415919 272237
rect 416037 272236 416103 272237
rect 455781 272236 455847 272237
rect 99373 272234 99420 272236
rect 99328 272232 99420 272234
rect 99328 272176 99378 272232
rect 99328 272174 99420 272176
rect 99373 272172 99420 272174
rect 99484 272172 99490 272236
rect 265157 272234 265204 272236
rect 265112 272232 265204 272234
rect 265112 272176 265162 272232
rect 265112 272174 265204 272176
rect 265157 272172 265204 272174
rect 265268 272172 265274 272236
rect 401685 272234 401732 272236
rect 401640 272232 401732 272234
rect 401640 272176 401690 272232
rect 401640 272174 401732 272176
rect 401685 272172 401732 272174
rect 401796 272172 401802 272236
rect 415853 272234 415900 272236
rect 415808 272232 415900 272234
rect 415808 272176 415858 272232
rect 415808 272174 415900 272176
rect 415853 272172 415900 272174
rect 415964 272172 415970 272236
rect 416037 272232 416084 272236
rect 416148 272234 416154 272236
rect 455781 272234 455828 272236
rect 416037 272176 416042 272232
rect 416037 272172 416084 272176
rect 416148 272174 416194 272234
rect 455736 272232 455828 272234
rect 455736 272176 455786 272232
rect 455736 272174 455828 272176
rect 416148 272172 416154 272174
rect 455781 272172 455828 272174
rect 455892 272172 455898 272236
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 99373 272171 99439 272172
rect 265157 272171 265223 272172
rect 401685 272171 401751 272172
rect 415853 272171 415919 272172
rect 416037 272171 416103 272172
rect 455781 272171 455847 272172
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 47669 271826 47735 271829
rect 48037 271826 48103 271829
rect 53281 271828 53347 271829
rect 53230 271826 53236 271828
rect 47669 271824 48103 271826
rect 47669 271768 47674 271824
rect 47730 271768 48042 271824
rect 48098 271768 48103 271824
rect 47669 271766 48103 271768
rect 53190 271766 53236 271826
rect 53300 271824 53347 271828
rect 53342 271768 53347 271824
rect 47669 271763 47735 271766
rect 48037 271763 48103 271766
rect 53230 271764 53236 271766
rect 53300 271764 53347 271768
rect 83958 271764 83964 271828
rect 84028 271826 84034 271828
rect 84193 271826 84259 271829
rect 84028 271824 84259 271826
rect 84028 271768 84198 271824
rect 84254 271768 84259 271824
rect 84028 271766 84259 271768
rect 84028 271764 84034 271766
rect 53281 271763 53347 271764
rect 84193 271763 84259 271766
rect 96613 271826 96679 271829
rect 100753 271828 100819 271829
rect 97022 271826 97028 271828
rect 96613 271824 97028 271826
rect 96613 271768 96618 271824
rect 96674 271768 97028 271824
rect 96613 271766 97028 271768
rect 96613 271763 96679 271766
rect 97022 271764 97028 271766
rect 97092 271764 97098 271828
rect 100702 271764 100708 271828
rect 100772 271826 100819 271828
rect 106273 271826 106339 271829
rect 106406 271826 106412 271828
rect 100772 271824 100864 271826
rect 100814 271768 100864 271824
rect 100772 271766 100864 271768
rect 106273 271824 106412 271826
rect 106273 271768 106278 271824
rect 106334 271768 106412 271824
rect 106273 271766 106412 271768
rect 100772 271764 100819 271766
rect 100753 271763 100819 271764
rect 106273 271763 106339 271766
rect 106406 271764 106412 271766
rect 106476 271764 106482 271828
rect 106549 271826 106615 271829
rect 112345 271828 112411 271829
rect 107510 271826 107516 271828
rect 106549 271824 107516 271826
rect 106549 271768 106554 271824
rect 106610 271768 107516 271824
rect 106549 271766 107516 271768
rect 106549 271763 106615 271766
rect 107510 271764 107516 271766
rect 107580 271764 107586 271828
rect 112294 271826 112300 271828
rect 112254 271766 112300 271826
rect 112364 271824 112411 271828
rect 112406 271768 112411 271824
rect 112294 271764 112300 271766
rect 112364 271764 112411 271768
rect 112345 271763 112411 271764
rect 123109 271826 123175 271829
rect 123518 271826 123524 271828
rect 123109 271824 123524 271826
rect 123109 271768 123114 271824
rect 123170 271768 123524 271824
rect 123109 271766 123524 271768
rect 123109 271763 123175 271766
rect 123518 271764 123524 271766
rect 123588 271764 123594 271828
rect 125593 271826 125659 271829
rect 125910 271826 125916 271828
rect 125593 271824 125916 271826
rect 125593 271768 125598 271824
rect 125654 271768 125916 271824
rect 125593 271766 125916 271768
rect 125593 271763 125659 271766
rect 125910 271764 125916 271766
rect 125980 271764 125986 271828
rect 128353 271826 128419 271829
rect 128670 271826 128676 271828
rect 128353 271824 128676 271826
rect 128353 271768 128358 271824
rect 128414 271768 128676 271824
rect 128353 271766 128676 271768
rect 128353 271763 128419 271766
rect 128670 271764 128676 271766
rect 128740 271764 128746 271828
rect 150934 271764 150940 271828
rect 151004 271826 151010 271828
rect 151353 271826 151419 271829
rect 151004 271824 151419 271826
rect 151004 271768 151358 271824
rect 151414 271768 151419 271824
rect 151004 271766 151419 271768
rect 151004 271764 151010 271766
rect 151353 271763 151419 271766
rect 154062 271764 154068 271828
rect 154132 271826 154138 271828
rect 154481 271826 154547 271829
rect 154132 271824 154547 271826
rect 154132 271768 154486 271824
rect 154542 271768 154547 271824
rect 154132 271766 154547 271768
rect 154132 271764 154138 271766
rect 154481 271763 154547 271766
rect 155902 271764 155908 271828
rect 155972 271826 155978 271828
rect 157241 271826 157307 271829
rect 155972 271824 157307 271826
rect 155972 271768 157246 271824
rect 157302 271768 157307 271824
rect 155972 271766 157307 271768
rect 155972 271764 155978 271766
rect 157241 271763 157307 271766
rect 215845 271826 215911 271829
rect 216213 271826 216279 271829
rect 263593 271828 263659 271829
rect 215845 271824 216279 271826
rect 215845 271768 215850 271824
rect 215906 271768 216218 271824
rect 216274 271768 216279 271824
rect 215845 271766 216279 271768
rect 215845 271763 215911 271766
rect 216213 271763 216279 271766
rect 263542 271764 263548 271828
rect 263612 271826 263659 271828
rect 264973 271826 265039 271829
rect 265934 271826 265940 271828
rect 263612 271824 263704 271826
rect 263654 271768 263704 271824
rect 263612 271766 263704 271768
rect 264973 271824 265940 271826
rect 264973 271768 264978 271824
rect 265034 271768 265940 271824
rect 264973 271766 265940 271768
rect 263612 271764 263659 271766
rect 263593 271763 263659 271764
rect 264973 271763 265039 271766
rect 265934 271764 265940 271766
rect 266004 271764 266010 271828
rect 268009 271826 268075 271829
rect 268326 271826 268332 271828
rect 268009 271824 268332 271826
rect 268009 271768 268014 271824
rect 268070 271768 268332 271824
rect 268009 271766 268332 271768
rect 268009 271763 268075 271766
rect 268326 271764 268332 271766
rect 268396 271764 268402 271828
rect 270493 271826 270559 271829
rect 270902 271826 270908 271828
rect 270493 271824 270908 271826
rect 270493 271768 270498 271824
rect 270554 271768 270908 271824
rect 270493 271766 270908 271768
rect 270493 271763 270559 271766
rect 270902 271764 270908 271766
rect 270972 271764 270978 271828
rect 271873 271826 271939 271829
rect 272558 271826 272564 271828
rect 271873 271824 272564 271826
rect 271873 271768 271878 271824
rect 271934 271768 272564 271824
rect 271873 271766 272564 271768
rect 271873 271763 271939 271766
rect 272558 271764 272564 271766
rect 272628 271764 272634 271828
rect 276013 271826 276079 271829
rect 276238 271826 276244 271828
rect 276013 271824 276244 271826
rect 276013 271768 276018 271824
rect 276074 271768 276244 271824
rect 276013 271766 276244 271768
rect 276013 271763 276079 271766
rect 276238 271764 276244 271766
rect 276308 271764 276314 271828
rect 277945 271826 278011 271829
rect 278446 271826 278452 271828
rect 277945 271824 278452 271826
rect 277945 271768 277950 271824
rect 278006 271768 278452 271824
rect 277945 271766 278452 271768
rect 277945 271763 278011 271766
rect 278446 271764 278452 271766
rect 278516 271764 278522 271828
rect 278998 271764 279004 271828
rect 279068 271826 279074 271828
rect 280061 271826 280127 271829
rect 279068 271824 280127 271826
rect 279068 271768 280066 271824
rect 280122 271768 280127 271824
rect 279068 271766 280127 271768
rect 279068 271764 279074 271766
rect 280061 271763 280127 271766
rect 280245 271826 280311 271829
rect 280838 271826 280844 271828
rect 280245 271824 280844 271826
rect 280245 271768 280250 271824
rect 280306 271768 280844 271824
rect 280245 271766 280844 271768
rect 280245 271763 280311 271766
rect 280838 271764 280844 271766
rect 280908 271764 280914 271828
rect 307753 271826 307819 271829
rect 308622 271826 308628 271828
rect 307753 271824 308628 271826
rect 307753 271768 307758 271824
rect 307814 271768 308628 271824
rect 307753 271766 308628 271768
rect 307753 271763 307819 271766
rect 308622 271764 308628 271766
rect 308692 271764 308698 271828
rect 313273 271826 313339 271829
rect 313406 271826 313412 271828
rect 313273 271824 313412 271826
rect 313273 271768 313278 271824
rect 313334 271768 313412 271824
rect 313273 271766 313412 271768
rect 313273 271763 313339 271766
rect 313406 271764 313412 271766
rect 313476 271764 313482 271828
rect 379145 271826 379211 271829
rect 427813 271826 427879 271829
rect 428590 271826 428596 271828
rect 379145 271824 383670 271826
rect 379145 271768 379150 271824
rect 379206 271768 383670 271824
rect 379145 271766 383670 271768
rect 379145 271763 379211 271766
rect 47761 271690 47827 271693
rect 84653 271692 84719 271693
rect 98085 271692 98151 271693
rect 79542 271690 79548 271692
rect 47761 271688 79548 271690
rect 47761 271632 47766 271688
rect 47822 271632 79548 271688
rect 47761 271630 79548 271632
rect 47761 271627 47827 271630
rect 79542 271628 79548 271630
rect 79612 271628 79618 271692
rect 84653 271690 84700 271692
rect 84608 271688 84700 271690
rect 84608 271632 84658 271688
rect 84608 271630 84700 271632
rect 84653 271628 84700 271630
rect 84764 271628 84770 271692
rect 98085 271688 98132 271692
rect 98196 271690 98202 271692
rect 107653 271690 107719 271693
rect 115933 271692 115999 271693
rect 108246 271690 108252 271692
rect 98085 271632 98090 271688
rect 98085 271628 98132 271632
rect 98196 271630 98242 271690
rect 107653 271688 108252 271690
rect 107653 271632 107658 271688
rect 107714 271632 108252 271688
rect 107653 271630 108252 271632
rect 98196 271628 98202 271630
rect 84653 271627 84719 271628
rect 98085 271627 98151 271628
rect 107653 271627 107719 271630
rect 108246 271628 108252 271630
rect 108316 271628 108322 271692
rect 115933 271690 115980 271692
rect 115888 271688 115980 271690
rect 115888 271632 115938 271688
rect 115888 271630 115980 271632
rect 115933 271628 115980 271630
rect 116044 271628 116050 271692
rect 117313 271690 117379 271693
rect 118366 271690 118372 271692
rect 117313 271688 118372 271690
rect 117313 271632 117318 271688
rect 117374 271632 118372 271688
rect 117313 271630 118372 271632
rect 115933 271627 115999 271628
rect 117313 271627 117379 271630
rect 118366 271628 118372 271630
rect 118436 271628 118442 271692
rect 120073 271690 120139 271693
rect 120758 271690 120764 271692
rect 120073 271688 120764 271690
rect 120073 271632 120078 271688
rect 120134 271632 120764 271688
rect 120073 271630 120764 271632
rect 120073 271627 120139 271630
rect 120758 271628 120764 271630
rect 120828 271628 120834 271692
rect 158478 271628 158484 271692
rect 158548 271690 158554 271692
rect 158621 271690 158687 271693
rect 158548 271688 158687 271690
rect 158548 271632 158626 271688
rect 158682 271632 158687 271688
rect 158548 271630 158687 271632
rect 158548 271628 158554 271630
rect 158621 271627 158687 271630
rect 160870 271628 160876 271692
rect 160940 271690 160946 271692
rect 161289 271690 161355 271693
rect 160940 271688 161355 271690
rect 160940 271632 161294 271688
rect 161350 271632 161355 271688
rect 160940 271630 161355 271632
rect 160940 271628 160946 271630
rect 161289 271627 161355 271630
rect 163446 271628 163452 271692
rect 163516 271690 163522 271692
rect 164141 271690 164207 271693
rect 163516 271688 164207 271690
rect 163516 271632 164146 271688
rect 164202 271632 164207 271688
rect 163516 271630 164207 271632
rect 163516 271628 163522 271630
rect 164141 271627 164207 271630
rect 166022 271628 166028 271692
rect 166092 271690 166098 271692
rect 198774 271690 198780 271692
rect 166092 271630 198780 271690
rect 166092 271628 166098 271630
rect 198774 271628 198780 271630
rect 198844 271628 198850 271692
rect 212073 271690 212139 271693
rect 315062 271690 315068 271692
rect 212073 271688 315068 271690
rect 212073 271632 212078 271688
rect 212134 271632 315068 271688
rect 212073 271630 315068 271632
rect 212073 271627 212139 271630
rect 315062 271628 315068 271630
rect 315132 271628 315138 271692
rect 383610 271690 383670 271766
rect 427813 271824 428596 271826
rect 427813 271768 427818 271824
rect 427874 271768 428596 271824
rect 427813 271766 428596 271768
rect 427813 271763 427879 271766
rect 428590 271764 428596 271766
rect 428660 271764 428666 271828
rect 433333 271826 433399 271829
rect 433558 271826 433564 271828
rect 433333 271824 433564 271826
rect 433333 271768 433338 271824
rect 433394 271768 433564 271824
rect 433333 271766 433564 271768
rect 433333 271763 433399 271766
rect 433558 271764 433564 271766
rect 433628 271764 433634 271828
rect 436093 271826 436159 271829
rect 436870 271826 436876 271828
rect 436093 271824 436876 271826
rect 436093 271768 436098 271824
rect 436154 271768 436876 271824
rect 436093 271766 436876 271768
rect 436093 271763 436159 271766
rect 436870 271764 436876 271766
rect 436940 271764 436946 271828
rect 437473 271826 437539 271829
rect 438526 271826 438532 271828
rect 437473 271824 438532 271826
rect 437473 271768 437478 271824
rect 437534 271768 438532 271824
rect 437473 271766 438532 271768
rect 437473 271763 437539 271766
rect 438526 271764 438532 271766
rect 438596 271764 438602 271828
rect 442993 271826 443059 271829
rect 443494 271826 443500 271828
rect 442993 271824 443500 271826
rect 442993 271768 442998 271824
rect 443054 271768 443500 271824
rect 442993 271766 443500 271768
rect 442993 271763 443059 271766
rect 443494 271764 443500 271766
rect 443564 271764 443570 271828
rect 445753 271826 445819 271829
rect 445886 271826 445892 271828
rect 445753 271824 445892 271826
rect 445753 271768 445758 271824
rect 445814 271768 445892 271824
rect 445753 271766 445892 271768
rect 445753 271763 445819 271766
rect 445886 271764 445892 271766
rect 445956 271764 445962 271828
rect 447133 271826 447199 271829
rect 448278 271826 448284 271828
rect 447133 271824 448284 271826
rect 447133 271768 447138 271824
rect 447194 271768 448284 271824
rect 447133 271766 448284 271768
rect 447133 271763 447199 271766
rect 448278 271764 448284 271766
rect 448348 271764 448354 271828
rect 449893 271826 449959 271829
rect 451038 271826 451044 271828
rect 449893 271824 451044 271826
rect 449893 271768 449898 271824
rect 449954 271768 451044 271824
rect 449893 271766 451044 271768
rect 449893 271763 449959 271766
rect 451038 271764 451044 271766
rect 451108 271764 451114 271828
rect 458173 271826 458239 271829
rect 458398 271826 458404 271828
rect 458173 271824 458404 271826
rect 458173 271768 458178 271824
rect 458234 271768 458404 271824
rect 458173 271766 458404 271768
rect 458173 271763 458239 271766
rect 458398 271764 458404 271766
rect 458468 271764 458474 271828
rect 465942 271690 465948 271692
rect 383610 271630 465948 271690
rect 465942 271628 465948 271630
rect 466012 271628 466018 271692
rect 503110 271628 503116 271692
rect 503180 271690 503186 271692
rect 503621 271690 503687 271693
rect 503180 271688 503687 271690
rect 503180 271632 503626 271688
rect 503682 271632 503687 271688
rect 503180 271630 503687 271632
rect 503180 271628 503186 271630
rect 503621 271627 503687 271630
rect 42241 271554 42307 271557
rect 61101 271554 61167 271557
rect 42241 271552 61167 271554
rect 42241 271496 42246 271552
rect 42302 271496 61106 271552
rect 61162 271496 61167 271552
rect 42241 271494 61167 271496
rect 42241 271491 42307 271494
rect 61101 271491 61167 271494
rect 100753 271554 100819 271557
rect 115841 271556 115907 271557
rect 101070 271554 101076 271556
rect 100753 271552 101076 271554
rect 100753 271496 100758 271552
rect 100814 271496 101076 271552
rect 100753 271494 101076 271496
rect 100753 271491 100819 271494
rect 101070 271492 101076 271494
rect 101140 271492 101146 271556
rect 115790 271554 115796 271556
rect 115750 271494 115796 271554
rect 115860 271552 115907 271556
rect 115902 271496 115907 271552
rect 115790 271492 115796 271494
rect 115860 271492 115907 271496
rect 115841 271491 115907 271492
rect 213177 271554 213243 271557
rect 213637 271554 213703 271557
rect 213177 271552 215402 271554
rect 213177 271496 213182 271552
rect 213238 271496 213642 271552
rect 213698 271496 215402 271552
rect 213177 271494 215402 271496
rect 213177 271491 213243 271494
rect 213637 271491 213703 271494
rect 47577 271418 47643 271421
rect 49141 271418 49207 271421
rect 104893 271418 104959 271421
rect 105854 271418 105860 271420
rect 47577 271416 55230 271418
rect 47577 271360 47582 271416
rect 47638 271360 49146 271416
rect 49202 271360 55230 271416
rect 47577 271358 55230 271360
rect 47577 271355 47643 271358
rect 49141 271355 49207 271358
rect 55170 271282 55230 271358
rect 104893 271416 105860 271418
rect 104893 271360 104898 271416
rect 104954 271360 105860 271416
rect 104893 271358 105860 271360
rect 104893 271355 104959 271358
rect 105854 271356 105860 271358
rect 105924 271356 105930 271420
rect 109217 271418 109283 271421
rect 109534 271418 109540 271420
rect 109217 271416 109540 271418
rect 109217 271360 109222 271416
rect 109278 271360 109540 271416
rect 109217 271358 109540 271360
rect 109217 271355 109283 271358
rect 109534 271356 109540 271358
rect 109604 271356 109610 271420
rect 113265 271418 113331 271421
rect 114318 271418 114324 271420
rect 113265 271416 114324 271418
rect 113265 271360 113270 271416
rect 113326 271360 114324 271416
rect 113265 271358 114324 271360
rect 113265 271355 113331 271358
rect 114318 271356 114324 271358
rect 114388 271356 114394 271420
rect 183134 271356 183140 271420
rect 183204 271418 183210 271420
rect 183461 271418 183527 271421
rect 183204 271416 183527 271418
rect 183204 271360 183466 271416
rect 183522 271360 183527 271416
rect 183204 271358 183527 271360
rect 215342 271418 215402 271494
rect 217174 271492 217180 271556
rect 217244 271554 217250 271556
rect 273478 271554 273484 271556
rect 217244 271494 273484 271554
rect 217244 271492 217250 271494
rect 273478 271492 273484 271494
rect 273548 271492 273554 271556
rect 276974 271492 276980 271556
rect 277044 271554 277050 271556
rect 277209 271554 277275 271557
rect 277044 271552 277275 271554
rect 277044 271496 277214 271552
rect 277270 271496 277275 271552
rect 277044 271494 277275 271496
rect 277044 271492 277050 271494
rect 277209 271491 277275 271494
rect 343398 271492 343404 271556
rect 343468 271554 343474 271556
rect 343541 271554 343607 271557
rect 343468 271552 343607 271554
rect 343468 271496 343546 271552
rect 343602 271496 343607 271552
rect 343468 271494 343607 271496
rect 343468 271492 343474 271494
rect 343541 271491 343607 271494
rect 376385 271554 376451 271557
rect 460974 271554 460980 271556
rect 376385 271552 460980 271554
rect 376385 271496 376390 271552
rect 376446 271496 460980 271552
rect 376385 271494 460980 271496
rect 376385 271491 376451 271494
rect 460974 271492 460980 271494
rect 461044 271492 461050 271556
rect 236494 271418 236500 271420
rect 215342 271358 236500 271418
rect 183204 271356 183210 271358
rect 183461 271355 183527 271358
rect 236494 271356 236500 271358
rect 236564 271356 236570 271420
rect 343214 271356 343220 271420
rect 343284 271418 343290 271420
rect 343449 271418 343515 271421
rect 343284 271416 343515 271418
rect 343284 271360 343454 271416
rect 343510 271360 343515 271416
rect 343284 271358 343515 271360
rect 343284 271356 343290 271358
rect 343449 271355 343515 271358
rect 377254 271356 377260 271420
rect 377324 271418 377330 271420
rect 408166 271418 408172 271420
rect 377324 271358 408172 271418
rect 377324 271356 377330 271358
rect 408166 271356 408172 271358
rect 408236 271356 408242 271420
rect 440233 271418 440299 271421
rect 440918 271418 440924 271420
rect 440233 271416 440924 271418
rect 440233 271360 440238 271416
rect 440294 271360 440924 271416
rect 440233 271358 440924 271360
rect 440233 271355 440299 271358
rect 440918 271356 440924 271358
rect 440988 271356 440994 271420
rect 88333 271284 88399 271285
rect 81934 271282 81940 271284
rect 55170 271222 81940 271282
rect 81934 271220 81940 271222
rect 82004 271220 82010 271284
rect 88333 271282 88380 271284
rect 88288 271280 88380 271282
rect 88288 271224 88338 271280
rect 88288 271222 88380 271224
rect 88333 271220 88380 271222
rect 88444 271220 88450 271284
rect 103513 271282 103579 271285
rect 103830 271282 103836 271284
rect 103513 271280 103836 271282
rect 103513 271224 103518 271280
rect 103574 271224 103836 271280
rect 103513 271222 103836 271224
rect 88333 271219 88399 271220
rect 103513 271219 103579 271222
rect 103830 271220 103836 271222
rect 103900 271220 103906 271284
rect 110413 271282 110479 271285
rect 113173 271284 113239 271285
rect 111006 271282 111012 271284
rect 110413 271280 111012 271282
rect 110413 271224 110418 271280
rect 110474 271224 111012 271280
rect 110413 271222 111012 271224
rect 110413 271219 110479 271222
rect 111006 271220 111012 271222
rect 111076 271220 111082 271284
rect 113173 271282 113220 271284
rect 113128 271280 113220 271282
rect 113128 271224 113178 271280
rect 113128 271222 113220 271224
rect 113173 271220 113220 271222
rect 113284 271220 113290 271284
rect 216213 271282 216279 271285
rect 237046 271282 237052 271284
rect 216213 271280 237052 271282
rect 216213 271224 216218 271280
rect 216274 271224 237052 271280
rect 216213 271222 237052 271224
rect 113173 271219 113239 271220
rect 216213 271219 216279 271222
rect 237046 271220 237052 271222
rect 237116 271220 237122 271284
rect 258257 271282 258323 271285
rect 258390 271282 258396 271284
rect 258257 271280 258396 271282
rect 258257 271224 258262 271280
rect 258318 271224 258396 271280
rect 258257 271222 258396 271224
rect 258257 271219 258323 271222
rect 258390 271220 258396 271222
rect 258460 271220 258466 271284
rect 260833 271282 260899 271285
rect 260966 271282 260972 271284
rect 260833 271280 260972 271282
rect 260833 271224 260838 271280
rect 260894 271224 260972 271280
rect 260833 271222 260972 271224
rect 260833 271219 260899 271222
rect 260966 271220 260972 271222
rect 261036 271220 261042 271284
rect 270493 271282 270559 271285
rect 271270 271282 271276 271284
rect 270493 271280 271276 271282
rect 270493 271224 270498 271280
rect 270554 271224 271276 271280
rect 270493 271222 271276 271224
rect 270493 271219 270559 271222
rect 271270 271220 271276 271222
rect 271340 271220 271346 271284
rect 376569 271282 376635 271285
rect 396022 271282 396028 271284
rect 376569 271280 396028 271282
rect 376569 271224 376574 271280
rect 376630 271224 396028 271280
rect 376569 271222 396028 271224
rect 376569 271219 376635 271222
rect 396022 271220 396028 271222
rect 396092 271220 396098 271284
rect 434713 271282 434779 271285
rect 503529 271284 503595 271285
rect 435950 271282 435956 271284
rect 434713 271280 435956 271282
rect 434713 271224 434718 271280
rect 434774 271224 435956 271280
rect 434713 271222 435956 271224
rect 434713 271219 434779 271222
rect 435950 271220 435956 271222
rect 436020 271220 436026 271284
rect 503478 271220 503484 271284
rect 503548 271282 503595 271284
rect 503548 271280 503640 271282
rect 503590 271224 503640 271280
rect 503548 271222 503640 271224
rect 503548 271220 503595 271222
rect 503529 271219 503595 271220
rect 48129 271146 48195 271149
rect 59813 271146 59879 271149
rect 48129 271144 59879 271146
rect 48129 271088 48134 271144
rect 48190 271088 59818 271144
rect 59874 271088 59879 271144
rect 48129 271086 59879 271088
rect 48129 271083 48195 271086
rect 59813 271083 59879 271086
rect 61561 271146 61627 271149
rect 62113 271146 62179 271149
rect 183461 271148 183527 271149
rect 119102 271146 119108 271148
rect 61561 271144 119108 271146
rect 61561 271088 61566 271144
rect 61622 271088 62118 271144
rect 62174 271088 119108 271144
rect 61561 271086 119108 271088
rect 61561 271083 61627 271086
rect 62113 271083 62179 271086
rect 119102 271084 119108 271086
rect 119172 271084 119178 271148
rect 183461 271146 183508 271148
rect 183416 271144 183508 271146
rect 183416 271088 183466 271144
rect 183416 271086 183508 271088
rect 183461 271084 183508 271086
rect 183572 271084 183578 271148
rect 247033 271146 247099 271149
rect 248270 271146 248276 271148
rect 247033 271144 248276 271146
rect 247033 271088 247038 271144
rect 247094 271088 248276 271144
rect 247033 271086 248276 271088
rect 183461 271083 183527 271084
rect 247033 271083 247099 271086
rect 248270 271084 248276 271086
rect 248340 271084 248346 271148
rect 252553 271146 252619 271149
rect 253606 271146 253612 271148
rect 252553 271144 253612 271146
rect 252553 271088 252558 271144
rect 252614 271088 253612 271144
rect 252553 271086 253612 271088
rect 252553 271083 252619 271086
rect 253606 271084 253612 271086
rect 253676 271084 253682 271148
rect 255313 271146 255379 271149
rect 256182 271146 256188 271148
rect 255313 271144 256188 271146
rect 255313 271088 255318 271144
rect 255374 271088 256188 271144
rect 255313 271086 256188 271088
rect 255313 271083 255379 271086
rect 256182 271084 256188 271086
rect 256252 271084 256258 271148
rect 379789 271146 379855 271149
rect 380157 271146 380223 271149
rect 397126 271146 397132 271148
rect 379789 271144 397132 271146
rect 379789 271088 379794 271144
rect 379850 271088 380162 271144
rect 380218 271088 397132 271144
rect 379789 271086 397132 271088
rect 379789 271083 379855 271086
rect 380157 271083 380223 271086
rect 397126 271084 397132 271086
rect 397196 271084 397202 271148
rect 409873 271146 409939 271149
rect 410742 271146 410748 271148
rect 409873 271144 410748 271146
rect 409873 271088 409878 271144
rect 409934 271088 410748 271144
rect 409873 271086 410748 271088
rect 409873 271083 409939 271086
rect 410742 271084 410748 271086
rect 410812 271084 410818 271148
rect 412725 271146 412791 271149
rect 413686 271146 413692 271148
rect 412725 271144 413692 271146
rect 412725 271088 412730 271144
rect 412786 271088 413692 271144
rect 412725 271086 413692 271088
rect 412725 271083 412791 271086
rect 413686 271084 413692 271086
rect 413756 271084 413762 271148
rect 418153 271146 418219 271149
rect 418470 271146 418476 271148
rect 418153 271144 418476 271146
rect 418153 271088 418158 271144
rect 418214 271088 418476 271144
rect 418153 271086 418476 271088
rect 418153 271083 418219 271086
rect 418470 271084 418476 271086
rect 418540 271084 418546 271148
rect 48037 271010 48103 271013
rect 77293 271010 77359 271013
rect 78254 271010 78260 271012
rect 48037 271008 64890 271010
rect 48037 270952 48042 271008
rect 48098 270952 64890 271008
rect 48037 270950 64890 270952
rect 48037 270947 48103 270950
rect 64830 270874 64890 270950
rect 77293 271008 78260 271010
rect 77293 270952 77298 271008
rect 77354 270952 78260 271008
rect 77293 270950 78260 270952
rect 77293 270947 77359 270950
rect 78254 270948 78260 270950
rect 78324 270948 78330 271012
rect 129733 271010 129799 271013
rect 130878 271010 130884 271012
rect 129733 271008 130884 271010
rect 129733 270952 129738 271008
rect 129794 270952 130884 271008
rect 129733 270950 130884 270952
rect 129733 270947 129799 270950
rect 130878 270948 130884 270950
rect 130948 270948 130954 271012
rect 210693 271010 210759 271013
rect 325550 271010 325556 271012
rect 210693 271008 325556 271010
rect 210693 270952 210698 271008
rect 210754 270952 325556 271008
rect 210693 270950 325556 270952
rect 210693 270947 210759 270950
rect 325550 270948 325556 270950
rect 325620 270948 325626 271012
rect 373533 271010 373599 271013
rect 462630 271010 462636 271012
rect 373533 271008 462636 271010
rect 373533 270952 373538 271008
rect 373594 270952 462636 271008
rect 373533 270950 462636 270952
rect 373533 270947 373599 270950
rect 462630 270948 462636 270950
rect 462700 270948 462706 271012
rect 80462 270874 80468 270876
rect 64830 270814 80468 270874
rect 80462 270812 80468 270814
rect 80532 270812 80538 270876
rect 88333 270874 88399 270877
rect 88742 270874 88748 270876
rect 88333 270872 88748 270874
rect 88333 270816 88338 270872
rect 88394 270816 88748 270872
rect 88333 270814 88748 270816
rect 88333 270811 88399 270814
rect 88742 270812 88748 270814
rect 88812 270812 88818 270876
rect 253933 270874 253999 270877
rect 254526 270874 254532 270876
rect 253933 270872 254532 270874
rect 253933 270816 253938 270872
rect 253994 270816 254532 270872
rect 253933 270814 254532 270816
rect 253933 270811 253999 270814
rect 254526 270812 254532 270814
rect 254596 270812 254602 270876
rect 267917 270874 267983 270877
rect 268694 270874 268700 270876
rect 267917 270872 268700 270874
rect 267917 270816 267922 270872
rect 267978 270816 268700 270872
rect 267917 270814 268700 270816
rect 267917 270811 267983 270814
rect 268694 270812 268700 270814
rect 268764 270812 268770 270876
rect 277393 270874 277459 270877
rect 278078 270874 278084 270876
rect 277393 270872 278084 270874
rect 277393 270816 277398 270872
rect 277454 270816 278084 270872
rect 277393 270814 278084 270816
rect 277393 270811 277459 270814
rect 278078 270812 278084 270814
rect 278148 270812 278154 270876
rect 405733 270874 405799 270877
rect 406510 270874 406516 270876
rect 405733 270872 406516 270874
rect 405733 270816 405738 270872
rect 405794 270816 406516 270872
rect 405733 270814 406516 270816
rect 405733 270811 405799 270814
rect 406510 270812 406516 270814
rect 406580 270812 406586 270876
rect 431953 270874 432019 270877
rect 432270 270874 432276 270876
rect 431953 270872 432276 270874
rect 431953 270816 431958 270872
rect 432014 270816 432276 270872
rect 431953 270814 432276 270816
rect 431953 270811 432019 270814
rect 432270 270812 432276 270814
rect 432340 270812 432346 270876
rect 433333 270874 433399 270877
rect 434662 270874 434668 270876
rect 433333 270872 434668 270874
rect 433333 270816 433338 270872
rect 433394 270816 434668 270872
rect 433333 270814 434668 270816
rect 433333 270811 433399 270814
rect 434662 270812 434668 270814
rect 434732 270812 434738 270876
rect 437473 270874 437539 270877
rect 438342 270874 438348 270876
rect 437473 270872 438348 270874
rect 437473 270816 437478 270872
rect 437534 270816 438348 270872
rect 437473 270814 438348 270816
rect 437473 270811 437539 270814
rect 438342 270812 438348 270814
rect 438412 270812 438418 270876
rect 438853 270874 438919 270877
rect 439078 270874 439084 270876
rect 438853 270872 439084 270874
rect 438853 270816 438858 270872
rect 438914 270816 439084 270872
rect 438853 270814 439084 270816
rect 438853 270811 438919 270814
rect 439078 270812 439084 270814
rect 439148 270812 439154 270876
rect 89713 270738 89779 270741
rect 90030 270738 90036 270740
rect 89713 270736 90036 270738
rect 89713 270680 89718 270736
rect 89774 270680 90036 270736
rect 89713 270678 90036 270680
rect 89713 270675 89779 270678
rect 90030 270676 90036 270678
rect 90100 270676 90106 270740
rect 92473 270738 92539 270741
rect 93342 270738 93348 270740
rect 92473 270736 93348 270738
rect 92473 270680 92478 270736
rect 92534 270680 93348 270736
rect 92473 270678 93348 270680
rect 92473 270675 92539 270678
rect 93342 270676 93348 270678
rect 93412 270676 93418 270740
rect 104893 270738 104959 270741
rect 105302 270738 105308 270740
rect 104893 270736 105308 270738
rect 104893 270680 104898 270736
rect 104954 270680 105308 270736
rect 104893 270678 105308 270680
rect 104893 270675 104959 270678
rect 105302 270676 105308 270678
rect 105372 270676 105378 270740
rect 147673 270738 147739 270741
rect 148542 270738 148548 270740
rect 147673 270736 148548 270738
rect 147673 270680 147678 270736
rect 147734 270680 148548 270736
rect 147673 270678 148548 270680
rect 147673 270675 147739 270678
rect 148542 270676 148548 270678
rect 148612 270676 148618 270740
rect 244222 270676 244228 270740
rect 244292 270738 244298 270740
rect 244365 270738 244431 270741
rect 244292 270736 244431 270738
rect 244292 270680 244370 270736
rect 244426 270680 244431 270736
rect 244292 270678 244431 270680
rect 244292 270676 244298 270678
rect 244365 270675 244431 270678
rect 251265 270738 251331 270741
rect 252318 270738 252324 270740
rect 251265 270736 252324 270738
rect 251265 270680 251270 270736
rect 251326 270680 252324 270736
rect 251265 270678 252324 270680
rect 251265 270675 251331 270678
rect 252318 270676 252324 270678
rect 252388 270676 252394 270740
rect 255313 270738 255379 270741
rect 255814 270738 255820 270740
rect 255313 270736 255820 270738
rect 255313 270680 255318 270736
rect 255374 270680 255820 270736
rect 255313 270678 255820 270680
rect 255313 270675 255379 270678
rect 255814 270676 255820 270678
rect 255884 270676 255890 270740
rect 259545 270738 259611 270741
rect 411345 270740 411411 270741
rect 260598 270738 260604 270740
rect 259545 270736 260604 270738
rect 259545 270680 259550 270736
rect 259606 270680 260604 270736
rect 259545 270678 260604 270680
rect 259545 270675 259611 270678
rect 260598 270676 260604 270678
rect 260668 270676 260674 270740
rect 411294 270676 411300 270740
rect 411364 270738 411411 270740
rect 429193 270738 429259 270741
rect 429694 270738 429700 270740
rect 411364 270736 411456 270738
rect 411406 270680 411456 270736
rect 411364 270678 411456 270680
rect 429193 270736 429700 270738
rect 429193 270680 429198 270736
rect 429254 270680 429700 270736
rect 429193 270678 429700 270680
rect 411364 270676 411411 270678
rect 411345 270675 411411 270676
rect 429193 270675 429259 270678
rect 429694 270676 429700 270678
rect 429764 270676 429770 270740
rect 59813 270602 59879 270605
rect 62205 270602 62271 270605
rect 59813 270600 62271 270602
rect 59813 270544 59818 270600
rect 59874 270544 62210 270600
rect 62266 270544 62271 270600
rect 59813 270542 62271 270544
rect 59813 270539 59879 270542
rect 62205 270539 62271 270542
rect 85573 270602 85639 270605
rect 86534 270602 86540 270604
rect 85573 270600 86540 270602
rect 85573 270544 85578 270600
rect 85634 270544 86540 270600
rect 85573 270542 86540 270544
rect 85573 270539 85639 270542
rect 86534 270540 86540 270542
rect 86604 270540 86610 270604
rect 91093 270602 91159 270605
rect 91318 270602 91324 270604
rect 91093 270600 91324 270602
rect 91093 270544 91098 270600
rect 91154 270544 91324 270600
rect 91093 270542 91324 270544
rect 91093 270539 91159 270542
rect 91318 270540 91324 270542
rect 91388 270540 91394 270604
rect 107653 270602 107719 270605
rect 108614 270602 108620 270604
rect 107653 270600 108620 270602
rect 107653 270544 107658 270600
rect 107714 270544 108620 270600
rect 107653 270542 108620 270544
rect 107653 270539 107719 270542
rect 108614 270540 108620 270542
rect 108684 270540 108690 270604
rect 110413 270602 110479 270605
rect 111190 270602 111196 270604
rect 110413 270600 111196 270602
rect 110413 270544 110418 270600
rect 110474 270544 111196 270600
rect 110413 270542 111196 270544
rect 110413 270539 110479 270542
rect 111190 270540 111196 270542
rect 111260 270540 111266 270604
rect 237373 270602 237439 270605
rect 242893 270604 242959 270605
rect 238150 270602 238156 270604
rect 237373 270600 238156 270602
rect 237373 270544 237378 270600
rect 237434 270544 238156 270600
rect 237373 270542 238156 270544
rect 237373 270539 237439 270542
rect 238150 270540 238156 270542
rect 238220 270540 238226 270604
rect 242893 270602 242940 270604
rect 242848 270600 242940 270602
rect 242848 270544 242898 270600
rect 242848 270542 242940 270544
rect 242893 270540 242940 270542
rect 243004 270540 243010 270604
rect 244273 270602 244339 270605
rect 245326 270602 245332 270604
rect 244273 270600 245332 270602
rect 244273 270544 244278 270600
rect 244334 270544 245332 270600
rect 244273 270542 245332 270544
rect 242893 270539 242959 270540
rect 244273 270539 244339 270542
rect 245326 270540 245332 270542
rect 245396 270540 245402 270604
rect 245653 270602 245719 270605
rect 246430 270602 246436 270604
rect 245653 270600 246436 270602
rect 245653 270544 245658 270600
rect 245714 270544 246436 270600
rect 245653 270542 246436 270544
rect 245653 270539 245719 270542
rect 246430 270540 246436 270542
rect 246500 270540 246506 270604
rect 247033 270602 247099 270605
rect 247718 270602 247724 270604
rect 247033 270600 247724 270602
rect 247033 270544 247038 270600
rect 247094 270544 247724 270600
rect 247033 270542 247724 270544
rect 247033 270539 247099 270542
rect 247718 270540 247724 270542
rect 247788 270540 247794 270604
rect 248505 270602 248571 270605
rect 248638 270602 248644 270604
rect 248505 270600 248644 270602
rect 248505 270544 248510 270600
rect 248566 270544 248644 270600
rect 248505 270542 248644 270544
rect 248505 270539 248571 270542
rect 248638 270540 248644 270542
rect 248708 270540 248714 270604
rect 249793 270602 249859 270605
rect 251173 270604 251239 270605
rect 250110 270602 250116 270604
rect 249793 270600 250116 270602
rect 249793 270544 249798 270600
rect 249854 270544 250116 270600
rect 249793 270542 250116 270544
rect 249793 270539 249859 270542
rect 250110 270540 250116 270542
rect 250180 270540 250186 270604
rect 251173 270602 251220 270604
rect 251128 270600 251220 270602
rect 251128 270544 251178 270600
rect 251128 270542 251220 270544
rect 251173 270540 251220 270542
rect 251284 270540 251290 270604
rect 252553 270602 252619 270605
rect 253422 270602 253428 270604
rect 252553 270600 253428 270602
rect 252553 270544 252558 270600
rect 252614 270544 253428 270600
rect 252553 270542 253428 270544
rect 251173 270539 251239 270540
rect 252553 270539 252619 270542
rect 253422 270540 253428 270542
rect 253492 270540 253498 270604
rect 256693 270602 256759 270605
rect 256918 270602 256924 270604
rect 256693 270600 256924 270602
rect 256693 270544 256698 270600
rect 256754 270544 256924 270600
rect 256693 270542 256924 270544
rect 256693 270539 256759 270542
rect 256918 270540 256924 270542
rect 256988 270540 256994 270604
rect 258073 270602 258139 270605
rect 259453 270604 259519 270605
rect 258390 270602 258396 270604
rect 258073 270600 258396 270602
rect 258073 270544 258078 270600
rect 258134 270544 258396 270600
rect 258073 270542 258396 270544
rect 258073 270539 258139 270542
rect 258390 270540 258396 270542
rect 258460 270540 258466 270604
rect 259453 270602 259500 270604
rect 259408 270600 259500 270602
rect 259408 270544 259458 270600
rect 259408 270542 259500 270544
rect 259453 270540 259500 270542
rect 259564 270540 259570 270604
rect 260833 270602 260899 270605
rect 262070 270602 262076 270604
rect 260833 270600 262076 270602
rect 260833 270544 260838 270600
rect 260894 270544 262076 270600
rect 260833 270542 262076 270544
rect 259453 270539 259519 270540
rect 260833 270539 260899 270542
rect 262070 270540 262076 270542
rect 262140 270540 262146 270604
rect 262213 270602 262279 270605
rect 262806 270602 262812 270604
rect 262213 270600 262812 270602
rect 262213 270544 262218 270600
rect 262274 270544 262812 270600
rect 262213 270542 262812 270544
rect 262213 270539 262279 270542
rect 262806 270540 262812 270542
rect 262876 270540 262882 270604
rect 263593 270602 263659 270605
rect 263910 270602 263916 270604
rect 263593 270600 263916 270602
rect 263593 270544 263598 270600
rect 263654 270544 263916 270600
rect 263593 270542 263916 270544
rect 263593 270539 263659 270542
rect 263910 270540 263916 270542
rect 263980 270540 263986 270604
rect 266353 270602 266419 270605
rect 267590 270602 267596 270604
rect 266353 270600 267596 270602
rect 266353 270544 266358 270600
rect 266414 270544 267596 270600
rect 266353 270542 267596 270544
rect 266353 270539 266419 270542
rect 267590 270540 267596 270542
rect 267660 270540 267666 270604
rect 269113 270602 269179 270605
rect 269798 270602 269804 270604
rect 269113 270600 269804 270602
rect 269113 270544 269118 270600
rect 269174 270544 269804 270600
rect 269113 270542 269804 270544
rect 269113 270539 269179 270542
rect 269798 270540 269804 270542
rect 269868 270540 269874 270604
rect 273161 270602 273227 270605
rect 274398 270602 274404 270604
rect 273161 270600 274404 270602
rect 273161 270544 273166 270600
rect 273222 270544 274404 270600
rect 273161 270542 274404 270544
rect 273161 270539 273227 270542
rect 274398 270540 274404 270542
rect 274468 270540 274474 270604
rect 274633 270602 274699 270605
rect 275318 270602 275324 270604
rect 274633 270600 275324 270602
rect 274633 270544 274638 270600
rect 274694 270544 275324 270600
rect 274633 270542 275324 270544
rect 274633 270539 274699 270542
rect 275318 270540 275324 270542
rect 275388 270540 275394 270604
rect 375741 270602 375807 270605
rect 376569 270602 376635 270605
rect 397453 270604 397519 270605
rect 397453 270602 397500 270604
rect 375741 270600 376635 270602
rect 375741 270544 375746 270600
rect 375802 270544 376574 270600
rect 376630 270544 376635 270600
rect 375741 270542 376635 270544
rect 397408 270600 397500 270602
rect 397408 270544 397458 270600
rect 397408 270542 397500 270544
rect 375741 270539 375807 270542
rect 376569 270539 376635 270542
rect 397453 270540 397500 270542
rect 397564 270540 397570 270604
rect 398833 270602 398899 270605
rect 399518 270602 399524 270604
rect 398833 270600 399524 270602
rect 398833 270544 398838 270600
rect 398894 270544 399524 270600
rect 398833 270542 399524 270544
rect 397453 270539 397519 270540
rect 398833 270539 398899 270542
rect 399518 270540 399524 270542
rect 399588 270540 399594 270604
rect 400213 270602 400279 270605
rect 402973 270604 403039 270605
rect 400438 270602 400444 270604
rect 400213 270600 400444 270602
rect 400213 270544 400218 270600
rect 400274 270544 400444 270600
rect 400213 270542 400444 270544
rect 400213 270539 400279 270542
rect 400438 270540 400444 270542
rect 400508 270540 400514 270604
rect 402973 270600 403020 270604
rect 403084 270602 403090 270604
rect 403341 270602 403407 270605
rect 404118 270602 404124 270604
rect 402973 270544 402978 270600
rect 402973 270540 403020 270544
rect 403084 270542 403130 270602
rect 403341 270600 404124 270602
rect 403341 270544 403346 270600
rect 403402 270544 404124 270600
rect 403341 270542 404124 270544
rect 403084 270540 403090 270542
rect 402973 270539 403039 270540
rect 403341 270539 403407 270542
rect 404118 270540 404124 270542
rect 404188 270540 404194 270604
rect 404353 270602 404419 270605
rect 405038 270602 405044 270604
rect 404353 270600 405044 270602
rect 404353 270544 404358 270600
rect 404414 270544 405044 270600
rect 404353 270542 405044 270544
rect 404353 270539 404419 270542
rect 405038 270540 405044 270542
rect 405108 270540 405114 270604
rect 407113 270602 407179 270605
rect 407614 270602 407620 270604
rect 407113 270600 407620 270602
rect 407113 270544 407118 270600
rect 407174 270544 407620 270600
rect 407113 270542 407620 270544
rect 407113 270539 407179 270542
rect 407614 270540 407620 270542
rect 407684 270540 407690 270604
rect 408493 270602 408559 270605
rect 408718 270602 408724 270604
rect 408493 270600 408724 270602
rect 408493 270544 408498 270600
rect 408554 270544 408724 270600
rect 408493 270542 408724 270544
rect 408493 270539 408559 270542
rect 408718 270540 408724 270542
rect 408788 270540 408794 270604
rect 409873 270602 409939 270605
rect 410006 270602 410012 270604
rect 409873 270600 410012 270602
rect 409873 270544 409878 270600
rect 409934 270544 410012 270600
rect 409873 270542 410012 270544
rect 409873 270539 409939 270542
rect 410006 270540 410012 270542
rect 410076 270540 410082 270604
rect 411253 270602 411319 270605
rect 412398 270602 412404 270604
rect 411253 270600 412404 270602
rect 411253 270544 411258 270600
rect 411314 270544 412404 270600
rect 411253 270542 412404 270544
rect 411253 270539 411319 270542
rect 412398 270540 412404 270542
rect 412468 270540 412474 270604
rect 413001 270602 413067 270605
rect 413318 270602 413324 270604
rect 413001 270600 413324 270602
rect 413001 270544 413006 270600
rect 413062 270544 413324 270600
rect 413001 270542 413324 270544
rect 413001 270539 413067 270542
rect 413318 270540 413324 270542
rect 413388 270540 413394 270604
rect 414013 270602 414079 270605
rect 414422 270602 414428 270604
rect 414013 270600 414428 270602
rect 414013 270544 414018 270600
rect 414074 270544 414428 270600
rect 414013 270542 414428 270544
rect 414013 270539 414079 270542
rect 414422 270540 414428 270542
rect 414492 270540 414498 270604
rect 416773 270602 416839 270605
rect 418153 270604 418219 270605
rect 416998 270602 417004 270604
rect 416773 270600 417004 270602
rect 416773 270544 416778 270600
rect 416834 270544 417004 270600
rect 416773 270542 417004 270544
rect 416773 270539 416839 270542
rect 416998 270540 417004 270542
rect 417068 270540 417074 270604
rect 418102 270540 418108 270604
rect 418172 270602 418219 270604
rect 419533 270602 419599 270605
rect 420678 270602 420684 270604
rect 418172 270600 418264 270602
rect 418214 270544 418264 270600
rect 418172 270542 418264 270544
rect 419533 270600 420684 270602
rect 419533 270544 419538 270600
rect 419594 270544 420684 270600
rect 419533 270542 420684 270544
rect 418172 270540 418219 270542
rect 418153 270539 418219 270540
rect 419533 270539 419599 270542
rect 420678 270540 420684 270542
rect 420748 270540 420754 270604
rect 420913 270602 420979 270605
rect 421782 270602 421788 270604
rect 420913 270600 421788 270602
rect 420913 270544 420918 270600
rect 420974 270544 421788 270600
rect 420913 270542 421788 270544
rect 420913 270539 420979 270542
rect 421782 270540 421788 270542
rect 421852 270540 421858 270604
rect 91502 270466 91508 270468
rect 64830 270406 91508 270466
rect 51809 270330 51875 270333
rect 57646 270330 57652 270332
rect 51809 270328 57652 270330
rect 51809 270272 51814 270328
rect 51870 270272 57652 270328
rect 51809 270270 57652 270272
rect 51809 270267 51875 270270
rect 57646 270268 57652 270270
rect 57716 270330 57722 270332
rect 64830 270330 64890 270406
rect 91502 270404 91508 270406
rect 91572 270404 91578 270468
rect 206185 270466 206251 270469
rect 206737 270466 206803 270469
rect 209405 270466 209471 270469
rect 323342 270466 323348 270468
rect 206185 270464 207674 270466
rect 206185 270408 206190 270464
rect 206246 270408 206742 270464
rect 206798 270408 207674 270464
rect 206185 270406 207674 270408
rect 206185 270403 206251 270406
rect 206737 270403 206803 270406
rect 57716 270270 64890 270330
rect 207614 270330 207674 270406
rect 209405 270464 323348 270466
rect 209405 270408 209410 270464
rect 209466 270408 323348 270464
rect 209405 270406 323348 270408
rect 209405 270403 209471 270406
rect 323342 270404 323348 270406
rect 323412 270404 323418 270468
rect 379421 270466 379487 270469
rect 379789 270466 379855 270469
rect 435766 270466 435772 270468
rect 379421 270464 379855 270466
rect 379421 270408 379426 270464
rect 379482 270408 379794 270464
rect 379850 270408 379855 270464
rect 379421 270406 379855 270408
rect 379421 270403 379487 270406
rect 379789 270403 379855 270406
rect 383610 270406 435772 270466
rect 239254 270330 239260 270332
rect 207614 270270 239260 270330
rect 57716 270268 57722 270270
rect 239254 270268 239260 270270
rect 239324 270268 239330 270332
rect 376477 270330 376543 270333
rect 383610 270330 383670 270406
rect 435766 270404 435772 270406
rect 435836 270404 435842 270468
rect 376477 270328 383670 270330
rect 376477 270272 376482 270328
rect 376538 270272 383670 270328
rect 376477 270270 383670 270272
rect 376477 270267 376543 270270
rect 217542 269996 217548 270060
rect 217612 270058 217618 270060
rect 219617 270058 219683 270061
rect 220721 270058 220787 270061
rect 217612 270056 220787 270058
rect 217612 270000 219622 270056
rect 219678 270000 220726 270056
rect 220782 270000 220787 270056
rect 217612 269998 220787 270000
rect 217612 269996 217618 269998
rect 219617 269995 219683 269998
rect 220721 269995 220787 269998
rect 372521 270058 372587 270061
rect 376385 270058 376451 270061
rect 372521 270056 379530 270058
rect 372521 270000 372526 270056
rect 372582 270000 376390 270056
rect 376446 270000 379530 270056
rect 372521 269998 379530 270000
rect 372521 269995 372587 269998
rect 376385 269995 376451 269998
rect 209497 269922 209563 269925
rect 213545 269922 213611 269925
rect 241646 269922 241652 269924
rect 209497 269920 241652 269922
rect 209497 269864 209502 269920
rect 209558 269864 213550 269920
rect 213606 269864 241652 269920
rect 209497 269862 241652 269864
rect 209497 269859 209563 269862
rect 213545 269859 213611 269862
rect 241646 269860 241652 269862
rect 241716 269860 241722 269924
rect 374913 269922 374979 269925
rect 376477 269922 376543 269925
rect 374913 269920 376543 269922
rect 374913 269864 374918 269920
rect 374974 269864 376482 269920
rect 376538 269864 376543 269920
rect 374913 269862 376543 269864
rect 379470 269922 379530 269998
rect 419206 269922 419212 269924
rect 379470 269862 419212 269922
rect 374913 269859 374979 269862
rect 376477 269859 376543 269862
rect 419206 269860 419212 269862
rect 419276 269860 419282 269924
rect 208117 269786 208183 269789
rect 210969 269786 211035 269789
rect 240542 269786 240548 269788
rect 208117 269784 240548 269786
rect 208117 269728 208122 269784
rect 208178 269728 210974 269784
rect 211030 269728 240548 269784
rect 208117 269726 240548 269728
rect 208117 269723 208183 269726
rect 210969 269723 211035 269726
rect 240542 269724 240548 269726
rect 240612 269724 240618 269788
rect 379789 269786 379855 269789
rect 427670 269786 427676 269788
rect 379789 269784 427676 269786
rect 379789 269728 379794 269784
rect 379850 269728 427676 269784
rect 379789 269726 427676 269728
rect 379789 269723 379855 269726
rect 427670 269724 427676 269726
rect 427740 269724 427746 269788
rect 375833 269378 375899 269381
rect 376753 269378 376819 269381
rect 387885 269378 387951 269381
rect 375833 269376 387951 269378
rect 375833 269320 375838 269376
rect 375894 269320 376758 269376
rect 376814 269320 387890 269376
rect 387946 269320 387951 269376
rect 375833 269318 387951 269320
rect 375833 269315 375899 269318
rect 376753 269315 376819 269318
rect 387885 269315 387951 269318
rect 372981 269242 373047 269245
rect 378685 269242 378751 269245
rect 390553 269242 390619 269245
rect 372981 269240 390619 269242
rect 372981 269184 372986 269240
rect 373042 269184 378690 269240
rect 378746 269184 390558 269240
rect 390614 269184 390619 269240
rect 372981 269182 390619 269184
rect 372981 269179 373047 269182
rect 378685 269179 378751 269182
rect 390553 269179 390619 269182
rect 44950 268500 44956 268564
rect 45020 268562 45026 268564
rect 46381 268562 46447 268565
rect 77385 268562 77451 268565
rect 45020 268560 77451 268562
rect 45020 268504 46386 268560
rect 46442 268504 77390 268560
rect 77446 268504 77451 268560
rect 45020 268502 77451 268504
rect 45020 268500 45026 268502
rect 46381 268499 46447 268502
rect 77385 268499 77451 268502
rect 44766 268364 44772 268428
rect 44836 268426 44842 268428
rect 46473 268426 46539 268429
rect 85757 268426 85823 268429
rect 44836 268424 85823 268426
rect 44836 268368 46478 268424
rect 46534 268368 85762 268424
rect 85818 268368 85823 268424
rect 44836 268366 85823 268368
rect 44836 268364 44842 268366
rect 46473 268363 46539 268366
rect 85757 268363 85823 268366
rect 376886 267548 376892 267612
rect 376956 267610 376962 267612
rect 377438 267610 377444 267612
rect 376956 267550 377444 267610
rect 376956 267548 376962 267550
rect 377438 267548 377444 267550
rect 377508 267610 377514 267612
rect 377673 267610 377739 267613
rect 377508 267608 377739 267610
rect 377508 267552 377678 267608
rect 377734 267552 377739 267608
rect 377508 267550 377739 267552
rect 377508 267548 377514 267550
rect 377673 267547 377739 267550
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 54334 254010 54340 254012
rect 6870 253950 54340 254010
rect 54334 253948 54340 253950
rect 54404 253948 54410 254012
rect 190862 253676 190868 253740
rect 190932 253738 190938 253740
rect 191741 253738 191807 253741
rect 190932 253736 191807 253738
rect 190932 253680 191746 253736
rect 191802 253680 191807 253736
rect 190932 253678 191807 253680
rect 190932 253676 190938 253678
rect 191741 253675 191807 253678
rect 338430 253540 338436 253604
rect 338500 253602 338506 253604
rect 339401 253602 339467 253605
rect 338500 253600 339467 253602
rect 338500 253544 339406 253600
rect 339462 253544 339467 253600
rect 338500 253542 339467 253544
rect 338500 253540 338506 253542
rect 339401 253539 339467 253542
rect 499798 253268 499804 253332
rect 499868 253330 499874 253332
rect 500861 253330 500927 253333
rect 499868 253328 500927 253330
rect 499868 253272 500866 253328
rect 500922 253272 500927 253328
rect 499868 253270 500927 253272
rect 499868 253268 499874 253270
rect 500861 253267 500927 253270
rect 178534 253132 178540 253196
rect 178604 253194 178610 253196
rect 179321 253194 179387 253197
rect 178604 253192 179387 253194
rect 178604 253136 179326 253192
rect 179382 253136 179387 253192
rect 178604 253134 179387 253136
rect 178604 253132 178610 253134
rect 179321 253131 179387 253134
rect 179638 253132 179644 253196
rect 179708 253194 179714 253196
rect 180517 253194 180583 253197
rect 179708 253192 180583 253194
rect 179708 253136 180522 253192
rect 180578 253136 180583 253192
rect 179708 253134 180583 253136
rect 179708 253132 179714 253134
rect 180517 253131 180583 253134
rect 350942 253132 350948 253196
rect 351012 253194 351018 253196
rect 351821 253194 351887 253197
rect 351012 253192 351887 253194
rect 351012 253136 351826 253192
rect 351882 253136 351887 253192
rect 351012 253134 351887 253136
rect 351012 253132 351018 253134
rect 351821 253131 351887 253134
rect 339718 252996 339724 253060
rect 339788 253058 339794 253060
rect 340781 253058 340847 253061
rect 339788 253056 340847 253058
rect 339788 253000 340786 253056
rect 340842 253000 340847 253056
rect 339788 252998 340847 253000
rect 339788 252996 339794 252998
rect 340781 252995 340847 252998
rect 498510 252724 498516 252788
rect 498580 252786 498586 252788
rect 499205 252786 499271 252789
rect 498580 252784 499271 252786
rect 498580 252728 499210 252784
rect 499266 252728 499271 252784
rect 498580 252726 499271 252728
rect 498580 252724 498586 252726
rect 499205 252723 499271 252726
rect 510889 252652 510955 252653
rect 510838 252650 510844 252652
rect 510798 252590 510844 252650
rect 510908 252648 510955 252652
rect 510950 252592 510955 252648
rect 510838 252588 510844 252590
rect 510908 252588 510955 252592
rect 510889 252587 510955 252588
rect 57646 252452 57652 252516
rect 57716 252514 57722 252516
rect 60733 252514 60799 252517
rect 57716 252512 60799 252514
rect 57716 252456 60738 252512
rect 60794 252456 60799 252512
rect 57716 252454 60799 252456
rect 57716 252452 57722 252454
rect 60733 252451 60799 252454
rect 216990 252452 216996 252516
rect 217060 252514 217066 252516
rect 217961 252514 218027 252517
rect 217060 252512 218027 252514
rect 217060 252456 217966 252512
rect 218022 252456 218027 252512
rect 217060 252454 218027 252456
rect 217060 252452 217066 252454
rect 217961 252451 218027 252454
rect 377673 252514 377739 252517
rect 377990 252514 377996 252516
rect 377673 252512 377996 252514
rect 377673 252456 377678 252512
rect 377734 252456 377996 252512
rect 377673 252454 377996 252456
rect 377673 252451 377739 252454
rect 377990 252452 377996 252454
rect 378060 252452 378066 252516
rect 198825 246258 198891 246261
rect 358905 246258 358971 246261
rect 519261 246258 519327 246261
rect 196558 246256 198891 246258
rect 196558 246200 198830 246256
rect 198886 246200 198891 246256
rect 196558 246198 198891 246200
rect 196558 246190 196618 246198
rect 198825 246195 198891 246198
rect 356562 246256 358971 246258
rect 356562 246200 358910 246256
rect 358966 246200 358971 246256
rect 356562 246198 358971 246200
rect 356562 246190 356622 246198
rect 358905 246195 358971 246198
rect 516558 246256 519327 246258
rect 516558 246200 519266 246256
rect 519322 246200 519327 246256
rect 516558 246198 519327 246200
rect 516558 246190 516618 246198
rect 519261 246195 519327 246198
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 57237 204234 57303 204237
rect 57605 204234 57671 204237
rect 57237 204232 60062 204234
rect 57237 204176 57242 204232
rect 57298 204176 57610 204232
rect 57666 204176 60062 204232
rect 57237 204174 60062 204176
rect 57237 204171 57303 204174
rect 57605 204171 57671 204174
rect 60002 203894 60062 204174
rect 217409 203962 217475 203965
rect 217869 203962 217935 203965
rect 377213 203962 377279 203965
rect 377397 203962 377463 203965
rect 217409 203960 219450 203962
rect 217409 203904 217414 203960
rect 217470 203904 217874 203960
rect 217930 203924 219450 203960
rect 377213 203960 379530 203962
rect 217930 203904 220064 203924
rect 217409 203902 220064 203904
rect 217409 203899 217475 203902
rect 217869 203899 217935 203902
rect 219390 203864 220064 203902
rect 377213 203904 377218 203960
rect 377274 203904 377402 203960
rect 377458 203924 379530 203960
rect 377458 203904 380052 203924
rect 377213 203902 380052 203904
rect 377213 203899 377279 203902
rect 377397 203899 377463 203902
rect 379470 203864 380052 203902
rect 56869 203418 56935 203421
rect 57513 203418 57579 203421
rect 56869 203416 60062 203418
rect 56869 203360 56874 203416
rect 56930 203360 57518 203416
rect 57574 203360 60062 203416
rect 56869 203358 60062 203360
rect 56869 203355 56935 203358
rect 57513 203355 57579 203358
rect 60002 202942 60062 203358
rect 216857 203010 216923 203013
rect 217869 203010 217935 203013
rect 377029 203010 377095 203013
rect 216857 203008 219450 203010
rect 216857 202952 216862 203008
rect 216918 202952 217874 203008
rect 217930 202972 219450 203008
rect 377029 203008 379530 203010
rect 217930 202952 220064 202972
rect 216857 202950 220064 202952
rect 216857 202947 216923 202950
rect 217869 202947 217935 202950
rect 219390 202912 220064 202950
rect 377029 202952 377034 203008
rect 377090 202972 379530 203008
rect 377090 202952 380052 202972
rect 377029 202950 380052 202952
rect 377029 202947 377095 202950
rect 379470 202912 380052 202950
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 376845 201378 376911 201381
rect 377581 201378 377647 201381
rect 376845 201376 377647 201378
rect 376845 201320 376850 201376
rect 376906 201320 377586 201376
rect 377642 201320 377647 201376
rect 376845 201318 377647 201320
rect 376845 201315 376911 201318
rect 377581 201315 377647 201318
rect 57605 200834 57671 200837
rect 217593 200834 217659 200837
rect 377581 200834 377647 200837
rect 57605 200832 60062 200834
rect 57605 200776 57610 200832
rect 57666 200776 60062 200832
rect 57605 200774 60062 200776
rect 57605 200771 57671 200774
rect 60002 200766 60062 200774
rect 217593 200832 219450 200834
rect 217593 200776 217598 200832
rect 217654 200796 219450 200832
rect 377581 200832 379530 200834
rect 217654 200776 220064 200796
rect 217593 200774 220064 200776
rect 217593 200771 217659 200774
rect 219390 200736 220064 200774
rect 377581 200776 377586 200832
rect 377642 200796 379530 200832
rect 377642 200776 380052 200796
rect 377581 200774 380052 200776
rect 377581 200771 377647 200774
rect 379470 200736 380052 200774
rect 57697 199882 57763 199885
rect 217685 199882 217751 199885
rect 376937 199882 377003 199885
rect 57697 199880 60062 199882
rect 57697 199824 57702 199880
rect 57758 199824 60062 199880
rect 57697 199822 60062 199824
rect 57697 199819 57763 199822
rect 60002 199814 60062 199822
rect 217685 199880 219450 199882
rect 217685 199824 217690 199880
rect 217746 199844 219450 199880
rect 376937 199880 379530 199882
rect 217746 199824 220064 199844
rect 217685 199822 220064 199824
rect 217685 199819 217751 199822
rect 219390 199784 220064 199822
rect 376937 199824 376942 199880
rect 376998 199844 379530 199880
rect 376998 199824 380052 199844
rect 376937 199822 380052 199824
rect 376937 199819 377003 199822
rect 379470 199784 380052 199822
rect 57421 198794 57487 198797
rect 57697 198794 57763 198797
rect 57421 198792 57763 198794
rect 57421 198736 57426 198792
rect 57482 198736 57702 198792
rect 57758 198736 57763 198792
rect 57421 198734 57763 198736
rect 57421 198731 57487 198734
rect 57697 198731 57763 198734
rect 216857 198794 216923 198797
rect 217685 198794 217751 198797
rect 216857 198792 217751 198794
rect 216857 198736 216862 198792
rect 216918 198736 217690 198792
rect 217746 198736 217751 198792
rect 216857 198734 217751 198736
rect 216857 198731 216923 198734
rect 217685 198731 217751 198734
rect 57697 198114 57763 198117
rect 217777 198114 217843 198117
rect 377673 198114 377739 198117
rect 57697 198112 60062 198114
rect 57697 198056 57702 198112
rect 57758 198056 60062 198112
rect 57697 198054 60062 198056
rect 57697 198051 57763 198054
rect 60002 198046 60062 198054
rect 217777 198112 219450 198114
rect 217777 198056 217782 198112
rect 217838 198076 219450 198112
rect 377673 198112 379530 198114
rect 217838 198056 220064 198076
rect 217777 198054 220064 198056
rect 217777 198051 217843 198054
rect 219390 198016 220064 198054
rect 377673 198056 377678 198112
rect 377734 198076 379530 198112
rect 377734 198056 380052 198076
rect 377673 198054 380052 198056
rect 377673 198051 377739 198054
rect 379470 198016 380052 198054
rect 57329 197026 57395 197029
rect 217501 197026 217567 197029
rect 377857 197026 377923 197029
rect 57329 197024 60062 197026
rect 57329 196968 57334 197024
rect 57390 196968 60062 197024
rect 57329 196966 60062 196968
rect 57329 196963 57395 196966
rect 60002 196958 60062 196966
rect 217501 197024 219450 197026
rect 217501 196968 217506 197024
rect 217562 196988 219450 197024
rect 377857 197024 379530 197026
rect 217562 196968 220064 196988
rect 217501 196966 220064 196968
rect 217501 196963 217567 196966
rect 219390 196928 220064 196966
rect 377857 196968 377862 197024
rect 377918 196988 379530 197024
rect 377918 196968 380052 196988
rect 377857 196966 380052 196968
rect 377857 196963 377923 196966
rect 379470 196928 380052 196966
rect 57053 195258 57119 195261
rect 57789 195258 57855 195261
rect 216949 195258 217015 195261
rect 217685 195258 217751 195261
rect 377305 195258 377371 195261
rect 377765 195258 377831 195261
rect 57053 195256 60062 195258
rect 57053 195200 57058 195256
rect 57114 195200 57794 195256
rect 57850 195200 60062 195256
rect 57053 195198 60062 195200
rect 57053 195195 57119 195198
rect 57789 195195 57855 195198
rect 60002 195190 60062 195198
rect 216949 195256 219450 195258
rect 216949 195200 216954 195256
rect 217010 195200 217690 195256
rect 217746 195220 219450 195256
rect 377305 195256 379530 195258
rect 217746 195200 220064 195220
rect 216949 195198 220064 195200
rect 216949 195195 217015 195198
rect 217685 195195 217751 195198
rect 219390 195160 220064 195198
rect 377305 195200 377310 195256
rect 377366 195200 377770 195256
rect 377826 195220 379530 195256
rect 377826 195200 380052 195220
rect 377305 195198 380052 195200
rect 377305 195195 377371 195198
rect 377765 195195 377831 195198
rect 379470 195160 380052 195198
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 199285 186418 199351 186421
rect 358813 186418 358879 186421
rect 359273 186418 359339 186421
rect 518893 186418 518959 186421
rect 519353 186418 519419 186421
rect 196558 186416 199351 186418
rect 196558 186360 199290 186416
rect 199346 186360 199351 186416
rect 196558 186358 199351 186360
rect 196558 186350 196618 186358
rect 199285 186355 199351 186358
rect 356562 186416 359339 186418
rect 356562 186360 358818 186416
rect 358874 186360 359278 186416
rect 359334 186360 359339 186416
rect 356562 186358 359339 186360
rect 356562 186350 356622 186358
rect 358813 186355 358879 186358
rect 359273 186355 359339 186358
rect 516558 186416 519419 186418
rect 516558 186360 518898 186416
rect 518954 186360 519358 186416
rect 519414 186360 519419 186416
rect 516558 186358 519419 186360
rect 516558 186350 516618 186358
rect 518893 186355 518959 186358
rect 519353 186355 519419 186358
rect 199009 184922 199075 184925
rect 359089 184922 359155 184925
rect 196558 184920 199075 184922
rect 196558 184864 199014 184920
rect 199070 184864 199075 184920
rect 196558 184862 199075 184864
rect 196558 184718 196618 184862
rect 199009 184859 199075 184862
rect 356562 184920 359155 184922
rect 356562 184864 359094 184920
rect 359150 184864 359155 184920
rect 356562 184862 359155 184864
rect 356562 184718 356622 184862
rect 359089 184859 359155 184862
rect 519629 184786 519695 184789
rect 520181 184786 520247 184789
rect 516558 184784 520247 184786
rect 516558 184728 519634 184784
rect 519690 184728 520186 184784
rect 520242 184728 520247 184784
rect 516558 184726 520247 184728
rect 516558 184718 516618 184726
rect 519629 184723 519695 184726
rect 520181 184723 520247 184726
rect 199009 183562 199075 183565
rect 199193 183562 199259 183565
rect 196558 183560 199259 183562
rect 196558 183504 199014 183560
rect 199070 183504 199198 183560
rect 199254 183504 199259 183560
rect 196558 183502 199259 183504
rect 196558 183358 196618 183502
rect 199009 183499 199075 183502
rect 199193 183499 199259 183502
rect 359365 183426 359431 183429
rect 519445 183426 519511 183429
rect 520089 183426 520155 183429
rect 356562 183424 359431 183426
rect 356562 183368 359370 183424
rect 359426 183368 359431 183424
rect 356562 183366 359431 183368
rect 356562 183358 356622 183366
rect 359365 183363 359431 183366
rect 516558 183424 520155 183426
rect 516558 183368 519450 183424
rect 519506 183368 520094 183424
rect 520150 183368 520155 183424
rect 516558 183366 520155 183368
rect 516558 183358 516618 183366
rect 519445 183363 519511 183366
rect 520089 183363 520155 183366
rect 358997 182066 359063 182069
rect 359273 182066 359339 182069
rect 356562 182064 359339 182066
rect 356562 182008 359002 182064
rect 359058 182008 359278 182064
rect 359334 182008 359339 182064
rect 356562 182006 359339 182008
rect 198733 181930 198799 181933
rect 196558 181928 198799 181930
rect 196558 181872 198738 181928
rect 198794 181872 198799 181928
rect 196558 181870 198799 181872
rect 196558 181862 196618 181870
rect 198733 181867 198799 181870
rect 356562 181862 356622 182006
rect 358997 182003 359063 182006
rect 359273 182003 359339 182006
rect 519169 181930 519235 181933
rect 519353 181930 519419 181933
rect 516558 181928 519419 181930
rect 516558 181872 519174 181928
rect 519230 181872 519358 181928
rect 519414 181872 519419 181928
rect 516558 181870 519419 181872
rect 516558 181862 516618 181870
rect 519169 181867 519235 181870
rect 519353 181867 519419 181870
rect 199193 180706 199259 180709
rect 359181 180706 359247 180709
rect 518985 180706 519051 180709
rect 196558 180704 199259 180706
rect 196558 180648 199198 180704
rect 199254 180648 199259 180704
rect 196558 180646 199259 180648
rect 196558 180638 196618 180646
rect 199193 180643 199259 180646
rect 356562 180704 359247 180706
rect 356562 180648 359186 180704
rect 359242 180648 359247 180704
rect 356562 180646 359247 180648
rect 356562 180638 356622 180646
rect 359181 180643 359247 180646
rect 516558 180704 519051 180706
rect 516558 180648 518990 180704
rect 519046 180648 519051 180704
rect 516558 180646 519051 180648
rect 516558 180638 516618 180646
rect 518985 180643 519051 180646
rect 583520 179060 584960 179300
rect 58801 177578 58867 177581
rect 58801 177576 60062 177578
rect 58801 177520 58806 177576
rect 58862 177520 60062 177576
rect 58801 177518 60062 177520
rect 58801 177515 58867 177518
rect 60002 176966 60062 177518
rect 216765 177034 216831 177037
rect 376937 177034 377003 177037
rect 216765 177032 219450 177034
rect 216765 176976 216770 177032
rect 216826 176996 219450 177032
rect 376937 177032 379530 177034
rect 216826 176976 220064 176996
rect 216765 176974 220064 176976
rect 216765 176971 216831 176974
rect 219390 176936 220064 176974
rect 376937 176976 376942 177032
rect 376998 176996 379530 177032
rect 376998 176976 380052 176996
rect 376937 176974 380052 176976
rect 376937 176971 377003 176974
rect 379470 176936 380052 176974
rect -960 175796 480 176036
rect 57881 175810 57947 175813
rect 57881 175808 60062 175810
rect 57881 175752 57886 175808
rect 57942 175752 60062 175808
rect 57881 175750 60062 175752
rect 57881 175747 57947 175750
rect 60002 175334 60062 175750
rect 216673 175402 216739 175405
rect 376937 175402 377003 175405
rect 216673 175400 219450 175402
rect 216673 175344 216678 175400
rect 216734 175364 219450 175400
rect 376937 175400 379530 175402
rect 216734 175344 220064 175364
rect 216673 175342 220064 175344
rect 216673 175339 216739 175342
rect 219390 175304 220064 175342
rect 376937 175344 376942 175400
rect 376998 175364 379530 175400
rect 376998 175344 380052 175364
rect 376937 175342 380052 175344
rect 376937 175339 377003 175342
rect 379470 175304 380052 175342
rect 57053 175130 57119 175133
rect 217041 175130 217107 175133
rect 376937 175130 377003 175133
rect 57053 175128 59554 175130
rect 57053 175072 57058 175128
rect 57114 175092 59554 175128
rect 217041 175128 219450 175130
rect 57114 175072 60032 175092
rect 57053 175070 60032 175072
rect 57053 175067 57119 175070
rect 59494 175032 60032 175070
rect 217041 175072 217046 175128
rect 217102 175092 219450 175128
rect 376937 175128 379530 175130
rect 217102 175072 220064 175092
rect 217041 175070 220064 175072
rect 217041 175067 217107 175070
rect 219390 175032 220064 175070
rect 376937 175072 376942 175128
rect 376998 175092 379530 175128
rect 376998 175072 380052 175092
rect 376937 175070 380052 175072
rect 376937 175067 377003 175070
rect 379470 175032 380052 175070
rect 57830 166908 57836 166972
rect 57900 166970 57906 166972
rect 57900 166910 143572 166970
rect 57900 166908 57906 166910
rect 98453 166836 98519 166837
rect 101029 166836 101095 166837
rect 105813 166836 105879 166837
rect 108205 166836 108271 166837
rect 138473 166836 138539 166837
rect 140865 166836 140931 166837
rect 143512 166836 143572 166910
rect 198038 166908 198044 166972
rect 198108 166970 198114 166972
rect 198108 166910 313500 166970
rect 198108 166908 198114 166910
rect 145925 166836 145991 166837
rect 313440 166836 313500 166910
rect 370630 166908 370636 166972
rect 370700 166970 370706 166972
rect 370700 166910 473500 166970
rect 370700 166908 370706 166910
rect 418429 166836 418495 166837
rect 421005 166836 421071 166837
rect 423397 166836 423463 166837
rect 428181 166836 428247 166837
rect 445845 166836 445911 166837
rect 470961 166836 471027 166837
rect 473440 166836 473500 166910
rect 475837 166836 475903 166837
rect 478413 166836 478479 166837
rect 480897 166836 480963 166837
rect 47894 166772 47900 166836
rect 47964 166834 47970 166836
rect 93710 166834 93716 166836
rect 47964 166774 93716 166834
rect 47964 166772 47970 166774
rect 93710 166772 93716 166774
rect 93780 166772 93786 166836
rect 98453 166834 98500 166836
rect 98408 166832 98500 166834
rect 98408 166776 98458 166832
rect 98408 166774 98500 166776
rect 98453 166772 98500 166774
rect 98564 166772 98570 166836
rect 101029 166834 101076 166836
rect 100984 166832 101076 166834
rect 100984 166776 101034 166832
rect 100984 166774 101076 166776
rect 101029 166772 101076 166774
rect 101140 166772 101146 166836
rect 105813 166834 105860 166836
rect 105768 166832 105860 166834
rect 105768 166776 105818 166832
rect 105768 166774 105860 166776
rect 105813 166772 105860 166774
rect 105924 166772 105930 166836
rect 108205 166834 108252 166836
rect 108160 166832 108252 166834
rect 108160 166776 108210 166832
rect 108160 166774 108252 166776
rect 108205 166772 108252 166774
rect 108316 166772 108322 166836
rect 138472 166772 138478 166836
rect 138542 166834 138548 166836
rect 138542 166774 138630 166834
rect 140865 166832 140926 166836
rect 140865 166776 140870 166832
rect 138542 166772 138548 166774
rect 140865 166772 140926 166776
rect 140990 166834 140996 166836
rect 140990 166774 141022 166834
rect 140990 166772 140996 166774
rect 143504 166772 143510 166836
rect 143574 166772 143580 166836
rect 145925 166832 145958 166836
rect 146022 166834 146028 166836
rect 145925 166776 145930 166832
rect 145925 166772 145958 166776
rect 146022 166774 146082 166834
rect 146022 166772 146028 166774
rect 205030 166772 205036 166836
rect 205100 166834 205106 166836
rect 305952 166834 305958 166836
rect 205100 166774 305958 166834
rect 205100 166772 205106 166774
rect 305952 166772 305958 166774
rect 306022 166772 306028 166836
rect 313432 166772 313438 166836
rect 313502 166772 313508 166836
rect 418429 166834 418476 166836
rect 418384 166832 418476 166834
rect 418384 166776 418434 166832
rect 418384 166774 418476 166776
rect 418429 166772 418476 166774
rect 418540 166772 418546 166836
rect 421005 166834 421052 166836
rect 420960 166832 421052 166834
rect 420960 166776 421010 166832
rect 420960 166774 421052 166776
rect 421005 166772 421052 166774
rect 421116 166772 421122 166836
rect 423397 166834 423444 166836
rect 423352 166832 423444 166834
rect 423352 166776 423402 166832
rect 423352 166774 423444 166776
rect 423397 166772 423444 166774
rect 423508 166772 423514 166836
rect 428181 166834 428228 166836
rect 428136 166832 428228 166834
rect 428136 166776 428186 166832
rect 428136 166774 428228 166776
rect 428181 166772 428228 166774
rect 428292 166772 428298 166836
rect 445845 166834 445892 166836
rect 445800 166832 445892 166834
rect 445800 166776 445850 166832
rect 445800 166774 445892 166776
rect 445845 166772 445892 166774
rect 445956 166772 445962 166836
rect 470961 166832 470990 166836
rect 471054 166834 471060 166836
rect 470961 166776 470966 166832
rect 470961 166772 470990 166776
rect 471054 166774 471118 166834
rect 471054 166772 471060 166774
rect 473432 166772 473438 166836
rect 473502 166772 473508 166836
rect 475837 166832 475886 166836
rect 475950 166834 475956 166836
rect 475837 166776 475842 166832
rect 475837 166772 475886 166776
rect 475950 166774 475994 166834
rect 478413 166832 478470 166836
rect 478534 166834 478540 166836
rect 478413 166776 478418 166832
rect 475950 166772 475956 166774
rect 478413 166772 478470 166776
rect 478534 166774 478570 166834
rect 480897 166832 480918 166836
rect 480982 166834 480988 166836
rect 480897 166776 480902 166832
rect 478534 166772 478540 166774
rect 480897 166772 480918 166776
rect 480982 166774 481054 166834
rect 480982 166772 480988 166774
rect 98453 166771 98519 166772
rect 101029 166771 101095 166772
rect 105813 166771 105879 166772
rect 108205 166771 108271 166772
rect 138473 166771 138539 166772
rect 140865 166771 140931 166772
rect 145925 166771 145991 166772
rect 418429 166771 418495 166772
rect 421005 166771 421071 166772
rect 423397 166771 423463 166772
rect 428181 166771 428247 166772
rect 445845 166771 445911 166772
rect 470961 166771 471027 166772
rect 475837 166771 475903 166772
rect 478413 166771 478479 166772
rect 480897 166771 480963 166772
rect 163313 166700 163379 166701
rect 165889 166700 165955 166701
rect 303521 166700 303587 166701
rect 483381 166700 483447 166701
rect 485957 166700 486023 166701
rect 163313 166696 163366 166700
rect 163430 166698 163436 166700
rect 163313 166640 163318 166696
rect 163313 166636 163366 166640
rect 163430 166638 163470 166698
rect 165889 166696 165950 166700
rect 165889 166640 165894 166696
rect 163430 166636 163436 166638
rect 165889 166636 165950 166640
rect 166014 166698 166020 166700
rect 166014 166638 166046 166698
rect 166014 166636 166020 166638
rect 213494 166636 213500 166700
rect 213564 166698 213570 166700
rect 298472 166698 298478 166700
rect 213564 166638 298478 166698
rect 213564 166636 213570 166638
rect 298472 166636 298478 166638
rect 298542 166636 298548 166700
rect 303504 166698 303510 166700
rect 303430 166638 303510 166698
rect 303574 166696 303587 166700
rect 483360 166698 483366 166700
rect 303582 166640 303587 166696
rect 303504 166636 303510 166638
rect 303574 166636 303587 166640
rect 483290 166638 483366 166698
rect 483430 166696 483447 166700
rect 485944 166698 485950 166700
rect 483442 166640 483447 166696
rect 483360 166636 483366 166638
rect 483430 166636 483447 166640
rect 485866 166638 485950 166698
rect 486014 166696 486023 166700
rect 486018 166640 486023 166696
rect 485944 166636 485950 166638
rect 486014 166636 486023 166640
rect 163313 166635 163379 166636
rect 165889 166635 165955 166636
rect 303521 166635 303587 166636
rect 483381 166635 483447 166636
rect 485957 166635 486023 166636
rect 114369 166564 114435 166565
rect 116945 166564 117011 166565
rect 148501 166564 148567 166565
rect 153285 166564 153351 166565
rect 183277 166564 183343 166565
rect 285949 166564 286015 166565
rect 288249 166564 288315 166565
rect 293401 166564 293467 166565
rect 295885 166564 295951 166565
rect 503253 166564 503319 166565
rect 114369 166560 114406 166564
rect 114470 166562 114476 166564
rect 114369 166504 114374 166560
rect 114369 166500 114406 166504
rect 114470 166502 114526 166562
rect 116945 166560 116990 166564
rect 117054 166562 117060 166564
rect 148501 166562 148548 166564
rect 116945 166504 116950 166560
rect 114470 166500 114476 166502
rect 116945 166500 116990 166504
rect 117054 166502 117102 166562
rect 148456 166560 148548 166562
rect 148456 166504 148506 166560
rect 148456 166502 148548 166504
rect 117054 166500 117060 166502
rect 148501 166500 148548 166502
rect 148612 166500 148618 166564
rect 153285 166562 153332 166564
rect 153240 166560 153332 166562
rect 153240 166504 153290 166560
rect 153240 166502 153332 166504
rect 153285 166500 153332 166502
rect 153396 166500 153402 166564
rect 183216 166562 183222 166564
rect 183186 166502 183222 166562
rect 183286 166560 183343 166564
rect 183338 166504 183343 166560
rect 183216 166500 183222 166502
rect 183286 166500 183343 166504
rect 207974 166500 207980 166564
rect 208044 166562 208050 166564
rect 208044 166502 273270 166562
rect 208044 166500 208050 166502
rect 114369 166499 114435 166500
rect 116945 166499 117011 166500
rect 148501 166499 148567 166500
rect 153285 166499 153351 166500
rect 183277 166499 183343 166500
rect 260925 166428 260991 166429
rect 265893 166428 265959 166429
rect 196566 166364 196572 166428
rect 196636 166426 196642 166428
rect 260925 166426 260972 166428
rect 196636 166366 253950 166426
rect 260880 166424 260972 166426
rect 260880 166368 260930 166424
rect 260880 166366 260972 166368
rect 196636 166364 196642 166366
rect 96061 166292 96127 166293
rect 96061 166290 96108 166292
rect 96016 166288 96108 166290
rect 96016 166232 96066 166288
rect 96016 166230 96108 166232
rect 96061 166228 96108 166230
rect 96172 166228 96178 166292
rect 253890 166290 253950 166366
rect 260925 166364 260972 166366
rect 261036 166364 261042 166428
rect 265893 166426 265940 166428
rect 265848 166424 265940 166426
rect 265848 166368 265898 166424
rect 265848 166366 265940 166368
rect 265893 166364 265940 166366
rect 266004 166364 266010 166428
rect 273210 166426 273270 166502
rect 285949 166560 285966 166564
rect 286030 166562 286036 166564
rect 285949 166504 285954 166560
rect 285949 166500 285966 166504
rect 286030 166502 286106 166562
rect 288249 166560 288278 166564
rect 288342 166562 288348 166564
rect 288249 166504 288254 166560
rect 286030 166500 286036 166502
rect 288249 166500 288278 166504
rect 288342 166502 288406 166562
rect 288342 166500 288348 166502
rect 290992 166500 290998 166564
rect 291062 166500 291068 166564
rect 293401 166560 293446 166564
rect 293510 166562 293516 166564
rect 293401 166504 293406 166560
rect 293401 166500 293446 166504
rect 293510 166502 293558 166562
rect 295885 166560 295894 166564
rect 295958 166562 295964 166564
rect 503216 166562 503222 166564
rect 295885 166504 295890 166560
rect 293510 166500 293516 166502
rect 295885 166500 295894 166504
rect 295958 166502 296042 166562
rect 503162 166502 503222 166562
rect 503286 166560 503319 166564
rect 503314 166504 503319 166560
rect 295958 166500 295964 166502
rect 503216 166500 503222 166502
rect 503286 166500 503319 166504
rect 285949 166499 286015 166500
rect 288249 166499 288315 166500
rect 291000 166426 291060 166500
rect 293401 166499 293467 166500
rect 295885 166499 295951 166500
rect 503253 166499 503319 166500
rect 273210 166366 291060 166426
rect 260925 166363 260991 166364
rect 265893 166363 265959 166364
rect 270902 166290 270908 166292
rect 253890 166230 270908 166290
rect 270902 166228 270908 166230
rect 270972 166228 270978 166292
rect 96061 166227 96127 166228
rect 583520 165732 584960 165972
rect 81433 165610 81499 165613
rect 81750 165610 81756 165612
rect 81433 165608 81756 165610
rect 81433 165552 81438 165608
rect 81494 165552 81756 165608
rect 81433 165550 81756 165552
rect 81433 165547 81499 165550
rect 81750 165548 81756 165550
rect 81820 165548 81826 165612
rect 84193 165610 84259 165613
rect 85430 165610 85436 165612
rect 84193 165608 85436 165610
rect 84193 165552 84198 165608
rect 84254 165552 85436 165608
rect 84193 165550 85436 165552
rect 84193 165547 84259 165550
rect 85430 165548 85436 165550
rect 85500 165548 85506 165612
rect 89989 165610 90055 165613
rect 90766 165610 90772 165612
rect 89989 165608 90772 165610
rect 89989 165552 89994 165608
rect 90050 165552 90772 165608
rect 89989 165550 90772 165552
rect 89989 165547 90055 165550
rect 90766 165548 90772 165550
rect 90836 165548 90842 165612
rect 91093 165610 91159 165613
rect 92422 165610 92428 165612
rect 91093 165608 92428 165610
rect 91093 165552 91098 165608
rect 91154 165552 92428 165608
rect 91093 165550 92428 165552
rect 91093 165547 91159 165550
rect 92422 165548 92428 165550
rect 92492 165548 92498 165612
rect 95233 165610 95299 165613
rect 99373 165612 99439 165613
rect 103513 165612 103579 165613
rect 95734 165610 95740 165612
rect 95233 165608 95740 165610
rect 95233 165552 95238 165608
rect 95294 165552 95740 165608
rect 95233 165550 95740 165552
rect 95233 165547 95299 165550
rect 95734 165548 95740 165550
rect 95804 165548 95810 165612
rect 99373 165608 99420 165612
rect 99484 165610 99490 165612
rect 99373 165552 99378 165608
rect 99373 165548 99420 165552
rect 99484 165550 99530 165610
rect 99484 165548 99490 165550
rect 103462 165548 103468 165612
rect 103532 165610 103579 165612
rect 109493 165610 109559 165613
rect 109718 165610 109724 165612
rect 103532 165608 103624 165610
rect 103574 165552 103624 165608
rect 103532 165550 103624 165552
rect 109493 165608 109724 165610
rect 109493 165552 109498 165608
rect 109554 165552 109724 165608
rect 109493 165550 109724 165552
rect 103532 165548 103579 165550
rect 99373 165547 99439 165548
rect 103513 165547 103579 165548
rect 109493 165547 109559 165550
rect 109718 165548 109724 165550
rect 109788 165548 109794 165612
rect 110873 165610 110939 165613
rect 111149 165612 111215 165613
rect 111006 165610 111012 165612
rect 110873 165608 111012 165610
rect 110873 165552 110878 165608
rect 110934 165552 111012 165608
rect 110873 165550 111012 165552
rect 110873 165547 110939 165550
rect 111006 165548 111012 165550
rect 111076 165548 111082 165612
rect 111149 165608 111196 165612
rect 111260 165610 111266 165612
rect 111149 165552 111154 165608
rect 111149 165548 111196 165552
rect 111260 165550 111306 165610
rect 111260 165548 111266 165550
rect 112294 165548 112300 165612
rect 112364 165610 112370 165612
rect 113173 165610 113239 165613
rect 112364 165608 113239 165610
rect 112364 165552 113178 165608
rect 113234 165552 113239 165608
rect 112364 165550 113239 165552
rect 112364 165548 112370 165550
rect 111149 165547 111215 165548
rect 113173 165547 113239 165550
rect 113541 165612 113607 165613
rect 115933 165612 115999 165613
rect 117957 165612 118023 165613
rect 118325 165612 118391 165613
rect 113541 165608 113588 165612
rect 113652 165610 113658 165612
rect 113541 165552 113546 165608
rect 113541 165548 113588 165552
rect 113652 165550 113698 165610
rect 115933 165608 115980 165612
rect 116044 165610 116050 165612
rect 115933 165552 115938 165608
rect 113652 165548 113658 165550
rect 115933 165548 115980 165552
rect 116044 165550 116090 165610
rect 117957 165608 118004 165612
rect 118068 165610 118074 165612
rect 117957 165552 117962 165608
rect 116044 165548 116050 165550
rect 117957 165548 118004 165552
rect 118068 165550 118114 165610
rect 118325 165608 118372 165612
rect 118436 165610 118442 165612
rect 118969 165610 119035 165613
rect 120901 165612 120967 165613
rect 123477 165612 123543 165613
rect 125869 165612 125935 165613
rect 119102 165610 119108 165612
rect 118325 165552 118330 165608
rect 118068 165548 118074 165550
rect 118325 165548 118372 165552
rect 118436 165550 118482 165610
rect 118969 165608 119108 165610
rect 118969 165552 118974 165608
rect 119030 165552 119108 165608
rect 118969 165550 119108 165552
rect 118436 165548 118442 165550
rect 113541 165547 113607 165548
rect 115933 165547 115999 165548
rect 117957 165547 118023 165548
rect 118325 165547 118391 165548
rect 118969 165547 119035 165550
rect 119102 165548 119108 165550
rect 119172 165548 119178 165612
rect 120901 165608 120948 165612
rect 121012 165610 121018 165612
rect 120901 165552 120906 165608
rect 120901 165548 120948 165552
rect 121012 165550 121058 165610
rect 123477 165608 123524 165612
rect 123588 165610 123594 165612
rect 123477 165552 123482 165608
rect 121012 165548 121018 165550
rect 123477 165548 123524 165552
rect 123588 165550 123634 165610
rect 125869 165608 125916 165612
rect 125980 165610 125986 165612
rect 128353 165610 128419 165613
rect 128486 165610 128492 165612
rect 125869 165552 125874 165608
rect 123588 165548 123594 165550
rect 125869 165548 125916 165552
rect 125980 165550 126026 165610
rect 128353 165608 128492 165610
rect 128353 165552 128358 165608
rect 128414 165552 128492 165608
rect 128353 165550 128492 165552
rect 125980 165548 125986 165550
rect 120901 165547 120967 165548
rect 123477 165547 123543 165548
rect 125869 165547 125935 165548
rect 128353 165547 128419 165550
rect 128486 165548 128492 165550
rect 128556 165548 128562 165612
rect 129733 165610 129799 165613
rect 130878 165610 130884 165612
rect 129733 165608 130884 165610
rect 129733 165552 129738 165608
rect 129794 165552 130884 165608
rect 129733 165550 130884 165552
rect 129733 165547 129799 165550
rect 130878 165548 130884 165550
rect 130948 165548 130954 165612
rect 132493 165610 132559 165613
rect 183369 165612 183435 165613
rect 235993 165612 236059 165613
rect 133454 165610 133460 165612
rect 132493 165608 133460 165610
rect 132493 165552 132498 165608
rect 132554 165552 133460 165608
rect 132493 165550 133460 165552
rect 132493 165547 132559 165550
rect 133454 165548 133460 165550
rect 133524 165548 133530 165612
rect 183318 165548 183324 165612
rect 183388 165610 183435 165612
rect 183388 165608 183480 165610
rect 183430 165552 183480 165608
rect 183388 165550 183480 165552
rect 183388 165548 183435 165550
rect 235942 165548 235948 165612
rect 236012 165610 236059 165612
rect 238753 165610 238819 165613
rect 239622 165610 239628 165612
rect 236012 165608 236104 165610
rect 236054 165552 236104 165608
rect 236012 165550 236104 165552
rect 238753 165608 239628 165610
rect 238753 165552 238758 165608
rect 238814 165552 239628 165608
rect 238753 165550 239628 165552
rect 236012 165548 236059 165550
rect 183369 165547 183435 165548
rect 235993 165547 236059 165548
rect 238753 165547 238819 165550
rect 239622 165548 239628 165550
rect 239692 165548 239698 165612
rect 242893 165610 242959 165613
rect 243118 165610 243124 165612
rect 242893 165608 243124 165610
rect 242893 165552 242898 165608
rect 242954 165552 243124 165608
rect 242893 165550 243124 165552
rect 242893 165547 242959 165550
rect 243118 165548 243124 165550
rect 243188 165548 243194 165612
rect 247033 165610 247099 165613
rect 247534 165610 247540 165612
rect 247033 165608 247540 165610
rect 247033 165552 247038 165608
rect 247094 165552 247540 165608
rect 247033 165550 247540 165552
rect 247033 165547 247099 165550
rect 247534 165548 247540 165550
rect 247604 165548 247610 165612
rect 247677 165610 247743 165613
rect 248270 165610 248276 165612
rect 247677 165608 248276 165610
rect 247677 165552 247682 165608
rect 247738 165552 248276 165608
rect 247677 165550 248276 165552
rect 247677 165547 247743 165550
rect 248270 165548 248276 165550
rect 248340 165548 248346 165612
rect 249793 165610 249859 165613
rect 250662 165610 250668 165612
rect 249793 165608 250668 165610
rect 249793 165552 249798 165608
rect 249854 165552 250668 165608
rect 249793 165550 250668 165552
rect 249793 165547 249859 165550
rect 250662 165548 250668 165550
rect 250732 165548 250738 165612
rect 252553 165610 252619 165613
rect 253606 165610 253612 165612
rect 252553 165608 253612 165610
rect 252553 165552 252558 165608
rect 252614 165552 253612 165608
rect 252553 165550 253612 165552
rect 252553 165547 252619 165550
rect 253606 165548 253612 165550
rect 253676 165548 253682 165612
rect 258073 165610 258139 165613
rect 258390 165610 258396 165612
rect 258073 165608 258396 165610
rect 258073 165552 258078 165608
rect 258134 165552 258396 165608
rect 258073 165550 258396 165552
rect 258073 165547 258139 165550
rect 258390 165548 258396 165550
rect 258460 165548 258466 165612
rect 260833 165610 260899 165613
rect 261702 165610 261708 165612
rect 260833 165608 261708 165610
rect 260833 165552 260838 165608
rect 260894 165552 261708 165608
rect 260833 165550 261708 165552
rect 260833 165547 260899 165550
rect 261702 165548 261708 165550
rect 261772 165548 261778 165612
rect 264973 165610 265039 165613
rect 265198 165610 265204 165612
rect 264973 165608 265204 165610
rect 264973 165552 264978 165608
rect 265034 165552 265204 165608
rect 264973 165550 265204 165552
rect 264973 165547 265039 165550
rect 265198 165548 265204 165550
rect 265268 165548 265274 165612
rect 267733 165610 267799 165613
rect 268326 165610 268332 165612
rect 267733 165608 268332 165610
rect 267733 165552 267738 165608
rect 267794 165552 268332 165608
rect 267733 165550 268332 165552
rect 267733 165547 267799 165550
rect 268326 165548 268332 165550
rect 268396 165548 268402 165612
rect 271873 165610 271939 165613
rect 273437 165612 273503 165613
rect 275921 165612 275987 165613
rect 272190 165610 272196 165612
rect 271873 165608 272196 165610
rect 271873 165552 271878 165608
rect 271934 165552 272196 165608
rect 271873 165550 272196 165552
rect 271873 165547 271939 165550
rect 272190 165548 272196 165550
rect 272260 165548 272266 165612
rect 273437 165610 273484 165612
rect 273392 165608 273484 165610
rect 273392 165552 273442 165608
rect 273392 165550 273484 165552
rect 273437 165548 273484 165550
rect 273548 165548 273554 165612
rect 275870 165610 275876 165612
rect 275830 165550 275876 165610
rect 275940 165608 275987 165612
rect 275982 165552 275987 165608
rect 275870 165548 275876 165550
rect 275940 165548 275987 165552
rect 276054 165548 276060 165612
rect 276124 165610 276130 165612
rect 276197 165610 276263 165613
rect 276124 165608 276263 165610
rect 276124 165552 276202 165608
rect 276258 165552 276263 165608
rect 276124 165550 276263 165552
rect 276124 165548 276130 165550
rect 273437 165547 273503 165548
rect 275921 165547 275987 165548
rect 276197 165547 276263 165550
rect 277393 165610 277459 165613
rect 278446 165610 278452 165612
rect 277393 165608 278452 165610
rect 277393 165552 277398 165608
rect 277454 165552 278452 165608
rect 277393 165550 278452 165552
rect 277393 165547 277459 165550
rect 278446 165548 278452 165550
rect 278516 165548 278522 165612
rect 279182 165548 279188 165612
rect 279252 165610 279258 165612
rect 280061 165610 280127 165613
rect 279252 165608 280127 165610
rect 279252 165552 280066 165608
rect 280122 165552 280127 165608
rect 279252 165550 280127 165552
rect 279252 165548 279258 165550
rect 280061 165547 280127 165550
rect 280245 165610 280311 165613
rect 283373 165612 283439 165613
rect 300853 165612 300919 165613
rect 323301 165612 323367 165613
rect 343449 165612 343515 165613
rect 280838 165610 280844 165612
rect 280245 165608 280844 165610
rect 280245 165552 280250 165608
rect 280306 165552 280844 165608
rect 280245 165550 280844 165552
rect 280245 165547 280311 165550
rect 280838 165548 280844 165550
rect 280908 165548 280914 165612
rect 283373 165608 283420 165612
rect 283484 165610 283490 165612
rect 283373 165552 283378 165608
rect 283373 165548 283420 165552
rect 283484 165550 283530 165610
rect 300853 165608 300900 165612
rect 300964 165610 300970 165612
rect 300853 165552 300858 165608
rect 283484 165548 283490 165550
rect 300853 165548 300900 165552
rect 300964 165550 301010 165610
rect 323301 165608 323348 165612
rect 323412 165610 323418 165612
rect 343398 165610 343404 165612
rect 323301 165552 323306 165608
rect 300964 165548 300970 165550
rect 323301 165548 323348 165552
rect 323412 165550 323458 165610
rect 343358 165550 343404 165610
rect 343468 165608 343515 165612
rect 343510 165552 343515 165608
rect 323412 165548 323418 165550
rect 343398 165548 343404 165550
rect 343468 165548 343515 165552
rect 283373 165547 283439 165548
rect 300853 165547 300919 165548
rect 323301 165547 323367 165548
rect 343449 165547 343515 165548
rect 376293 165610 376359 165613
rect 380525 165610 380591 165613
rect 376293 165608 380591 165610
rect 376293 165552 376298 165608
rect 376354 165552 380530 165608
rect 380586 165552 380591 165608
rect 376293 165550 380591 165552
rect 376293 165547 376359 165550
rect 380525 165547 380591 165550
rect 397453 165610 397519 165613
rect 398230 165610 398236 165612
rect 397453 165608 398236 165610
rect 397453 165552 397458 165608
rect 397514 165552 398236 165608
rect 397453 165550 398236 165552
rect 397453 165547 397519 165550
rect 398230 165548 398236 165550
rect 398300 165548 398306 165612
rect 401593 165610 401659 165613
rect 401726 165610 401732 165612
rect 401593 165608 401732 165610
rect 401593 165552 401598 165608
rect 401654 165552 401732 165608
rect 401593 165550 401732 165552
rect 401593 165547 401659 165550
rect 401726 165548 401732 165550
rect 401796 165548 401802 165612
rect 404353 165610 404419 165613
rect 405406 165610 405412 165612
rect 404353 165608 405412 165610
rect 404353 165552 404358 165608
rect 404414 165552 405412 165608
rect 404353 165550 405412 165552
rect 404353 165547 404419 165550
rect 405406 165548 405412 165550
rect 405476 165548 405482 165612
rect 409873 165610 409939 165613
rect 410742 165610 410748 165612
rect 409873 165608 410748 165610
rect 409873 165552 409878 165608
rect 409934 165552 410748 165608
rect 409873 165550 410748 165552
rect 409873 165547 409939 165550
rect 410742 165548 410748 165550
rect 410812 165548 410818 165612
rect 415485 165610 415551 165613
rect 416037 165612 416103 165613
rect 415894 165610 415900 165612
rect 415485 165608 415900 165610
rect 415485 165552 415490 165608
rect 415546 165552 415900 165608
rect 415485 165550 415900 165552
rect 415485 165547 415551 165550
rect 415894 165548 415900 165550
rect 415964 165548 415970 165612
rect 416037 165608 416084 165612
rect 416148 165610 416154 165612
rect 418521 165610 418587 165613
rect 423765 165612 423831 165613
rect 419390 165610 419396 165612
rect 416037 165552 416042 165608
rect 416037 165548 416084 165552
rect 416148 165550 416194 165610
rect 418521 165608 419396 165610
rect 418521 165552 418526 165608
rect 418582 165552 419396 165608
rect 418521 165550 419396 165552
rect 416148 165548 416154 165550
rect 416037 165547 416103 165548
rect 418521 165547 418587 165550
rect 419390 165548 419396 165550
rect 419460 165548 419466 165612
rect 423765 165610 423812 165612
rect 423720 165608 423812 165610
rect 423720 165552 423770 165608
rect 423720 165550 423812 165552
rect 423765 165548 423812 165550
rect 423876 165548 423882 165612
rect 433425 165610 433491 165613
rect 434294 165610 434300 165612
rect 433425 165608 434300 165610
rect 433425 165552 433430 165608
rect 433486 165552 434300 165608
rect 433425 165550 434300 165552
rect 423765 165547 423831 165548
rect 433425 165547 433491 165550
rect 434294 165548 434300 165550
rect 434364 165548 434370 165612
rect 434713 165610 434779 165613
rect 435950 165610 435956 165612
rect 434713 165608 435956 165610
rect 434713 165552 434718 165608
rect 434774 165552 435956 165608
rect 434713 165550 435956 165552
rect 434713 165547 434779 165550
rect 435950 165548 435956 165550
rect 436020 165548 436026 165612
rect 436093 165610 436159 165613
rect 437749 165612 437815 165613
rect 436870 165610 436876 165612
rect 436093 165608 436876 165610
rect 436093 165552 436098 165608
rect 436154 165552 436876 165608
rect 436093 165550 436876 165552
rect 436093 165547 436159 165550
rect 436870 165548 436876 165550
rect 436940 165548 436946 165612
rect 437749 165610 437796 165612
rect 437704 165608 437796 165610
rect 437704 165552 437754 165608
rect 437704 165550 437796 165552
rect 437749 165548 437796 165550
rect 437860 165548 437866 165612
rect 438025 165610 438091 165613
rect 438526 165610 438532 165612
rect 438025 165608 438532 165610
rect 438025 165552 438030 165608
rect 438086 165552 438532 165608
rect 438025 165550 438532 165552
rect 437749 165547 437815 165548
rect 438025 165547 438091 165550
rect 438526 165548 438532 165550
rect 438596 165548 438602 165612
rect 439262 165548 439268 165612
rect 439332 165610 439338 165612
rect 440141 165610 440207 165613
rect 439332 165608 440207 165610
rect 439332 165552 440146 165608
rect 440202 165552 440207 165608
rect 439332 165550 440207 165552
rect 439332 165548 439338 165550
rect 440141 165547 440207 165550
rect 442993 165610 443059 165613
rect 443494 165610 443500 165612
rect 442993 165608 443500 165610
rect 442993 165552 442998 165608
rect 443054 165552 443500 165608
rect 442993 165550 443500 165552
rect 442993 165547 443059 165550
rect 443494 165548 443500 165550
rect 443564 165548 443570 165612
rect 447317 165610 447383 165613
rect 448278 165610 448284 165612
rect 447317 165608 448284 165610
rect 447317 165552 447322 165608
rect 447378 165552 448284 165608
rect 447317 165550 448284 165552
rect 447317 165547 447383 165550
rect 448278 165548 448284 165550
rect 448348 165548 448354 165612
rect 449893 165610 449959 165613
rect 451038 165610 451044 165612
rect 449893 165608 451044 165610
rect 449893 165552 449898 165608
rect 449954 165552 451044 165608
rect 449893 165550 451044 165552
rect 449893 165547 449959 165550
rect 451038 165548 451044 165550
rect 451108 165548 451114 165612
rect 452653 165610 452719 165613
rect 453430 165610 453436 165612
rect 452653 165608 453436 165610
rect 452653 165552 452658 165608
rect 452714 165552 453436 165608
rect 452653 165550 453436 165552
rect 452653 165547 452719 165550
rect 453430 165548 453436 165550
rect 453500 165548 453506 165612
rect 455413 165610 455479 165613
rect 458357 165612 458423 165613
rect 503345 165612 503411 165613
rect 455822 165610 455828 165612
rect 455413 165608 455828 165610
rect 455413 165552 455418 165608
rect 455474 165552 455828 165608
rect 455413 165550 455828 165552
rect 455413 165547 455479 165550
rect 455822 165548 455828 165550
rect 455892 165548 455898 165612
rect 458357 165608 458404 165612
rect 458468 165610 458474 165612
rect 458357 165552 458362 165608
rect 458357 165548 458404 165552
rect 458468 165550 458514 165610
rect 458468 165548 458474 165550
rect 503294 165548 503300 165612
rect 503364 165610 503411 165612
rect 503364 165608 503456 165610
rect 503406 165552 503456 165608
rect 503364 165550 503456 165552
rect 503364 165548 503411 165550
rect 458357 165547 458423 165548
rect 503345 165547 503411 165548
rect 49325 165474 49391 165477
rect 158478 165474 158484 165476
rect 49325 165472 158484 165474
rect 49325 165416 49330 165472
rect 49386 165416 158484 165472
rect 49325 165414 158484 165416
rect 49325 165411 49391 165414
rect 158478 165412 158484 165414
rect 158548 165412 158554 165476
rect 208894 165412 208900 165476
rect 208964 165474 208970 165476
rect 325918 165474 325924 165476
rect 208964 165414 325924 165474
rect 208964 165412 208970 165414
rect 325918 165412 325924 165414
rect 325988 165412 325994 165476
rect 343214 165412 343220 165476
rect 343284 165474 343290 165476
rect 343541 165474 343607 165477
rect 343284 165472 343607 165474
rect 343284 165416 343546 165472
rect 343602 165416 343607 165472
rect 343284 165414 343607 165416
rect 343284 165412 343290 165414
rect 343541 165411 343607 165414
rect 378961 165474 379027 165477
rect 468518 165474 468524 165476
rect 378961 165472 468524 165474
rect 378961 165416 378966 165472
rect 379022 165416 468524 165472
rect 378961 165414 468524 165416
rect 378961 165411 379027 165414
rect 468518 165412 468524 165414
rect 468588 165412 468594 165476
rect 50889 165338 50955 165341
rect 155902 165338 155908 165340
rect 50889 165336 155908 165338
rect 50889 165280 50894 165336
rect 50950 165280 155908 165336
rect 50889 165278 155908 165280
rect 50889 165275 50955 165278
rect 155902 165276 155908 165278
rect 155972 165276 155978 165340
rect 204846 165276 204852 165340
rect 204916 165338 204922 165340
rect 315798 165338 315804 165340
rect 204916 165278 315804 165338
rect 204916 165276 204922 165278
rect 315798 165276 315804 165278
rect 315868 165276 315874 165340
rect 378777 165338 378843 165341
rect 380525 165338 380591 165341
rect 463550 165338 463556 165340
rect 378777 165336 380450 165338
rect 378777 165280 378782 165336
rect 378838 165280 380450 165336
rect 378777 165278 380450 165280
rect 378777 165275 378843 165278
rect 59905 165202 59971 165205
rect 150934 165202 150940 165204
rect 59905 165200 150940 165202
rect 59905 165144 59910 165200
rect 59966 165144 150940 165200
rect 59905 165142 150940 165144
rect 59905 165139 59971 165142
rect 150934 165140 150940 165142
rect 151004 165140 151010 165204
rect 213310 165140 213316 165204
rect 213380 165202 213386 165204
rect 311014 165202 311020 165204
rect 213380 165142 311020 165202
rect 213380 165140 213386 165142
rect 311014 165140 311020 165142
rect 311084 165140 311090 165204
rect 379646 165140 379652 165204
rect 379716 165140 379722 165204
rect 380390 165202 380450 165278
rect 380525 165336 463556 165338
rect 380525 165280 380530 165336
rect 380586 165280 463556 165336
rect 380525 165278 463556 165280
rect 380525 165275 380591 165278
rect 463550 165276 463556 165278
rect 463620 165276 463626 165340
rect 460974 165202 460980 165204
rect 380390 165142 460980 165202
rect 460974 165140 460980 165142
rect 461044 165140 461050 165204
rect 56041 165066 56107 165069
rect 136030 165066 136036 165068
rect 56041 165064 136036 165066
rect 56041 165008 56046 165064
rect 56102 165008 136036 165064
rect 56041 165006 136036 165008
rect 56041 165003 56107 165006
rect 136030 165004 136036 165006
rect 136100 165004 136106 165068
rect 216254 165004 216260 165068
rect 216324 165066 216330 165068
rect 308622 165066 308628 165068
rect 216324 165006 308628 165066
rect 216324 165004 216330 165006
rect 308622 165004 308628 165006
rect 308692 165004 308698 165068
rect 379654 165066 379714 165140
rect 426014 165066 426020 165068
rect 379654 165006 426020 165066
rect 426014 165004 426020 165006
rect 426084 165004 426090 165068
rect 440325 165066 440391 165069
rect 440918 165066 440924 165068
rect 440325 165064 440924 165066
rect 440325 165008 440330 165064
rect 440386 165008 440924 165064
rect 440325 165006 440924 165008
rect 440325 165003 440391 165006
rect 440918 165004 440924 165006
rect 440988 165004 440994 165068
rect 88333 164932 88399 164933
rect 88333 164930 88380 164932
rect 88288 164928 88380 164930
rect 88288 164872 88338 164928
rect 88288 164870 88380 164872
rect 88333 164868 88380 164870
rect 88444 164868 88450 164932
rect 107653 164930 107719 164933
rect 108614 164930 108620 164932
rect 107653 164928 108620 164930
rect 107653 164872 107658 164928
rect 107714 164872 108620 164928
rect 107653 164870 108620 164872
rect 88333 164867 88399 164868
rect 107653 164867 107719 164870
rect 108614 164868 108620 164870
rect 108684 164868 108690 164932
rect 206502 164868 206508 164932
rect 206572 164930 206578 164932
rect 263726 164930 263732 164932
rect 206572 164870 263732 164930
rect 206572 164868 206578 164870
rect 263726 164868 263732 164870
rect 263796 164868 263802 164932
rect 407113 164930 407179 164933
rect 408166 164930 408172 164932
rect 407113 164928 408172 164930
rect 407113 164872 407118 164928
rect 407174 164872 408172 164928
rect 407113 164870 408172 164872
rect 407113 164867 407179 164870
rect 408166 164868 408172 164870
rect 408236 164868 408242 164932
rect 433333 164930 433399 164933
rect 433558 164930 433564 164932
rect 433333 164928 433564 164930
rect 433333 164872 433338 164928
rect 433394 164872 433564 164928
rect 433333 164870 433564 164872
rect 433333 164867 433399 164870
rect 433558 164868 433564 164870
rect 433628 164868 433634 164932
rect 106273 164794 106339 164797
rect 107510 164794 107516 164796
rect 106273 164792 107516 164794
rect 106273 164736 106278 164792
rect 106334 164736 107516 164792
rect 106273 164734 107516 164736
rect 106273 164731 106339 164734
rect 107510 164732 107516 164734
rect 107580 164732 107586 164796
rect 200982 164732 200988 164796
rect 201052 164794 201058 164796
rect 256182 164794 256188 164796
rect 201052 164734 256188 164794
rect 201052 164732 201058 164734
rect 256182 164732 256188 164734
rect 256252 164732 256258 164796
rect 412633 164794 412699 164797
rect 413686 164794 413692 164796
rect 412633 164792 413692 164794
rect 412633 164736 412638 164792
rect 412694 164736 413692 164792
rect 412633 164734 413692 164736
rect 412633 164731 412699 164734
rect 413686 164732 413692 164734
rect 413756 164732 413762 164796
rect 420913 164794 420979 164797
rect 421782 164794 421788 164796
rect 420913 164792 421788 164794
rect 420913 164736 420918 164792
rect 420974 164736 421788 164792
rect 420913 164734 421788 164736
rect 420913 164731 420979 164734
rect 421782 164732 421788 164734
rect 421852 164732 421858 164796
rect 430665 164794 430731 164797
rect 431166 164794 431172 164796
rect 430665 164792 431172 164794
rect 430665 164736 430670 164792
rect 430726 164736 431172 164792
rect 430665 164734 431172 164736
rect 430665 164731 430731 164734
rect 431166 164732 431172 164734
rect 431236 164732 431242 164796
rect 50470 164596 50476 164660
rect 50540 164658 50546 164660
rect 160870 164658 160876 164660
rect 50540 164598 160876 164658
rect 50540 164596 50546 164598
rect 160870 164596 160876 164598
rect 160940 164596 160946 164660
rect 266353 164658 266419 164661
rect 267590 164658 267596 164660
rect 266353 164656 267596 164658
rect 266353 164600 266358 164656
rect 266414 164600 267596 164656
rect 266353 164598 267596 164600
rect 266353 164595 266419 164598
rect 267590 164596 267596 164598
rect 267660 164596 267666 164660
rect 376109 164658 376175 164661
rect 465942 164658 465948 164660
rect 376109 164656 465948 164658
rect 376109 164600 376114 164656
rect 376170 164600 465948 164656
rect 376109 164598 465948 164600
rect 376109 164595 376175 164598
rect 465942 164596 465948 164598
rect 466012 164596 466018 164660
rect 100753 164524 100819 164525
rect 100702 164460 100708 164524
rect 100772 164522 100819 164524
rect 100772 164520 100864 164522
rect 100814 164464 100864 164520
rect 100772 164462 100864 164464
rect 100772 164460 100819 164462
rect 113214 164460 113220 164524
rect 113284 164522 113290 164524
rect 114553 164522 114619 164525
rect 113284 164520 114619 164522
rect 113284 164464 114558 164520
rect 114614 164464 114619 164520
rect 113284 164462 114619 164464
rect 113284 164460 113290 164462
rect 100753 164459 100819 164460
rect 114553 164459 114619 164462
rect 115790 164460 115796 164524
rect 115860 164522 115866 164524
rect 115933 164522 115999 164525
rect 115860 164520 115999 164522
rect 115860 164464 115938 164520
rect 115994 164464 115999 164520
rect 115860 164462 115999 164464
rect 115860 164460 115866 164462
rect 115933 164459 115999 164462
rect 244365 164524 244431 164525
rect 244365 164520 244412 164524
rect 244476 164522 244482 164524
rect 251265 164522 251331 164525
rect 252318 164522 252324 164524
rect 244365 164464 244370 164520
rect 244365 164460 244412 164464
rect 244476 164462 244522 164522
rect 251265 164520 252324 164522
rect 251265 164464 251270 164520
rect 251326 164464 252324 164520
rect 251265 164462 252324 164464
rect 244476 164460 244482 164462
rect 244365 164459 244431 164460
rect 251265 164459 251331 164462
rect 252318 164460 252324 164462
rect 252388 164460 252394 164524
rect 259545 164522 259611 164525
rect 260598 164522 260604 164524
rect 259545 164520 260604 164522
rect 259545 164464 259550 164520
rect 259606 164464 260604 164520
rect 259545 164462 260604 164464
rect 259545 164459 259611 164462
rect 260598 164460 260604 164462
rect 260668 164460 260674 164524
rect 266486 164460 266492 164524
rect 266556 164522 266562 164524
rect 267641 164522 267707 164525
rect 266556 164520 267707 164522
rect 266556 164464 267646 164520
rect 267702 164464 267707 164520
rect 266556 164462 267707 164464
rect 266556 164460 266562 164462
rect 267641 164459 267707 164462
rect 273294 164460 273300 164524
rect 273364 164522 273370 164524
rect 274449 164522 274515 164525
rect 273364 164520 274515 164522
rect 273364 164464 274454 164520
rect 274510 164464 274515 164520
rect 273364 164462 274515 164464
rect 273364 164460 273370 164462
rect 274449 164459 274515 164462
rect 76005 164386 76071 164389
rect 77150 164386 77156 164388
rect 76005 164384 77156 164386
rect 76005 164328 76010 164384
rect 76066 164328 77156 164384
rect 76005 164326 77156 164328
rect 76005 164323 76071 164326
rect 77150 164324 77156 164326
rect 77220 164324 77226 164388
rect 89897 164386 89963 164389
rect 90030 164386 90036 164388
rect 89897 164384 90036 164386
rect 89897 164328 89902 164384
rect 89958 164328 90036 164384
rect 89897 164326 90036 164328
rect 89897 164323 89963 164326
rect 90030 164324 90036 164326
rect 90100 164324 90106 164388
rect 202454 164324 202460 164388
rect 202524 164386 202530 164388
rect 320950 164386 320956 164388
rect 202524 164326 320956 164386
rect 202524 164324 202530 164326
rect 320950 164324 320956 164326
rect 321020 164324 321026 164388
rect 396165 164386 396231 164389
rect 397126 164386 397132 164388
rect 396165 164384 397132 164386
rect 396165 164328 396170 164384
rect 396226 164328 397132 164384
rect 396165 164326 397132 164328
rect 396165 164323 396231 164326
rect 397126 164324 397132 164326
rect 397196 164324 397202 164388
rect 402973 164386 403039 164389
rect 404118 164386 404124 164388
rect 402973 164384 404124 164386
rect 402973 164328 402978 164384
rect 403034 164328 404124 164384
rect 402973 164326 404124 164328
rect 402973 164323 403039 164326
rect 404118 164324 404124 164326
rect 404188 164324 404194 164388
rect 411253 164386 411319 164389
rect 412398 164386 412404 164388
rect 411253 164384 412404 164386
rect 411253 164328 411258 164384
rect 411314 164328 412404 164384
rect 411253 164326 412404 164328
rect 411253 164323 411319 164326
rect 412398 164324 412404 164326
rect 412468 164324 412474 164388
rect 426382 164324 426388 164388
rect 426452 164386 426458 164388
rect 426525 164386 426591 164389
rect 426452 164384 426591 164386
rect 426452 164328 426530 164384
rect 426586 164328 426591 164384
rect 426452 164326 426591 164328
rect 426452 164324 426458 164326
rect 426525 164323 426591 164326
rect 429285 164386 429351 164389
rect 429694 164386 429700 164388
rect 429285 164384 429700 164386
rect 429285 164328 429290 164384
rect 429346 164328 429700 164384
rect 429285 164326 429700 164328
rect 429285 164323 429351 164326
rect 429694 164324 429700 164326
rect 429764 164324 429770 164388
rect 75913 164250 75979 164253
rect 76046 164250 76052 164252
rect 75913 164248 76052 164250
rect 75913 164192 75918 164248
rect 75974 164192 76052 164248
rect 75913 164190 76052 164192
rect 75913 164187 75979 164190
rect 76046 164188 76052 164190
rect 76116 164188 76122 164252
rect 77293 164250 77359 164253
rect 78254 164250 78260 164252
rect 77293 164248 78260 164250
rect 77293 164192 77298 164248
rect 77354 164192 78260 164248
rect 77293 164190 78260 164192
rect 77293 164187 77359 164190
rect 78254 164188 78260 164190
rect 78324 164188 78330 164252
rect 78673 164250 78739 164253
rect 79542 164250 79548 164252
rect 78673 164248 79548 164250
rect 78673 164192 78678 164248
rect 78734 164192 79548 164248
rect 78673 164190 79548 164192
rect 78673 164187 78739 164190
rect 79542 164188 79548 164190
rect 79612 164188 79618 164252
rect 80053 164250 80119 164253
rect 80462 164250 80468 164252
rect 80053 164248 80468 164250
rect 80053 164192 80058 164248
rect 80114 164192 80468 164248
rect 80053 164190 80468 164192
rect 80053 164187 80119 164190
rect 80462 164188 80468 164190
rect 80532 164188 80538 164252
rect 82813 164250 82879 164253
rect 83038 164250 83044 164252
rect 82813 164248 83044 164250
rect 82813 164192 82818 164248
rect 82874 164192 83044 164248
rect 82813 164190 83044 164192
rect 82813 164187 82879 164190
rect 83038 164188 83044 164190
rect 83108 164188 83114 164252
rect 84142 164188 84148 164252
rect 84212 164250 84218 164252
rect 84285 164250 84351 164253
rect 84212 164248 84351 164250
rect 84212 164192 84290 164248
rect 84346 164192 84351 164248
rect 84212 164190 84351 164192
rect 84212 164188 84218 164190
rect 84285 164187 84351 164190
rect 85573 164250 85639 164253
rect 86534 164250 86540 164252
rect 85573 164248 86540 164250
rect 85573 164192 85578 164248
rect 85634 164192 86540 164248
rect 85573 164190 86540 164192
rect 85573 164187 85639 164190
rect 86534 164188 86540 164190
rect 86604 164188 86610 164252
rect 86953 164250 87019 164253
rect 87638 164250 87644 164252
rect 86953 164248 87644 164250
rect 86953 164192 86958 164248
rect 87014 164192 87644 164248
rect 86953 164190 87644 164192
rect 86953 164187 87019 164190
rect 87638 164188 87644 164190
rect 87708 164188 87714 164252
rect 88425 164250 88491 164253
rect 88742 164250 88748 164252
rect 88425 164248 88748 164250
rect 88425 164192 88430 164248
rect 88486 164192 88748 164248
rect 88425 164190 88748 164192
rect 88425 164187 88491 164190
rect 88742 164188 88748 164190
rect 88812 164188 88818 164252
rect 91185 164250 91251 164253
rect 91318 164250 91324 164252
rect 91185 164248 91324 164250
rect 91185 164192 91190 164248
rect 91246 164192 91324 164248
rect 91185 164190 91324 164192
rect 91185 164187 91251 164190
rect 91318 164188 91324 164190
rect 91388 164188 91394 164252
rect 92473 164250 92539 164253
rect 93342 164250 93348 164252
rect 92473 164248 93348 164250
rect 92473 164192 92478 164248
rect 92534 164192 93348 164248
rect 92473 164190 93348 164192
rect 92473 164187 92539 164190
rect 93342 164188 93348 164190
rect 93412 164188 93418 164252
rect 93853 164250 93919 164253
rect 94446 164250 94452 164252
rect 93853 164248 94452 164250
rect 93853 164192 93858 164248
rect 93914 164192 94452 164248
rect 93853 164190 94452 164192
rect 93853 164187 93919 164190
rect 94446 164188 94452 164190
rect 94516 164188 94522 164252
rect 96613 164250 96679 164253
rect 97022 164250 97028 164252
rect 96613 164248 97028 164250
rect 96613 164192 96618 164248
rect 96674 164192 97028 164248
rect 96613 164190 97028 164192
rect 96613 164187 96679 164190
rect 97022 164188 97028 164190
rect 97092 164188 97098 164252
rect 97993 164250 98059 164253
rect 98126 164250 98132 164252
rect 97993 164248 98132 164250
rect 97993 164192 97998 164248
rect 98054 164192 98132 164248
rect 97993 164190 98132 164192
rect 97993 164187 98059 164190
rect 98126 164188 98132 164190
rect 98196 164188 98202 164252
rect 100017 164250 100083 164253
rect 101806 164250 101812 164252
rect 100017 164248 101812 164250
rect 100017 164192 100022 164248
rect 100078 164192 101812 164248
rect 100017 164190 101812 164192
rect 100017 164187 100083 164190
rect 101806 164188 101812 164190
rect 101876 164188 101882 164252
rect 102133 164250 102199 164253
rect 102726 164250 102732 164252
rect 102133 164248 102732 164250
rect 102133 164192 102138 164248
rect 102194 164192 102732 164248
rect 102133 164190 102732 164192
rect 102133 164187 102199 164190
rect 102726 164188 102732 164190
rect 102796 164188 102802 164252
rect 103513 164250 103579 164253
rect 103830 164250 103836 164252
rect 103513 164248 103836 164250
rect 103513 164192 103518 164248
rect 103574 164192 103836 164248
rect 103513 164190 103836 164192
rect 103513 164187 103579 164190
rect 103830 164188 103836 164190
rect 103900 164188 103906 164252
rect 105302 164188 105308 164252
rect 105372 164250 105378 164252
rect 106181 164250 106247 164253
rect 105372 164248 106247 164250
rect 105372 164192 106186 164248
rect 106242 164192 106247 164248
rect 105372 164190 106247 164192
rect 105372 164188 105378 164190
rect 106181 164187 106247 164190
rect 106365 164252 106431 164253
rect 106365 164248 106412 164252
rect 106476 164250 106482 164252
rect 236085 164250 236151 164253
rect 237046 164250 237052 164252
rect 106365 164192 106370 164248
rect 106365 164188 106412 164192
rect 106476 164190 106522 164250
rect 236085 164248 237052 164250
rect 236085 164192 236090 164248
rect 236146 164192 237052 164248
rect 236085 164190 237052 164192
rect 106476 164188 106482 164190
rect 106365 164187 106431 164188
rect 236085 164187 236151 164190
rect 237046 164188 237052 164190
rect 237116 164188 237122 164252
rect 237373 164250 237439 164253
rect 238150 164250 238156 164252
rect 237373 164248 238156 164250
rect 237373 164192 237378 164248
rect 237434 164192 238156 164248
rect 237373 164190 238156 164192
rect 237373 164187 237439 164190
rect 238150 164188 238156 164190
rect 238220 164188 238226 164252
rect 240133 164250 240199 164253
rect 240542 164250 240548 164252
rect 240133 164248 240548 164250
rect 240133 164192 240138 164248
rect 240194 164192 240548 164248
rect 240133 164190 240548 164192
rect 240133 164187 240199 164190
rect 240542 164188 240548 164190
rect 240612 164188 240618 164252
rect 241513 164250 241579 164253
rect 241646 164250 241652 164252
rect 241513 164248 241652 164250
rect 241513 164192 241518 164248
rect 241574 164192 241652 164248
rect 241513 164190 241652 164192
rect 241513 164187 241579 164190
rect 241646 164188 241652 164190
rect 241716 164188 241722 164252
rect 244273 164250 244339 164253
rect 245326 164250 245332 164252
rect 244273 164248 245332 164250
rect 244273 164192 244278 164248
rect 244334 164192 245332 164248
rect 244273 164190 245332 164192
rect 244273 164187 244339 164190
rect 245326 164188 245332 164190
rect 245396 164188 245402 164252
rect 245653 164250 245719 164253
rect 246430 164250 246436 164252
rect 245653 164248 246436 164250
rect 245653 164192 245658 164248
rect 245714 164192 246436 164248
rect 245653 164190 246436 164192
rect 245653 164187 245719 164190
rect 246430 164188 246436 164190
rect 246500 164188 246506 164252
rect 248413 164250 248479 164253
rect 248638 164250 248644 164252
rect 248413 164248 248644 164250
rect 248413 164192 248418 164248
rect 248474 164192 248644 164248
rect 248413 164190 248644 164192
rect 248413 164187 248479 164190
rect 248638 164188 248644 164190
rect 248708 164188 248714 164252
rect 249793 164250 249859 164253
rect 251173 164252 251239 164253
rect 250110 164250 250116 164252
rect 249793 164248 250116 164250
rect 249793 164192 249798 164248
rect 249854 164192 250116 164248
rect 249793 164190 250116 164192
rect 249793 164187 249859 164190
rect 250110 164188 250116 164190
rect 250180 164188 250186 164252
rect 251173 164250 251220 164252
rect 251128 164248 251220 164250
rect 251128 164192 251178 164248
rect 251128 164190 251220 164192
rect 251173 164188 251220 164190
rect 251284 164188 251290 164252
rect 252553 164250 252619 164253
rect 253422 164250 253428 164252
rect 252553 164248 253428 164250
rect 252553 164192 252558 164248
rect 252614 164192 253428 164248
rect 252553 164190 253428 164192
rect 251173 164187 251239 164188
rect 252553 164187 252619 164190
rect 253422 164188 253428 164190
rect 253492 164188 253498 164252
rect 253933 164250 253999 164253
rect 254526 164250 254532 164252
rect 253933 164248 254532 164250
rect 253933 164192 253938 164248
rect 253994 164192 254532 164248
rect 253933 164190 254532 164192
rect 253933 164187 253999 164190
rect 254526 164188 254532 164190
rect 254596 164188 254602 164252
rect 255313 164250 255379 164253
rect 255814 164250 255820 164252
rect 255313 164248 255820 164250
rect 255313 164192 255318 164248
rect 255374 164192 255820 164248
rect 255313 164190 255820 164192
rect 255313 164187 255379 164190
rect 255814 164188 255820 164190
rect 255884 164188 255890 164252
rect 256693 164250 256759 164253
rect 256918 164250 256924 164252
rect 256693 164248 256924 164250
rect 256693 164192 256698 164248
rect 256754 164192 256924 164248
rect 256693 164190 256924 164192
rect 256693 164187 256759 164190
rect 256918 164188 256924 164190
rect 256988 164188 256994 164252
rect 258073 164250 258139 164253
rect 259453 164252 259519 164253
rect 258390 164250 258396 164252
rect 258073 164248 258396 164250
rect 258073 164192 258078 164248
rect 258134 164192 258396 164248
rect 258073 164190 258396 164192
rect 258073 164187 258139 164190
rect 258390 164188 258396 164190
rect 258460 164188 258466 164252
rect 259453 164250 259500 164252
rect 259408 164248 259500 164250
rect 259408 164192 259458 164248
rect 259408 164190 259500 164192
rect 259453 164188 259500 164190
rect 259564 164188 259570 164252
rect 262806 164188 262812 164252
rect 262876 164250 262882 164252
rect 263501 164250 263567 164253
rect 262876 164248 263567 164250
rect 262876 164192 263506 164248
rect 263562 164192 263567 164248
rect 262876 164190 263567 164192
rect 262876 164188 262882 164190
rect 259453 164187 259519 164188
rect 263501 164187 263567 164190
rect 263777 164250 263843 164253
rect 263910 164250 263916 164252
rect 263777 164248 263916 164250
rect 263777 164192 263782 164248
rect 263838 164192 263916 164248
rect 263777 164190 263916 164192
rect 263777 164187 263843 164190
rect 263910 164188 263916 164190
rect 263980 164188 263986 164252
rect 267825 164250 267891 164253
rect 268694 164250 268700 164252
rect 267825 164248 268700 164250
rect 267825 164192 267830 164248
rect 267886 164192 268700 164248
rect 267825 164190 268700 164192
rect 267825 164187 267891 164190
rect 268694 164188 268700 164190
rect 268764 164188 268770 164252
rect 269113 164250 269179 164253
rect 269798 164250 269804 164252
rect 269113 164248 269804 164250
rect 269113 164192 269118 164248
rect 269174 164192 269804 164248
rect 269113 164190 269804 164192
rect 269113 164187 269179 164190
rect 269798 164188 269804 164190
rect 269868 164188 269874 164252
rect 270493 164250 270559 164253
rect 271270 164250 271276 164252
rect 270493 164248 271276 164250
rect 270493 164192 270498 164248
rect 270554 164192 271276 164248
rect 270493 164190 271276 164192
rect 270493 164187 270559 164190
rect 271270 164188 271276 164190
rect 271340 164188 271346 164252
rect 274398 164188 274404 164252
rect 274468 164250 274474 164252
rect 274541 164250 274607 164253
rect 274468 164248 274607 164250
rect 274468 164192 274546 164248
rect 274602 164192 274607 164248
rect 274468 164190 274607 164192
rect 274468 164188 274474 164190
rect 274541 164187 274607 164190
rect 276013 164250 276079 164253
rect 276974 164250 276980 164252
rect 276013 164248 276980 164250
rect 276013 164192 276018 164248
rect 276074 164192 276980 164248
rect 276013 164190 276980 164192
rect 276013 164187 276079 164190
rect 276974 164188 276980 164190
rect 277044 164188 277050 164252
rect 277393 164250 277459 164253
rect 396073 164252 396139 164253
rect 278078 164250 278084 164252
rect 277393 164248 278084 164250
rect 277393 164192 277398 164248
rect 277454 164192 278084 164248
rect 277393 164190 278084 164192
rect 277393 164187 277459 164190
rect 278078 164188 278084 164190
rect 278148 164188 278154 164252
rect 318374 164250 318380 164252
rect 315990 164190 318380 164250
rect 57646 164052 57652 164116
rect 57716 164114 57722 164116
rect 58157 164114 58223 164117
rect 57716 164112 58223 164114
rect 57716 164056 58162 164112
rect 58218 164056 58223 164112
rect 57716 164054 58223 164056
rect 57716 164052 57722 164054
rect 58157 164051 58223 164054
rect 206318 164052 206324 164116
rect 206388 164114 206394 164116
rect 315990 164114 316050 164190
rect 318374 164188 318380 164190
rect 318444 164188 318450 164252
rect 396022 164250 396028 164252
rect 395982 164190 396028 164250
rect 396092 164248 396139 164252
rect 396134 164192 396139 164248
rect 396022 164188 396028 164190
rect 396092 164188 396139 164192
rect 396073 164187 396139 164188
rect 398833 164250 398899 164253
rect 399518 164250 399524 164252
rect 398833 164248 399524 164250
rect 398833 164192 398838 164248
rect 398894 164192 399524 164248
rect 398833 164190 399524 164192
rect 398833 164187 398899 164190
rect 399518 164188 399524 164190
rect 399588 164188 399594 164252
rect 400213 164250 400279 164253
rect 403065 164252 403131 164253
rect 400438 164250 400444 164252
rect 400213 164248 400444 164250
rect 400213 164192 400218 164248
rect 400274 164192 400444 164248
rect 400213 164190 400444 164192
rect 400213 164187 400279 164190
rect 400438 164188 400444 164190
rect 400508 164188 400514 164252
rect 403014 164188 403020 164252
rect 403084 164250 403131 164252
rect 405733 164250 405799 164253
rect 406510 164250 406516 164252
rect 403084 164248 403176 164250
rect 403126 164192 403176 164248
rect 403084 164190 403176 164192
rect 405733 164248 406516 164250
rect 405733 164192 405738 164248
rect 405794 164192 406516 164248
rect 405733 164190 406516 164192
rect 403084 164188 403131 164190
rect 403065 164187 403131 164188
rect 405733 164187 405799 164190
rect 406510 164188 406516 164190
rect 406580 164188 406586 164252
rect 407205 164250 407271 164253
rect 407614 164250 407620 164252
rect 407205 164248 407620 164250
rect 407205 164192 407210 164248
rect 407266 164192 407620 164248
rect 407205 164190 407620 164192
rect 407205 164187 407271 164190
rect 407614 164188 407620 164190
rect 407684 164188 407690 164252
rect 408493 164250 408559 164253
rect 408718 164250 408724 164252
rect 408493 164248 408724 164250
rect 408493 164192 408498 164248
rect 408554 164192 408724 164248
rect 408493 164190 408724 164192
rect 408493 164187 408559 164190
rect 408718 164188 408724 164190
rect 408788 164188 408794 164252
rect 409873 164250 409939 164253
rect 411345 164252 411411 164253
rect 410006 164250 410012 164252
rect 409873 164248 410012 164250
rect 409873 164192 409878 164248
rect 409934 164192 410012 164248
rect 409873 164190 410012 164192
rect 409873 164187 409939 164190
rect 410006 164188 410012 164190
rect 410076 164188 410082 164252
rect 411294 164250 411300 164252
rect 411254 164190 411300 164250
rect 411364 164248 411411 164252
rect 411406 164192 411411 164248
rect 411294 164188 411300 164190
rect 411364 164188 411411 164192
rect 411345 164187 411411 164188
rect 412725 164250 412791 164253
rect 413318 164250 413324 164252
rect 412725 164248 413324 164250
rect 412725 164192 412730 164248
rect 412786 164192 413324 164248
rect 412725 164190 413324 164192
rect 412725 164187 412791 164190
rect 413318 164188 413324 164190
rect 413388 164188 413394 164252
rect 414013 164250 414079 164253
rect 414422 164250 414428 164252
rect 414013 164248 414428 164250
rect 414013 164192 414018 164248
rect 414074 164192 414428 164248
rect 414013 164190 414428 164192
rect 414013 164187 414079 164190
rect 414422 164188 414428 164190
rect 414492 164188 414498 164252
rect 416773 164250 416839 164253
rect 416998 164250 417004 164252
rect 416773 164248 417004 164250
rect 416773 164192 416778 164248
rect 416834 164192 417004 164248
rect 416773 164190 417004 164192
rect 416773 164187 416839 164190
rect 416998 164188 417004 164190
rect 417068 164188 417074 164252
rect 418153 164250 418219 164253
rect 418286 164250 418292 164252
rect 418153 164248 418292 164250
rect 418153 164192 418158 164248
rect 418214 164192 418292 164248
rect 418153 164190 418292 164192
rect 418153 164187 418219 164190
rect 418286 164188 418292 164190
rect 418356 164188 418362 164252
rect 419533 164250 419599 164253
rect 420678 164250 420684 164252
rect 419533 164248 420684 164250
rect 419533 164192 419538 164248
rect 419594 164192 420684 164248
rect 419533 164190 420684 164192
rect 419533 164187 419599 164190
rect 420678 164188 420684 164190
rect 420748 164188 420754 164252
rect 422886 164188 422892 164252
rect 422956 164250 422962 164252
rect 423581 164250 423647 164253
rect 422956 164248 423647 164250
rect 422956 164192 423586 164248
rect 423642 164192 423647 164248
rect 422956 164190 423647 164192
rect 422956 164188 422962 164190
rect 423581 164187 423647 164190
rect 425278 164188 425284 164252
rect 425348 164250 425354 164252
rect 426341 164250 426407 164253
rect 427721 164252 427787 164253
rect 427670 164250 427676 164252
rect 425348 164248 426407 164250
rect 425348 164192 426346 164248
rect 426402 164192 426407 164248
rect 425348 164190 426407 164192
rect 427630 164190 427676 164250
rect 427740 164248 427787 164252
rect 427782 164192 427787 164248
rect 425348 164188 425354 164190
rect 426341 164187 426407 164190
rect 427670 164188 427676 164190
rect 427740 164188 427787 164192
rect 428774 164188 428780 164252
rect 428844 164250 428850 164252
rect 429101 164250 429167 164253
rect 428844 164248 429167 164250
rect 428844 164192 429106 164248
rect 429162 164192 429167 164248
rect 428844 164190 429167 164192
rect 428844 164188 428850 164190
rect 427721 164187 427787 164188
rect 429101 164187 429167 164190
rect 430573 164250 430639 164253
rect 430982 164250 430988 164252
rect 430573 164248 430988 164250
rect 430573 164192 430578 164248
rect 430634 164192 430988 164248
rect 430573 164190 430988 164192
rect 430573 164187 430639 164190
rect 430982 164188 430988 164190
rect 431052 164188 431058 164252
rect 431953 164250 432019 164253
rect 432270 164250 432276 164252
rect 431953 164248 432276 164250
rect 431953 164192 431958 164248
rect 432014 164192 432276 164248
rect 431953 164190 432276 164192
rect 431953 164187 432019 164190
rect 432270 164188 432276 164190
rect 432340 164188 432346 164252
rect 433374 164188 433380 164252
rect 433444 164250 433450 164252
rect 434621 164250 434687 164253
rect 433444 164248 434687 164250
rect 433444 164192 434626 164248
rect 434682 164192 434687 164248
rect 433444 164190 434687 164192
rect 433444 164188 433450 164190
rect 434621 164187 434687 164190
rect 434805 164250 434871 164253
rect 435766 164250 435772 164252
rect 434805 164248 435772 164250
rect 434805 164192 434810 164248
rect 434866 164192 435772 164248
rect 434805 164190 435772 164192
rect 434805 164187 434871 164190
rect 435766 164188 435772 164190
rect 435836 164188 435842 164252
rect 206388 164054 316050 164114
rect 375557 164114 375623 164117
rect 376886 164114 376892 164116
rect 375557 164112 376892 164114
rect 375557 164056 375562 164112
rect 375618 164056 376892 164112
rect 375557 164054 376892 164056
rect 206388 164052 206394 164054
rect 375557 164051 375623 164054
rect 376886 164052 376892 164054
rect 376956 164052 376962 164116
rect -960 162740 480 162980
rect 217174 162692 217180 162756
rect 217244 162754 217250 162756
rect 217961 162754 218027 162757
rect 217244 162752 218027 162754
rect 217244 162696 217966 162752
rect 218022 162696 218027 162752
rect 217244 162694 218027 162696
rect 217244 162692 217250 162694
rect 217961 162691 218027 162694
rect 376886 162692 376892 162756
rect 376956 162754 376962 162756
rect 437749 162754 437815 162757
rect 376956 162752 437815 162754
rect 376956 162696 437754 162752
rect 437810 162696 437815 162752
rect 376956 162694 437815 162696
rect 376956 162692 376962 162694
rect 437749 162691 437815 162694
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 363454 149154 363460 149156
rect 246 149094 363460 149154
rect 363454 149092 363460 149094
rect 363524 149092 363530 149156
rect 57646 147732 57652 147796
rect 57716 147794 57722 147796
rect 58065 147794 58131 147797
rect 57716 147792 58131 147794
rect 57716 147736 58070 147792
rect 58126 147736 58131 147792
rect 57716 147734 58131 147736
rect 57716 147732 57722 147734
rect 58065 147731 58131 147734
rect 377438 147732 377444 147796
rect 377508 147794 377514 147796
rect 379053 147794 379119 147797
rect 377508 147792 379119 147794
rect 377508 147736 379058 147792
rect 379114 147736 379119 147792
rect 377508 147734 379119 147736
rect 377508 147732 377514 147734
rect 379053 147731 379119 147734
rect 54201 146298 54267 146301
rect 54753 146298 54819 146301
rect 100017 146298 100083 146301
rect 54201 146296 100083 146298
rect 54201 146240 54206 146296
rect 54262 146240 54758 146296
rect 54814 146240 100022 146296
rect 100078 146240 100083 146296
rect 54201 146238 100083 146240
rect 54201 146235 54267 146238
rect 54753 146235 54819 146238
rect 100017 146235 100083 146238
rect 217317 146298 217383 146301
rect 217542 146298 217548 146300
rect 217317 146296 217548 146298
rect 217317 146240 217322 146296
rect 217378 146240 217548 146296
rect 217317 146238 217548 146240
rect 217317 146235 217383 146238
rect 217542 146236 217548 146238
rect 217612 146236 217618 146300
rect 218237 146298 218303 146301
rect 219893 146298 219959 146301
rect 267733 146298 267799 146301
rect 218237 146296 267799 146298
rect 218237 146240 218242 146296
rect 218298 146240 219898 146296
rect 219954 146240 267738 146296
rect 267794 146240 267799 146296
rect 218237 146238 267799 146240
rect 218237 146235 218303 146238
rect 219893 146235 219959 146238
rect 267733 146235 267799 146238
rect 377990 146236 377996 146300
rect 378060 146298 378066 146300
rect 378869 146298 378935 146301
rect 378060 146296 378935 146298
rect 378060 146240 378874 146296
rect 378930 146240 378935 146296
rect 378060 146238 378935 146240
rect 378060 146236 378066 146238
rect 378869 146235 378935 146238
rect 56133 146162 56199 146165
rect 59721 146162 59787 146165
rect 99373 146162 99439 146165
rect 56133 146160 99439 146162
rect 56133 146104 56138 146160
rect 56194 146104 59726 146160
rect 59782 146104 99378 146160
rect 99434 146104 99439 146160
rect 56133 146102 99439 146104
rect 56133 146099 56199 146102
rect 59721 146099 59787 146102
rect 99373 146099 99439 146102
rect 219893 146162 219959 146165
rect 220813 146162 220879 146165
rect 267825 146162 267891 146165
rect 219893 146160 267891 146162
rect 219893 146104 219898 146160
rect 219954 146104 220818 146160
rect 220874 146104 267830 146160
rect 267886 146104 267891 146160
rect 219893 146102 267891 146104
rect 219893 146099 219959 146102
rect 220813 146099 220879 146102
rect 267825 146099 267891 146102
rect 215845 146026 215911 146029
rect 219433 146026 219499 146029
rect 263593 146026 263659 146029
rect 215845 146024 263659 146026
rect 215845 145968 215850 146024
rect 215906 145968 219438 146024
rect 219494 145968 263598 146024
rect 263654 145968 263659 146024
rect 215845 145966 263659 145968
rect 215845 145963 215911 145966
rect 219433 145963 219499 145966
rect 263593 145963 263659 145966
rect 378869 146026 378935 146029
rect 415485 146026 415551 146029
rect 378869 146024 415551 146026
rect 378869 145968 378874 146024
rect 378930 145968 415490 146024
rect 415546 145968 415551 146024
rect 378869 145966 415551 145968
rect 378869 145963 378935 145966
rect 415485 145963 415551 145966
rect 369761 145890 369827 145893
rect 377622 145890 377628 145892
rect 369761 145888 377628 145890
rect 369761 145832 369766 145888
rect 369822 145832 377628 145888
rect 369761 145830 377628 145832
rect 369761 145827 369827 145830
rect 377622 145828 377628 145830
rect 377692 145890 377698 145892
rect 423673 145890 423739 145893
rect 377692 145888 423739 145890
rect 377692 145832 423678 145888
rect 423734 145832 423739 145888
rect 377692 145830 423739 145832
rect 377692 145828 377698 145830
rect 423673 145827 423739 145830
rect 58709 145754 58775 145757
rect 92473 145754 92539 145757
rect 58709 145752 92539 145754
rect 58709 145696 58714 145752
rect 58770 145696 92478 145752
rect 92534 145696 92539 145752
rect 58709 145694 92539 145696
rect 58709 145691 58775 145694
rect 92473 145691 92539 145694
rect 213269 145754 213335 145757
rect 237373 145754 237439 145757
rect 213269 145752 237439 145754
rect 213269 145696 213274 145752
rect 213330 145696 237378 145752
rect 237434 145696 237439 145752
rect 213269 145694 237439 145696
rect 213269 145691 213335 145694
rect 237373 145691 237439 145694
rect 371049 145754 371115 145757
rect 377489 145754 377555 145757
rect 423765 145754 423831 145757
rect 371049 145752 423831 145754
rect 371049 145696 371054 145752
rect 371110 145696 377494 145752
rect 377550 145696 423770 145752
rect 423826 145696 423831 145752
rect 371049 145694 423831 145696
rect 371049 145691 371115 145694
rect 377489 145691 377555 145694
rect 423765 145691 423831 145694
rect 58893 145618 58959 145621
rect 98637 145618 98703 145621
rect 58893 145616 98703 145618
rect 58893 145560 58898 145616
rect 58954 145560 98642 145616
rect 98698 145560 98703 145616
rect 58893 145558 98703 145560
rect 58893 145555 58959 145558
rect 98637 145555 98703 145558
rect 214465 145618 214531 145621
rect 269113 145618 269179 145621
rect 214465 145616 269179 145618
rect 214465 145560 214470 145616
rect 214526 145560 269118 145616
rect 269174 145560 269179 145616
rect 214465 145558 269179 145560
rect 214465 145555 214531 145558
rect 269113 145555 269179 145558
rect 371693 145618 371759 145621
rect 377806 145618 377812 145620
rect 371693 145616 377812 145618
rect 371693 145560 371698 145616
rect 371754 145560 377812 145616
rect 371693 145558 377812 145560
rect 371693 145555 371759 145558
rect 377806 145556 377812 145558
rect 377876 145618 377882 145620
rect 426433 145618 426499 145621
rect 377876 145616 426499 145618
rect 377876 145560 426438 145616
rect 426494 145560 426499 145616
rect 377876 145558 426499 145560
rect 377876 145556 377882 145558
rect 426433 145555 426499 145558
rect 510613 145482 510679 145485
rect 510838 145482 510844 145484
rect 510613 145480 510844 145482
rect 510613 145424 510618 145480
rect 510674 145424 510844 145480
rect 510613 145422 510844 145424
rect 510613 145419 510679 145422
rect 510838 145420 510844 145422
rect 510908 145420 510914 145484
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 190862 144876 190868 144940
rect 190932 144938 190938 144940
rect 191281 144938 191347 144941
rect 338481 144940 338547 144941
rect 338430 144938 338436 144940
rect 190932 144936 191347 144938
rect 190932 144880 191286 144936
rect 191342 144880 191347 144936
rect 190932 144878 191347 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 190932 144876 190938 144878
rect 179689 144875 179755 144876
rect 191281 144875 191347 144878
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144940
rect 499868 144938 499874 144940
rect 500217 144938 500283 144941
rect 499868 144936 500283 144938
rect 499868 144880 500222 144936
rect 500278 144880 500283 144936
rect 499868 144878 500283 144880
rect 499868 144876 499874 144878
rect 500217 144875 500283 144878
rect 57462 140796 57468 140860
rect 57532 140858 57538 140860
rect 59353 140858 59419 140861
rect 57532 140856 59419 140858
rect 57532 140800 59358 140856
rect 59414 140800 59419 140856
rect 57532 140798 59419 140800
rect 57532 140796 57538 140798
rect 59353 140795 59419 140798
rect 358905 139362 358971 139365
rect 519261 139362 519327 139365
rect 356562 139360 358971 139362
rect 356562 139304 358910 139360
rect 358966 139304 358971 139360
rect 356562 139302 358971 139304
rect 198825 139226 198891 139229
rect 197126 139224 198891 139226
rect 197126 139220 198830 139224
rect 196604 139168 198830 139220
rect 198886 139168 198891 139224
rect 356562 139190 356622 139302
rect 358905 139299 358971 139302
rect 516558 139360 519327 139362
rect 516558 139304 519266 139360
rect 519322 139304 519327 139360
rect 516558 139302 519327 139304
rect 516558 139190 516618 139302
rect 519261 139299 519327 139302
rect 583520 139212 584960 139452
rect 196604 139166 198891 139168
rect 196604 139160 197186 139166
rect 198825 139163 198891 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 57237 97474 57303 97477
rect 57237 97472 60062 97474
rect 57237 97416 57242 97472
rect 57298 97416 60062 97472
rect 57237 97414 60062 97416
rect 57237 97411 57303 97414
rect 60002 96894 60062 97414
rect 217409 96930 217475 96933
rect 377213 96930 377279 96933
rect 217409 96928 219450 96930
rect 217409 96872 217414 96928
rect 217470 96924 219450 96928
rect 377213 96928 379530 96930
rect 217470 96872 220064 96924
rect 217409 96870 220064 96872
rect 217409 96867 217475 96870
rect 219390 96864 220064 96870
rect 377213 96872 377218 96928
rect 377274 96924 379530 96928
rect 377274 96872 380052 96924
rect 377213 96870 380052 96872
rect 377213 96867 377279 96870
rect 379470 96864 380052 96870
rect 57513 96522 57579 96525
rect 57513 96520 60062 96522
rect 57513 96464 57518 96520
rect 57574 96464 60062 96520
rect 57513 96462 60062 96464
rect 57513 96459 57579 96462
rect 60002 95942 60062 96462
rect 217869 95978 217935 95981
rect 377029 95978 377095 95981
rect 217869 95976 219450 95978
rect 217869 95920 217874 95976
rect 217930 95972 219450 95976
rect 377029 95976 379530 95978
rect 217930 95920 220064 95972
rect 217869 95918 220064 95920
rect 217869 95915 217935 95918
rect 219390 95912 220064 95918
rect 377029 95920 377034 95976
rect 377090 95972 379530 95976
rect 377090 95920 380052 95972
rect 377029 95918 380052 95920
rect 377029 95915 377095 95918
rect 379470 95912 380052 95918
rect 57605 93802 57671 93805
rect 217593 93802 217659 93805
rect 377581 93802 377647 93805
rect 57605 93800 60062 93802
rect 57605 93744 57610 93800
rect 57666 93744 60062 93800
rect 57605 93742 60062 93744
rect 217593 93800 219450 93802
rect 217593 93744 217598 93800
rect 217654 93796 219450 93800
rect 377581 93800 379530 93802
rect 217654 93744 220064 93796
rect 217593 93742 220064 93744
rect 57605 93739 57671 93742
rect 217593 93739 217659 93742
rect 219390 93736 220064 93742
rect 377581 93744 377586 93800
rect 377642 93796 379530 93800
rect 377642 93744 380052 93796
rect 377581 93742 380052 93744
rect 377581 93739 377647 93742
rect 379470 93736 380052 93742
rect 57421 93394 57487 93397
rect 57421 93392 60062 93394
rect 57421 93336 57426 93392
rect 57482 93336 60062 93392
rect 57421 93334 60062 93336
rect 57421 93331 57487 93334
rect 60002 92814 60062 93334
rect 216857 92850 216923 92853
rect 376937 92850 377003 92853
rect 216857 92848 219450 92850
rect 216857 92792 216862 92848
rect 216918 92844 219450 92848
rect 376937 92848 379530 92850
rect 216918 92792 220064 92844
rect 216857 92790 220064 92792
rect 216857 92787 216923 92790
rect 219390 92784 220064 92790
rect 376937 92792 376942 92848
rect 376998 92844 379530 92848
rect 376998 92792 380052 92844
rect 376937 92790 380052 92792
rect 376937 92787 377003 92790
rect 379470 92784 380052 92790
rect 57697 91082 57763 91085
rect 217777 91082 217843 91085
rect 377673 91082 377739 91085
rect 57697 91080 60062 91082
rect 57697 91024 57702 91080
rect 57758 91024 60062 91080
rect 57697 91022 60062 91024
rect 217777 91080 219450 91082
rect 217777 91024 217782 91080
rect 217838 91076 219450 91080
rect 377673 91080 379530 91082
rect 217838 91024 220064 91076
rect 217777 91022 220064 91024
rect 57697 91019 57763 91022
rect 217777 91019 217843 91022
rect 219390 91016 220064 91022
rect 377673 91024 377678 91080
rect 377734 91076 379530 91080
rect 377734 91024 380052 91076
rect 377673 91022 380052 91024
rect 377673 91019 377739 91022
rect 379470 91016 380052 91022
rect 57329 90538 57395 90541
rect 57329 90536 60062 90538
rect 57329 90480 57334 90536
rect 57390 90480 60062 90536
rect 57329 90478 60062 90480
rect 57329 90475 57395 90478
rect 60002 89958 60062 90478
rect 217501 89994 217567 89997
rect 377857 89994 377923 89997
rect 217501 89992 219450 89994
rect 217501 89936 217506 89992
rect 217562 89988 219450 89992
rect 377857 89992 379530 89994
rect 217562 89936 220064 89988
rect 217501 89934 220064 89936
rect 217501 89931 217567 89934
rect 219390 89928 220064 89934
rect 377857 89936 377862 89992
rect 377918 89988 379530 89992
rect 377918 89936 380052 89988
rect 377857 89934 380052 89936
rect 377857 89931 377923 89934
rect 379470 89928 380052 89934
rect 57789 88226 57855 88229
rect 217685 88226 217751 88229
rect 377765 88226 377831 88229
rect 57789 88224 60062 88226
rect 57789 88168 57794 88224
rect 57850 88168 60062 88224
rect 57789 88166 60062 88168
rect 217685 88224 219450 88226
rect 217685 88168 217690 88224
rect 217746 88220 219450 88224
rect 377765 88224 379530 88226
rect 217746 88168 220064 88220
rect 217685 88166 220064 88168
rect 57789 88163 57855 88166
rect 217685 88163 217751 88166
rect 219390 88160 220064 88166
rect 377765 88168 377770 88224
rect 377826 88220 379530 88224
rect 377826 88168 380052 88220
rect 377765 88166 380052 88168
rect 377765 88163 377831 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 358813 79930 358879 79933
rect 518893 79930 518959 79933
rect 520181 79930 520247 79933
rect 356562 79928 358879 79930
rect 356562 79872 358818 79928
rect 358874 79872 358879 79928
rect 356562 79870 358879 79872
rect 199285 79386 199351 79389
rect 197126 79384 199351 79386
rect 197126 79380 199290 79384
rect 196604 79328 199290 79380
rect 199346 79328 199351 79384
rect 356562 79350 356622 79870
rect 358813 79867 358879 79870
rect 516558 79928 520247 79930
rect 516558 79872 518898 79928
rect 518954 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 518893 79867 518959 79870
rect 520181 79867 520247 79870
rect 196604 79326 199351 79328
rect 196604 79320 197186 79326
rect 199285 79323 199351 79326
rect 359089 78298 359155 78301
rect 519077 78298 519143 78301
rect 356562 78296 359155 78298
rect 356562 78240 359094 78296
rect 359150 78240 359155 78296
rect 356562 78238 359155 78240
rect 198917 77754 198983 77757
rect 197126 77752 198983 77754
rect 197126 77748 198922 77752
rect 196604 77696 198922 77748
rect 198978 77696 198983 77752
rect 356562 77718 356622 78238
rect 359089 78235 359155 78238
rect 516558 78296 519143 78298
rect 516558 78240 519082 78296
rect 519138 78240 519143 78296
rect 516558 78238 519143 78240
rect 516558 77718 516618 78238
rect 519077 78235 519143 78238
rect 196604 77694 198983 77696
rect 196604 77688 197186 77694
rect 198917 77691 198983 77694
rect 359365 76938 359431 76941
rect 356562 76936 359431 76938
rect 356562 76880 359370 76936
rect 359426 76880 359431 76936
rect 356562 76878 359431 76880
rect 199009 76394 199075 76397
rect 197126 76392 199075 76394
rect 197126 76388 199014 76392
rect 196604 76336 199014 76388
rect 199070 76336 199075 76392
rect 356562 76358 356622 76878
rect 359365 76875 359431 76878
rect 519445 76802 519511 76805
rect 516558 76800 519511 76802
rect 516558 76744 519450 76800
rect 519506 76744 519511 76800
rect 516558 76742 519511 76744
rect 516558 76358 516618 76742
rect 519445 76739 519511 76742
rect 196604 76334 199075 76336
rect 196604 76328 197186 76334
rect 199009 76331 199075 76334
rect 359273 75442 359339 75445
rect 519353 75442 519419 75445
rect 356562 75440 359339 75442
rect 356562 75384 359278 75440
rect 359334 75384 359339 75440
rect 356562 75382 359339 75384
rect 198733 74898 198799 74901
rect 197126 74896 198799 74898
rect 197126 74892 198738 74896
rect 196604 74840 198738 74892
rect 198794 74840 198799 74896
rect 356562 74862 356622 75382
rect 359273 75379 359339 75382
rect 516558 75440 519419 75442
rect 516558 75384 519358 75440
rect 519414 75384 519419 75440
rect 516558 75382 519419 75384
rect 516558 74862 516618 75382
rect 519353 75379 519419 75382
rect 196604 74838 198799 74840
rect 196604 74832 197186 74838
rect 198733 74835 198799 74838
rect 518985 74218 519051 74221
rect 516558 74216 519051 74218
rect 516558 74160 518990 74216
rect 519046 74160 519051 74216
rect 516558 74158 519051 74160
rect 359181 74082 359247 74085
rect 356562 74080 359247 74082
rect 356562 74024 359186 74080
rect 359242 74024 359247 74080
rect 356562 74022 359247 74024
rect 199193 73674 199259 73677
rect 197126 73672 199259 73674
rect 197126 73668 199198 73672
rect 196604 73616 199198 73668
rect 199254 73616 199259 73672
rect 356562 73638 356622 74022
rect 359181 74019 359247 74022
rect 516558 73638 516618 74158
rect 518985 74155 519051 74158
rect 196604 73614 199259 73616
rect 196604 73608 197186 73614
rect 199193 73611 199259 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 57605 70138 57671 70141
rect 57605 70136 60062 70138
rect 57605 70080 57610 70136
rect 57666 70080 60062 70136
rect 57605 70078 60062 70080
rect 57605 70075 57671 70078
rect 60002 69966 60062 70078
rect 216673 70002 216739 70005
rect 376937 70002 377003 70005
rect 216673 70000 219450 70002
rect 216673 69944 216678 70000
rect 216734 69996 219450 70000
rect 376937 70000 379530 70002
rect 216734 69944 220064 69996
rect 216673 69942 220064 69944
rect 216673 69939 216739 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 375414 68852 375420 68916
rect 375484 68914 375490 68916
rect 376661 68914 376727 68917
rect 375484 68912 376727 68914
rect 375484 68856 376666 68912
rect 376722 68856 376727 68912
rect 375484 68854 376727 68856
rect 375484 68852 375490 68854
rect 376661 68851 376727 68854
rect 216673 68370 216739 68373
rect 217961 68370 218027 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68312 217966 68368
rect 218022 68364 219450 68368
rect 376937 68368 379530 68370
rect 218022 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 217961 68307 218027 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 46790 67764 46796 67828
rect 46860 67826 46866 67828
rect 60002 67826 60062 68062
rect 214598 68036 214604 68100
rect 214668 68098 214674 68100
rect 376017 68098 376083 68101
rect 214668 68092 219450 68098
rect 376017 68096 379530 68098
rect 214668 68038 220064 68092
rect 214668 68036 214674 68038
rect 219390 68032 220064 68038
rect 376017 68040 376022 68096
rect 376078 68092 379530 68096
rect 376078 68040 380052 68092
rect 376017 68038 380052 68040
rect 376017 68035 376083 68038
rect 379470 68032 380052 68038
rect 46860 67766 60062 67826
rect 46860 67764 46866 67766
rect 218697 60620 218763 60621
rect 219249 60620 219315 60621
rect 218646 60618 218652 60620
rect 218606 60558 218652 60618
rect 218716 60616 218763 60620
rect 219198 60618 219204 60620
rect 218758 60560 218763 60616
rect 218646 60556 218652 60558
rect 218716 60556 218763 60560
rect 219158 60558 219204 60618
rect 219268 60616 219315 60620
rect 219310 60560 219315 60616
rect 219198 60556 219204 60558
rect 219268 60556 219315 60560
rect 218697 60555 218763 60556
rect 219249 60555 219315 60556
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 94497 59804 94563 59805
rect 101765 59804 101831 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 94497 59800 94550 59804
rect 94614 59802 94620 59804
rect 101752 59802 101758 59804
rect 94497 59744 94502 59800
rect 83190 59740 83196 59742
rect 94497 59740 94550 59744
rect 94614 59742 94654 59802
rect 101674 59742 101758 59802
rect 101822 59800 101831 59804
rect 101826 59744 101831 59800
rect 94614 59740 94620 59742
rect 101752 59740 101758 59742
rect 101822 59740 101831 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 94497 59739 94563 59740
rect 101765 59739 101831 59740
rect 102777 59804 102843 59805
rect 113541 59804 113607 59805
rect 237097 59804 237163 59805
rect 255865 59804 255931 59805
rect 256969 59804 257035 59805
rect 262857 59804 262923 59805
rect 102777 59800 102846 59804
rect 102777 59744 102782 59800
rect 102838 59744 102846 59800
rect 102777 59740 102846 59744
rect 102910 59802 102916 59804
rect 102910 59742 102934 59802
rect 113541 59800 113590 59804
rect 113654 59802 113660 59804
rect 113541 59744 113546 59800
rect 102910 59740 102916 59742
rect 113541 59740 113590 59744
rect 113654 59742 113698 59802
rect 237097 59800 237142 59804
rect 237206 59802 237212 59804
rect 237097 59744 237102 59800
rect 113654 59740 113660 59742
rect 237097 59740 237142 59744
rect 237206 59742 237254 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 255865 59744 255870 59800
rect 237206 59740 237212 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 256969 59800 256998 59804
rect 257062 59802 257068 59804
rect 262840 59802 262846 59804
rect 256969 59744 256974 59800
rect 255974 59740 255980 59742
rect 256969 59740 256998 59744
rect 257062 59742 257126 59802
rect 262766 59742 262846 59802
rect 262910 59800 262923 59804
rect 262918 59744 262923 59800
rect 257062 59740 257068 59742
rect 262840 59740 262846 59742
rect 262910 59740 262923 59744
rect 102777 59739 102843 59740
rect 113541 59739 113607 59740
rect 237097 59739 237163 59740
rect 255865 59739 255931 59740
rect 256969 59739 257035 59740
rect 262857 59739 262923 59740
rect 263869 59804 263935 59805
rect 396073 59804 396139 59805
rect 263869 59800 263934 59804
rect 263869 59744 263874 59800
rect 263930 59744 263934 59800
rect 263869 59740 263934 59744
rect 263998 59802 264004 59804
rect 396048 59802 396054 59804
rect 263998 59742 264026 59802
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 263998 59740 264004 59742
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 263869 59739 263935 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 416957 59804 417023 59805
rect 423489 59804 423555 59805
rect 423949 59804 424015 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 416957 59800 416998 59804
rect 417062 59802 417068 59804
rect 416957 59744 416962 59800
rect 397206 59740 397212 59742
rect 416957 59740 416998 59744
rect 417062 59742 417114 59802
rect 423489 59800 423526 59804
rect 423590 59802 423596 59804
rect 423928 59802 423934 59804
rect 423489 59744 423494 59800
rect 417062 59740 417068 59742
rect 423489 59740 423526 59744
rect 423590 59742 423646 59802
rect 423858 59742 423934 59802
rect 423998 59800 424015 59804
rect 424010 59744 424015 59800
rect 423590 59740 423596 59742
rect 423928 59740 423934 59742
rect 423998 59740 424015 59744
rect 397085 59739 397151 59740
rect 416957 59739 417023 59740
rect 423489 59739 423555 59740
rect 423949 59739 424015 59740
rect 107561 59668 107627 59669
rect 258073 59668 258139 59669
rect 260649 59668 260715 59669
rect 261753 59668 261819 59669
rect 308489 59668 308555 59669
rect 315849 59668 315915 59669
rect 403065 59668 403131 59669
rect 404169 59668 404235 59669
rect 105288 59666 105294 59668
rect 84150 59606 105294 59666
rect 57646 59468 57652 59532
rect 57716 59530 57722 59532
rect 84150 59530 84210 59606
rect 105288 59604 105294 59606
rect 105358 59604 105364 59668
rect 105968 59604 105974 59668
rect 106038 59604 106044 59668
rect 107561 59664 107606 59668
rect 107670 59666 107676 59668
rect 107561 59608 107566 59664
rect 107561 59604 107606 59608
rect 107670 59606 107718 59666
rect 258073 59664 258086 59668
rect 258150 59666 258156 59668
rect 258073 59608 258078 59664
rect 107670 59604 107676 59606
rect 258073 59604 258086 59608
rect 258150 59606 258230 59666
rect 260649 59664 260670 59668
rect 260734 59666 260740 59668
rect 260649 59608 260654 59664
rect 258150 59604 258156 59606
rect 260649 59604 260670 59608
rect 260734 59606 260806 59666
rect 260734 59604 260740 59606
rect 261752 59604 261758 59668
rect 261822 59666 261828 59668
rect 261822 59606 261910 59666
rect 308489 59664 308542 59668
rect 308606 59666 308612 59668
rect 308489 59608 308494 59664
rect 261822 59604 261828 59606
rect 308489 59604 308542 59608
rect 308606 59606 308646 59666
rect 315849 59664 315886 59668
rect 315950 59666 315956 59668
rect 315849 59608 315854 59664
rect 308606 59604 308612 59606
rect 315849 59604 315886 59608
rect 315950 59606 316006 59666
rect 403065 59664 403126 59668
rect 403065 59608 403070 59664
rect 315950 59604 315956 59606
rect 403065 59604 403126 59608
rect 403190 59666 403196 59668
rect 403190 59606 403222 59666
rect 404169 59664 404214 59668
rect 404278 59666 404284 59668
rect 412541 59666 412607 59669
rect 416037 59668 416103 59669
rect 419441 59668 419507 59669
rect 421741 59668 421807 59669
rect 458449 59668 458515 59669
rect 503253 59668 503319 59669
rect 413456 59666 413462 59668
rect 404169 59608 404174 59664
rect 403190 59604 403196 59606
rect 404169 59604 404214 59608
rect 404278 59606 404326 59666
rect 412541 59664 413462 59666
rect 412541 59608 412546 59664
rect 412602 59608 413462 59664
rect 412541 59606 413462 59608
rect 404278 59604 404284 59606
rect 57716 59470 84210 59530
rect 89989 59532 90055 59533
rect 95877 59532 95943 59533
rect 96981 59532 97047 59533
rect 98085 59532 98151 59533
rect 100753 59532 100819 59533
rect 89989 59528 90036 59532
rect 90100 59530 90106 59532
rect 89989 59472 89994 59528
rect 57716 59468 57722 59470
rect 89989 59468 90036 59472
rect 90100 59470 90146 59530
rect 95877 59528 95924 59532
rect 95988 59530 95994 59532
rect 95877 59472 95882 59528
rect 90100 59468 90106 59470
rect 95877 59468 95924 59472
rect 95988 59470 96034 59530
rect 96981 59528 97028 59532
rect 97092 59530 97098 59532
rect 96981 59472 96986 59528
rect 95988 59468 95994 59470
rect 96981 59468 97028 59472
rect 97092 59470 97138 59530
rect 98085 59528 98132 59532
rect 98196 59530 98202 59532
rect 100702 59530 100708 59532
rect 98085 59472 98090 59528
rect 97092 59468 97098 59470
rect 98085 59468 98132 59472
rect 98196 59470 98242 59530
rect 100662 59470 100708 59530
rect 100772 59528 100819 59532
rect 105976 59530 106036 59604
rect 107561 59603 107627 59604
rect 258073 59603 258139 59604
rect 260649 59603 260715 59604
rect 261753 59603 261819 59604
rect 308489 59603 308555 59604
rect 315849 59603 315915 59604
rect 403065 59603 403131 59604
rect 404169 59603 404235 59604
rect 412541 59603 412607 59606
rect 413456 59604 413462 59606
rect 413526 59604 413532 59668
rect 416037 59664 416046 59668
rect 416110 59666 416116 59668
rect 416037 59608 416042 59664
rect 416037 59604 416046 59608
rect 416110 59606 416194 59666
rect 416110 59604 416116 59606
rect 419440 59604 419446 59668
rect 419510 59666 419516 59668
rect 419510 59606 419598 59666
rect 421741 59664 421758 59668
rect 421822 59666 421828 59668
rect 421741 59608 421746 59664
rect 419510 59604 419516 59606
rect 421741 59604 421758 59608
rect 421822 59606 421898 59666
rect 458449 59664 458478 59668
rect 458542 59666 458548 59668
rect 503216 59666 503222 59668
rect 458449 59608 458454 59664
rect 421822 59604 421828 59606
rect 458449 59604 458478 59608
rect 458542 59606 458606 59666
rect 503162 59606 503222 59666
rect 503286 59664 503319 59668
rect 503314 59608 503319 59664
rect 458542 59604 458548 59606
rect 503216 59604 503222 59606
rect 503286 59604 503319 59608
rect 416037 59603 416103 59604
rect 419441 59603 419507 59604
rect 421741 59603 421807 59604
rect 458449 59603 458515 59604
rect 503253 59603 503319 59604
rect 100814 59472 100819 59528
rect 98196 59468 98202 59470
rect 100702 59468 100708 59470
rect 100772 59468 100819 59472
rect 89989 59467 90055 59468
rect 95877 59467 95943 59468
rect 96981 59467 97047 59468
rect 98085 59467 98151 59468
rect 100753 59467 100819 59468
rect 103470 59470 106036 59530
rect 410701 59532 410767 59533
rect 418153 59532 418219 59533
rect 410701 59528 410748 59532
rect 410812 59530 410818 59532
rect 418102 59530 418108 59532
rect 410701 59472 410706 59528
rect 46606 59332 46612 59396
rect 46676 59394 46682 59396
rect 103470 59394 103530 59470
rect 410701 59468 410748 59472
rect 410812 59470 410858 59530
rect 418062 59470 418108 59530
rect 418172 59528 418219 59532
rect 418214 59472 418219 59528
rect 410812 59468 410818 59470
rect 418102 59468 418108 59470
rect 418172 59468 418219 59472
rect 410701 59467 410767 59468
rect 418153 59467 418219 59468
rect 420637 59532 420703 59533
rect 420637 59528 420684 59532
rect 420748 59530 420754 59532
rect 420637 59472 420642 59528
rect 420637 59468 420684 59472
rect 420748 59470 420794 59530
rect 583520 59516 584960 59756
rect 420748 59468 420754 59470
rect 420637 59467 420703 59468
rect 46676 59334 103530 59394
rect 110965 59396 111031 59397
rect 279233 59396 279299 59397
rect 425973 59396 426039 59397
rect 428181 59396 428247 59397
rect 453389 59396 453455 59397
rect 110965 59392 111012 59396
rect 111076 59394 111082 59396
rect 110965 59336 110970 59392
rect 46676 59332 46682 59334
rect 110965 59332 111012 59336
rect 111076 59334 111122 59394
rect 111076 59332 111082 59334
rect 200798 59332 200804 59396
rect 200868 59394 200874 59396
rect 263542 59394 263548 59396
rect 200868 59334 263548 59394
rect 200868 59332 200874 59334
rect 263542 59332 263548 59334
rect 263612 59332 263618 59396
rect 279182 59394 279188 59396
rect 279142 59334 279188 59394
rect 279252 59392 279299 59396
rect 279294 59336 279299 59392
rect 279182 59332 279188 59334
rect 279252 59332 279299 59336
rect 377622 59332 377628 59396
rect 377692 59394 377698 59396
rect 422886 59394 422892 59396
rect 377692 59334 422892 59394
rect 377692 59332 377698 59334
rect 422886 59332 422892 59334
rect 422956 59332 422962 59396
rect 425973 59392 426020 59396
rect 426084 59394 426090 59396
rect 425973 59336 425978 59392
rect 425973 59332 426020 59336
rect 426084 59334 426130 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 426084 59332 426090 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 453389 59392 453436 59396
rect 453500 59394 453506 59396
rect 453389 59336 453394 59392
rect 428292 59332 428298 59334
rect 453389 59332 453436 59336
rect 453500 59334 453546 59394
rect 453500 59332 453506 59334
rect 110965 59331 111031 59332
rect 279233 59331 279299 59332
rect 425973 59331 426039 59332
rect 428181 59331 428247 59332
rect 453389 59331 453455 59332
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 290917 59260 290983 59261
rect 300853 59260 300919 59261
rect 320909 59260 320975 59261
rect 325877 59260 325943 59261
rect 54702 59196 54708 59260
rect 54772 59258 54778 59260
rect 143574 59258 143580 59260
rect 54772 59198 143580 59258
rect 54772 59196 54778 59198
rect 143574 59196 143580 59198
rect 143644 59196 143650 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 198406 59196 198412 59260
rect 198476 59258 198482 59260
rect 280838 59258 280844 59260
rect 198476 59198 280844 59258
rect 198476 59196 198482 59198
rect 280838 59196 280844 59198
rect 280908 59196 280914 59260
rect 290917 59256 290964 59260
rect 291028 59258 291034 59260
rect 290917 59200 290922 59256
rect 290917 59196 290964 59200
rect 291028 59198 291074 59258
rect 300853 59256 300900 59260
rect 300964 59258 300970 59260
rect 300853 59200 300858 59256
rect 291028 59196 291034 59198
rect 300853 59196 300900 59200
rect 300964 59198 301010 59258
rect 320909 59256 320956 59260
rect 321020 59258 321026 59260
rect 320909 59200 320914 59256
rect 300964 59196 300970 59198
rect 320909 59196 320956 59200
rect 321020 59198 321066 59258
rect 325877 59256 325924 59260
rect 325988 59258 325994 59260
rect 325877 59200 325882 59256
rect 321020 59196 321026 59198
rect 325877 59196 325924 59200
rect 325988 59198 326034 59258
rect 325988 59196 325994 59198
rect 357934 59196 357940 59260
rect 358004 59258 358010 59260
rect 480846 59258 480852 59260
rect 358004 59198 480852 59258
rect 358004 59196 358010 59198
rect 480846 59196 480852 59198
rect 480916 59196 480922 59260
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 290917 59195 290983 59196
rect 300853 59195 300919 59196
rect 320909 59195 320975 59196
rect 325877 59195 325943 59196
rect 55622 59060 55628 59124
rect 55692 59122 55698 59124
rect 140814 59122 140820 59124
rect 55692 59062 140820 59122
rect 55692 59060 55698 59062
rect 140814 59060 140820 59062
rect 140884 59060 140890 59124
rect 212390 59060 212396 59124
rect 212460 59122 212466 59124
rect 285990 59122 285996 59124
rect 212460 59062 285996 59122
rect 212460 59060 212466 59062
rect 285990 59060 285996 59062
rect 286060 59060 286066 59124
rect 371734 59060 371740 59124
rect 371804 59122 371810 59124
rect 483422 59122 483428 59124
rect 371804 59062 483428 59122
rect 371804 59060 371810 59062
rect 483422 59060 483428 59062
rect 483492 59060 483498 59124
rect 475837 58988 475903 58989
rect 53414 58924 53420 58988
rect 53484 58986 53490 58988
rect 138422 58986 138428 58988
rect 53484 58926 138428 58986
rect 53484 58924 53490 58926
rect 138422 58924 138428 58926
rect 138492 58924 138498 58988
rect 201350 58924 201356 58988
rect 201420 58986 201426 58988
rect 273478 58986 273484 58988
rect 201420 58926 273484 58986
rect 201420 58924 201426 58926
rect 273478 58924 273484 58926
rect 273548 58924 273554 58988
rect 367870 58924 367876 58988
rect 367940 58986 367946 58988
rect 468518 58986 468524 58988
rect 367940 58926 468524 58986
rect 367940 58924 367946 58926
rect 468518 58924 468524 58926
rect 468588 58924 468594 58988
rect 475837 58984 475884 58988
rect 475948 58986 475954 58988
rect 475837 58928 475842 58984
rect 475837 58924 475884 58928
rect 475948 58926 475994 58986
rect 475948 58924 475954 58926
rect 475837 58923 475903 58924
rect 52126 58788 52132 58852
rect 52196 58850 52202 58852
rect 135846 58850 135852 58852
rect 52196 58790 135852 58850
rect 52196 58788 52202 58790
rect 135846 58788 135852 58790
rect 135916 58788 135922 58852
rect 209630 58788 209636 58852
rect 209700 58850 209706 58852
rect 276054 58850 276060 58852
rect 209700 58790 276060 58850
rect 209700 58788 209706 58790
rect 276054 58788 276060 58790
rect 276124 58788 276130 58852
rect 375966 58788 375972 58852
rect 376036 58850 376042 58852
rect 473486 58850 473492 58852
rect 376036 58790 473492 58850
rect 376036 58788 376042 58790
rect 473486 58788 473492 58790
rect 473556 58788 473562 58852
rect -960 58578 480 58668
rect 59302 58652 59308 58716
rect 59372 58714 59378 58716
rect 120942 58714 120948 58716
rect 59372 58654 120948 58714
rect 59372 58652 59378 58654
rect 120942 58652 120948 58654
rect 121012 58652 121018 58716
rect 197854 58652 197860 58716
rect 197924 58714 197930 58716
rect 253606 58714 253612 58716
rect 197924 58654 253612 58714
rect 197924 58652 197930 58654
rect 253606 58652 253612 58654
rect 253676 58652 253682 58716
rect 374678 58652 374684 58716
rect 374748 58714 374754 58716
rect 463550 58714 463556 58716
rect 374748 58654 463556 58714
rect 374748 58652 374754 58654
rect 463550 58652 463556 58654
rect 463620 58652 463626 58716
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 48078 58516 48084 58580
rect 48148 58578 48154 58580
rect 108246 58578 108252 58580
rect 48148 58518 108252 58578
rect 48148 58516 48154 58518
rect 108246 58516 108252 58518
rect 108316 58516 108322 58580
rect 200614 58516 200620 58580
rect 200684 58578 200690 58580
rect 250662 58578 250668 58580
rect 200684 58518 250668 58578
rect 200684 58516 200690 58518
rect 250662 58516 250668 58518
rect 250732 58516 250738 58580
rect 59118 58380 59124 58444
rect 59188 58442 59194 58444
rect 101070 58442 101076 58444
rect 59188 58382 101076 58442
rect 59188 58380 59194 58382
rect 101070 58380 101076 58382
rect 101140 58380 101146 58444
rect 217358 58380 217364 58444
rect 217428 58442 217434 58444
rect 259494 58442 259500 58444
rect 217428 58382 259500 58442
rect 217428 58380 217434 58382
rect 259494 58380 259500 58382
rect 259564 58380 259570 58444
rect 85430 58108 85436 58172
rect 85500 58108 85506 58172
rect 92422 58108 92428 58172
rect 92492 58108 92498 58172
rect 99414 58108 99420 58172
rect 99484 58108 99490 58172
rect 113214 58108 113220 58172
rect 113284 58108 113290 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 235942 58108 235948 58172
rect 236012 58108 236018 58172
rect 265198 58108 265204 58172
rect 265268 58108 265274 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 398230 58108 398236 58172
rect 398300 58108 398306 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 405406 58108 405412 58172
rect 405476 58108 405482 58172
rect 455822 58108 455828 58172
rect 455892 58108 455898 58172
rect 83958 57972 83964 58036
rect 84028 58034 84034 58036
rect 84193 58034 84259 58037
rect 84028 58032 84259 58034
rect 84028 57976 84198 58032
rect 84254 57976 84259 58032
rect 84028 57974 84259 57976
rect 84028 57972 84034 57974
rect 84193 57971 84259 57974
rect 85438 57901 85498 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78673 57898 78739 57901
rect 80421 57900 80487 57901
rect 79542 57898 79548 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 78673 57896 79548 57898
rect 78673 57840 78678 57896
rect 78734 57840 79548 57896
rect 78673 57838 79548 57840
rect 78324 57836 78330 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 78673 57835 78739 57838
rect 79542 57836 79548 57838
rect 79612 57836 79618 57900
rect 80421 57896 80468 57900
rect 80532 57898 80538 57900
rect 81433 57898 81499 57901
rect 81934 57898 81940 57900
rect 80421 57840 80426 57896
rect 80421 57836 80468 57840
rect 80532 57838 80578 57898
rect 81433 57896 81940 57898
rect 81433 57840 81438 57896
rect 81494 57840 81940 57896
rect 81433 57838 81940 57840
rect 80532 57836 80538 57838
rect 80421 57835 80487 57836
rect 81433 57835 81499 57838
rect 81934 57836 81940 57838
rect 82004 57836 82010 57900
rect 85389 57896 85498 57901
rect 85389 57840 85394 57896
rect 85450 57840 85498 57896
rect 85389 57838 85498 57840
rect 86493 57900 86559 57901
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 88333 57900 88399 57901
rect 88701 57900 88767 57901
rect 90725 57900 90791 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 85389 57835 85455 57838
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88333 57896 88380 57900
rect 88444 57898 88450 57900
rect 88333 57840 88338 57896
rect 88333 57836 88380 57840
rect 88444 57838 88490 57898
rect 88701 57896 88748 57900
rect 88812 57898 88818 57900
rect 88701 57840 88706 57896
rect 88444 57836 88450 57838
rect 88701 57836 88748 57840
rect 88812 57838 88858 57898
rect 90725 57896 90772 57900
rect 90836 57898 90842 57900
rect 91093 57898 91159 57901
rect 91318 57898 91324 57900
rect 90725 57840 90730 57896
rect 88812 57836 88818 57838
rect 90725 57836 90772 57840
rect 90836 57838 90882 57898
rect 91093 57896 91324 57898
rect 91093 57840 91098 57896
rect 91154 57840 91324 57896
rect 91093 57838 91324 57840
rect 90836 57836 90842 57838
rect 88333 57835 88399 57836
rect 88701 57835 88767 57836
rect 90725 57835 90791 57836
rect 91093 57835 91159 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 91461 57898 91527 57901
rect 92430 57898 92490 58108
rect 99422 57901 99482 58108
rect 113222 57901 113282 58108
rect 153334 57901 153394 58108
rect 235950 57901 236010 58108
rect 93301 57900 93367 57901
rect 93669 57900 93735 57901
rect 93301 57898 93348 57900
rect 91461 57896 92490 57898
rect 91461 57840 91466 57896
rect 91522 57840 92490 57896
rect 91461 57838 92490 57840
rect 93256 57896 93348 57898
rect 93256 57840 93306 57896
rect 93256 57838 93348 57840
rect 91461 57835 91527 57838
rect 93301 57836 93348 57838
rect 93412 57836 93418 57900
rect 93669 57896 93716 57900
rect 93780 57898 93786 57900
rect 93669 57840 93674 57896
rect 93669 57836 93716 57840
rect 93780 57838 93826 57898
rect 99373 57896 99482 57901
rect 99373 57840 99378 57896
rect 99434 57840 99482 57896
rect 99373 57838 99482 57840
rect 103789 57900 103855 57901
rect 103789 57896 103836 57900
rect 103900 57898 103906 57900
rect 106273 57898 106339 57901
rect 106406 57898 106412 57900
rect 103789 57840 103794 57896
rect 93780 57836 93786 57838
rect 93301 57835 93367 57836
rect 93669 57835 93735 57836
rect 99373 57835 99439 57838
rect 103789 57836 103836 57840
rect 103900 57838 103946 57898
rect 106273 57896 106412 57898
rect 106273 57840 106278 57896
rect 106334 57840 106412 57896
rect 106273 57838 106412 57840
rect 103900 57836 103906 57838
rect 103789 57835 103855 57836
rect 106273 57835 106339 57838
rect 106406 57836 106412 57838
rect 106476 57836 106482 57900
rect 108205 57898 108271 57901
rect 108614 57898 108620 57900
rect 108205 57896 108620 57898
rect 108205 57840 108210 57896
rect 108266 57840 108620 57896
rect 108205 57838 108620 57840
rect 108205 57835 108271 57838
rect 108614 57836 108620 57838
rect 108684 57836 108690 57900
rect 109033 57898 109099 57901
rect 111149 57900 111215 57901
rect 112069 57900 112135 57901
rect 109534 57898 109540 57900
rect 109033 57896 109540 57898
rect 109033 57840 109038 57896
rect 109094 57840 109540 57896
rect 109033 57838 109540 57840
rect 109033 57835 109099 57838
rect 109534 57836 109540 57838
rect 109604 57836 109610 57900
rect 111149 57896 111196 57900
rect 111260 57898 111266 57900
rect 111149 57840 111154 57896
rect 111149 57836 111196 57840
rect 111260 57838 111306 57898
rect 112069 57896 112116 57900
rect 112180 57898 112186 57900
rect 112069 57840 112074 57896
rect 111260 57836 111266 57838
rect 112069 57836 112116 57840
rect 112180 57838 112226 57898
rect 113173 57896 113282 57901
rect 115749 57900 115815 57901
rect 115933 57900 115999 57901
rect 119061 57900 119127 57901
rect 130837 57900 130903 57901
rect 133413 57900 133479 57901
rect 145557 57900 145623 57901
rect 115749 57898 115796 57900
rect 113173 57840 113178 57896
rect 113234 57840 113282 57896
rect 113173 57838 113282 57840
rect 115704 57896 115796 57898
rect 115704 57840 115754 57896
rect 115704 57838 115796 57840
rect 112180 57836 112186 57838
rect 111149 57835 111215 57836
rect 112069 57835 112135 57836
rect 113173 57835 113239 57838
rect 115749 57836 115796 57838
rect 115860 57836 115866 57900
rect 115933 57896 115980 57900
rect 116044 57898 116050 57900
rect 115933 57840 115938 57896
rect 115933 57836 115980 57840
rect 116044 57838 116090 57898
rect 119061 57896 119108 57900
rect 119172 57898 119178 57900
rect 119061 57840 119066 57896
rect 116044 57836 116050 57838
rect 119061 57836 119108 57840
rect 119172 57838 119218 57898
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 130837 57840 130842 57896
rect 119172 57836 119178 57838
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 133413 57896 133460 57900
rect 133524 57898 133530 57900
rect 133413 57840 133418 57896
rect 130948 57836 130954 57838
rect 133413 57836 133460 57840
rect 133524 57838 133570 57898
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 133524 57836 133530 57838
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 183461 57900 183527 57901
rect 183461 57896 183508 57900
rect 183572 57898 183578 57900
rect 183461 57840 183466 57896
rect 145668 57836 145674 57838
rect 115749 57835 115815 57836
rect 115933 57835 115999 57836
rect 119061 57835 119127 57836
rect 130837 57835 130903 57836
rect 133413 57835 133479 57836
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 183461 57836 183508 57840
rect 183572 57838 183618 57898
rect 235950 57896 236059 57901
rect 235950 57840 235998 57896
rect 236054 57840 236059 57896
rect 235950 57838 236059 57840
rect 183572 57836 183578 57838
rect 183461 57835 183527 57836
rect 235993 57835 236059 57838
rect 237373 57898 237439 57901
rect 239213 57900 239279 57901
rect 238150 57898 238156 57900
rect 237373 57896 238156 57898
rect 237373 57840 237378 57896
rect 237434 57840 238156 57896
rect 237373 57838 238156 57840
rect 237373 57835 237439 57838
rect 238150 57836 238156 57838
rect 238220 57836 238226 57900
rect 239213 57896 239260 57900
rect 239324 57898 239330 57900
rect 240133 57898 240199 57901
rect 241605 57900 241671 57901
rect 242893 57900 242959 57901
rect 240542 57898 240548 57900
rect 239213 57840 239218 57896
rect 239213 57836 239260 57840
rect 239324 57838 239370 57898
rect 240133 57896 240548 57898
rect 240133 57840 240138 57896
rect 240194 57840 240548 57896
rect 240133 57838 240548 57840
rect 239324 57836 239330 57838
rect 239213 57835 239279 57836
rect 240133 57835 240199 57838
rect 240542 57836 240548 57838
rect 240612 57836 240618 57900
rect 241605 57896 241652 57900
rect 241716 57898 241722 57900
rect 241605 57840 241610 57896
rect 241605 57836 241652 57840
rect 241716 57838 241762 57898
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 242893 57840 242898 57896
rect 241716 57836 241722 57838
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 243004 57836 243010 57838
rect 244222 57836 244228 57900
rect 244292 57898 244298 57900
rect 244365 57898 244431 57901
rect 244292 57896 244431 57898
rect 244292 57840 244370 57896
rect 244426 57840 244431 57896
rect 244292 57838 244431 57840
rect 244292 57836 244298 57838
rect 241605 57835 241671 57836
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245285 57900 245351 57901
rect 245285 57896 245332 57900
rect 245396 57898 245402 57900
rect 245653 57898 245719 57901
rect 246430 57898 246436 57900
rect 245285 57840 245290 57896
rect 245285 57836 245332 57840
rect 245396 57838 245442 57898
rect 245653 57896 246436 57898
rect 245653 57840 245658 57896
rect 245714 57840 246436 57896
rect 245653 57838 246436 57840
rect 245396 57836 245402 57838
rect 245285 57835 245351 57836
rect 245653 57835 245719 57838
rect 246430 57836 246436 57838
rect 246500 57836 246506 57900
rect 247033 57898 247099 57901
rect 248229 57900 248295 57901
rect 248597 57900 248663 57901
rect 247718 57898 247724 57900
rect 247033 57896 247724 57898
rect 247033 57840 247038 57896
rect 247094 57840 247724 57896
rect 247033 57838 247724 57840
rect 247033 57835 247099 57838
rect 247718 57836 247724 57838
rect 247788 57836 247794 57900
rect 248229 57896 248276 57900
rect 248340 57898 248346 57900
rect 248229 57840 248234 57896
rect 248229 57836 248276 57840
rect 248340 57838 248386 57898
rect 248597 57896 248644 57900
rect 248708 57898 248714 57900
rect 249793 57898 249859 57901
rect 251173 57900 251239 57901
rect 250110 57898 250116 57900
rect 248597 57840 248602 57896
rect 248340 57836 248346 57838
rect 248597 57836 248644 57840
rect 248708 57838 248754 57898
rect 249793 57896 250116 57898
rect 249793 57840 249798 57896
rect 249854 57840 250116 57896
rect 249793 57838 250116 57840
rect 248708 57836 248714 57838
rect 248229 57835 248295 57836
rect 248597 57835 248663 57836
rect 249793 57835 249859 57838
rect 250110 57836 250116 57838
rect 250180 57836 250186 57900
rect 251173 57898 251220 57900
rect 251128 57896 251220 57898
rect 251128 57840 251178 57896
rect 251128 57838 251220 57840
rect 251173 57836 251220 57838
rect 251284 57836 251290 57900
rect 251357 57898 251423 57901
rect 253381 57900 253447 57901
rect 252318 57898 252324 57900
rect 251357 57896 252324 57898
rect 251357 57840 251362 57896
rect 251418 57840 252324 57896
rect 251357 57838 252324 57840
rect 251173 57835 251239 57836
rect 251357 57835 251423 57838
rect 252318 57836 252324 57838
rect 252388 57836 252394 57900
rect 253381 57896 253428 57900
rect 253492 57898 253498 57900
rect 253933 57898 253999 57901
rect 258349 57900 258415 57901
rect 254526 57898 254532 57900
rect 253381 57840 253386 57896
rect 253381 57836 253428 57840
rect 253492 57838 253538 57898
rect 253933 57896 254532 57898
rect 253933 57840 253938 57896
rect 253994 57840 254532 57896
rect 253933 57838 254532 57840
rect 253492 57836 253498 57838
rect 253381 57835 253447 57836
rect 253933 57835 253999 57838
rect 254526 57836 254532 57838
rect 254596 57836 254602 57900
rect 258349 57896 258396 57900
rect 258460 57898 258466 57900
rect 264973 57898 265039 57901
rect 265206 57898 265266 58108
rect 258349 57840 258354 57896
rect 258349 57836 258396 57840
rect 258460 57838 258506 57898
rect 264973 57896 265266 57898
rect 264973 57840 264978 57896
rect 265034 57840 265266 57896
rect 264973 57838 265266 57840
rect 266445 57898 266511 57901
rect 267590 57898 267596 57900
rect 266445 57896 267596 57898
rect 266445 57840 266450 57896
rect 266506 57840 267596 57896
rect 266445 57838 267596 57840
rect 258460 57836 258466 57838
rect 258349 57835 258415 57836
rect 264973 57835 265039 57838
rect 266445 57835 266511 57838
rect 267590 57836 267596 57838
rect 267660 57836 267666 57900
rect 268101 57898 268167 57901
rect 268694 57898 268700 57900
rect 268101 57896 268700 57898
rect 268101 57840 268106 57896
rect 268162 57840 268700 57896
rect 268101 57838 268700 57840
rect 268101 57835 268167 57838
rect 268694 57836 268700 57838
rect 268764 57836 268770 57900
rect 268929 57898 268995 57901
rect 271045 57900 271111 57901
rect 270902 57898 270908 57900
rect 268929 57896 270908 57898
rect 268929 57840 268934 57896
rect 268990 57840 270908 57896
rect 268929 57838 270908 57840
rect 268929 57835 268995 57838
rect 270902 57836 270908 57838
rect 270972 57836 270978 57900
rect 271045 57896 271092 57900
rect 271156 57898 271162 57900
rect 271873 57898 271939 57901
rect 272198 57898 272258 58108
rect 271045 57840 271050 57896
rect 271045 57836 271092 57840
rect 271156 57838 271202 57898
rect 271873 57896 272258 57898
rect 271873 57840 271878 57896
rect 271934 57840 272258 57896
rect 271873 57838 272258 57840
rect 273253 57900 273319 57901
rect 273253 57896 273300 57900
rect 273364 57898 273370 57900
rect 275093 57898 275159 57901
rect 275694 57898 275754 58108
rect 273253 57840 273258 57896
rect 271156 57836 271162 57838
rect 271045 57835 271111 57836
rect 271873 57835 271939 57838
rect 273253 57836 273300 57840
rect 273364 57838 273410 57898
rect 275093 57896 275754 57898
rect 275093 57840 275098 57896
rect 275154 57840 275754 57896
rect 275093 57838 275754 57840
rect 276933 57900 276999 57901
rect 276933 57896 276980 57900
rect 277044 57898 277050 57900
rect 278313 57898 278379 57901
rect 295885 57900 295951 57901
rect 278446 57898 278452 57900
rect 276933 57840 276938 57896
rect 273364 57836 273370 57838
rect 273253 57835 273319 57836
rect 275093 57835 275159 57838
rect 276933 57836 276980 57840
rect 277044 57838 277090 57898
rect 278313 57896 278452 57898
rect 278313 57840 278318 57896
rect 278374 57840 278452 57896
rect 278313 57838 278452 57840
rect 277044 57836 277050 57838
rect 276933 57835 276999 57836
rect 278313 57835 278379 57838
rect 278446 57836 278452 57838
rect 278516 57836 278522 57900
rect 295885 57896 295932 57900
rect 295996 57898 296002 57900
rect 298093 57898 298159 57901
rect 303429 57900 303495 57901
rect 305821 57900 305887 57901
rect 310973 57900 311039 57901
rect 313365 57900 313431 57901
rect 298502 57898 298508 57900
rect 295885 57840 295890 57896
rect 295885 57836 295932 57840
rect 295996 57838 296042 57898
rect 298093 57896 298508 57898
rect 298093 57840 298098 57896
rect 298154 57840 298508 57896
rect 298093 57838 298508 57840
rect 295996 57836 296002 57838
rect 295885 57835 295951 57836
rect 298093 57835 298159 57838
rect 298502 57836 298508 57838
rect 298572 57836 298578 57900
rect 303429 57896 303476 57900
rect 303540 57898 303546 57900
rect 303429 57840 303434 57896
rect 303429 57836 303476 57840
rect 303540 57838 303586 57898
rect 305821 57896 305868 57900
rect 305932 57898 305938 57900
rect 305821 57840 305826 57896
rect 303540 57836 303546 57838
rect 305821 57836 305868 57840
rect 305932 57838 305978 57898
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 305932 57836 305938 57838
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 313365 57896 313412 57900
rect 313476 57898 313482 57900
rect 318241 57898 318307 57901
rect 323301 57900 323367 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 318374 57898 318380 57900
rect 313365 57840 313370 57896
rect 311084 57836 311090 57838
rect 313365 57836 313412 57840
rect 313476 57838 313522 57898
rect 318241 57896 318380 57898
rect 318241 57840 318246 57896
rect 318302 57840 318380 57896
rect 318241 57838 318380 57840
rect 313476 57836 313482 57838
rect 303429 57835 303495 57836
rect 305821 57835 305887 57836
rect 310973 57835 311039 57836
rect 313365 57835 313431 57836
rect 318241 57835 318307 57838
rect 318374 57836 318380 57838
rect 318444 57836 318450 57900
rect 323301 57896 323348 57900
rect 323412 57898 323418 57900
rect 343173 57898 343220 57900
rect 323301 57840 323306 57896
rect 323301 57836 323348 57840
rect 323412 57838 323458 57898
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 323412 57836 323418 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 323301 57835 323367 57836
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 397453 57898 397519 57901
rect 398238 57898 398298 58108
rect 401734 57901 401794 58108
rect 397453 57896 398298 57898
rect 397453 57840 397458 57896
rect 397514 57840 398298 57896
rect 397453 57838 398298 57840
rect 399477 57900 399543 57901
rect 399477 57896 399524 57900
rect 399588 57898 399594 57900
rect 400213 57898 400279 57901
rect 400438 57898 400444 57900
rect 399477 57840 399482 57896
rect 397453 57835 397519 57838
rect 399477 57836 399524 57840
rect 399588 57838 399634 57898
rect 400213 57896 400444 57898
rect 400213 57840 400218 57896
rect 400274 57840 400444 57896
rect 400213 57838 400444 57840
rect 399588 57836 399594 57838
rect 399477 57835 399543 57836
rect 400213 57835 400279 57838
rect 400438 57836 400444 57838
rect 400508 57836 400514 57900
rect 401685 57896 401794 57901
rect 401685 57840 401690 57896
rect 401746 57840 401794 57896
rect 401685 57838 401794 57840
rect 404353 57898 404419 57901
rect 405414 57898 405474 58108
rect 404353 57896 405474 57898
rect 404353 57840 404358 57896
rect 404414 57840 405474 57896
rect 404353 57838 405474 57840
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 401685 57835 401751 57838
rect 404353 57835 404419 57838
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407205 57898 407271 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407205 57896 407620 57898
rect 407205 57840 407210 57896
rect 407266 57840 407620 57896
rect 407205 57838 407620 57840
rect 407205 57835 407271 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 414565 57900 414631 57901
rect 415485 57900 415551 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 414565 57896 414612 57900
rect 414676 57898 414682 57900
rect 414565 57840 414570 57896
rect 414565 57836 414612 57840
rect 414676 57838 414722 57898
rect 415485 57896 415532 57900
rect 415596 57898 415602 57900
rect 415485 57840 415490 57896
rect 414676 57836 414682 57838
rect 415485 57836 415532 57840
rect 415596 57838 415642 57898
rect 415596 57836 415602 57838
rect 426382 57836 426388 57900
rect 426452 57898 426458 57900
rect 426525 57898 426591 57901
rect 427629 57900 427695 57901
rect 427629 57898 427676 57900
rect 426452 57896 426591 57898
rect 426452 57840 426530 57896
rect 426586 57840 426591 57896
rect 426452 57838 426591 57840
rect 427584 57896 427676 57898
rect 427584 57840 427634 57896
rect 427584 57838 427676 57840
rect 426452 57836 426458 57838
rect 414565 57835 414631 57836
rect 415485 57835 415551 57836
rect 426525 57835 426591 57838
rect 427629 57836 427676 57838
rect 427740 57836 427746 57900
rect 427813 57898 427879 57901
rect 428590 57898 428596 57900
rect 427813 57896 428596 57898
rect 427813 57840 427818 57896
rect 427874 57840 428596 57896
rect 427813 57838 428596 57840
rect 427629 57835 427695 57836
rect 427813 57835 427879 57838
rect 428590 57836 428596 57838
rect 428660 57836 428666 57900
rect 429193 57898 429259 57901
rect 429694 57898 429700 57900
rect 429193 57896 429700 57898
rect 429193 57840 429198 57896
rect 429254 57840 429700 57896
rect 429193 57838 429700 57840
rect 429193 57835 429259 57838
rect 429694 57836 429700 57838
rect 429764 57836 429770 57900
rect 430573 57898 430639 57901
rect 432229 57900 432295 57901
rect 431166 57898 431172 57900
rect 430573 57896 431172 57898
rect 430573 57840 430578 57896
rect 430634 57840 431172 57896
rect 430573 57838 431172 57840
rect 430573 57835 430639 57838
rect 431166 57836 431172 57838
rect 431236 57836 431242 57900
rect 432229 57896 432276 57900
rect 432340 57898 432346 57900
rect 434437 57898 434503 57901
rect 435909 57900 435975 57901
rect 434662 57898 434668 57900
rect 432229 57840 432234 57896
rect 432229 57836 432276 57840
rect 432340 57838 432386 57898
rect 434437 57896 434668 57898
rect 434437 57840 434442 57896
rect 434498 57840 434668 57896
rect 434437 57838 434668 57840
rect 432340 57836 432346 57838
rect 432229 57835 432295 57836
rect 434437 57835 434503 57838
rect 434662 57836 434668 57838
rect 434732 57836 434738 57900
rect 435909 57896 435956 57900
rect 436020 57898 436026 57900
rect 436277 57898 436343 57901
rect 438485 57900 438551 57901
rect 445845 57900 445911 57901
rect 450997 57900 451063 57901
rect 436870 57898 436876 57900
rect 435909 57840 435914 57896
rect 435909 57836 435956 57840
rect 436020 57838 436066 57898
rect 436277 57896 436876 57898
rect 436277 57840 436282 57896
rect 436338 57840 436876 57896
rect 436277 57838 436876 57840
rect 436020 57836 436026 57838
rect 435909 57835 435975 57836
rect 436277 57835 436343 57838
rect 436870 57836 436876 57838
rect 436940 57836 436946 57900
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 438485 57840 438490 57896
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 445845 57896 445892 57900
rect 445956 57898 445962 57900
rect 445845 57840 445850 57896
rect 438596 57836 438602 57838
rect 445845 57836 445892 57840
rect 445956 57838 446002 57898
rect 450997 57896 451044 57900
rect 451108 57898 451114 57900
rect 455830 57898 455890 58108
rect 450997 57840 451002 57896
rect 445956 57836 445962 57838
rect 450997 57836 451044 57840
rect 451108 57838 451154 57898
rect 451230 57838 455890 57898
rect 460933 57900 460999 57901
rect 465901 57900 465967 57901
rect 470869 57900 470935 57901
rect 478413 57900 478479 57901
rect 485957 57900 486023 57901
rect 503345 57900 503411 57901
rect 460933 57896 460980 57900
rect 461044 57898 461050 57900
rect 460933 57840 460938 57896
rect 451108 57836 451114 57838
rect 438485 57835 438551 57836
rect 445845 57835 445911 57836
rect 450997 57835 451063 57836
rect 183185 57764 183251 57765
rect 60222 57700 60228 57764
rect 60292 57762 60298 57764
rect 125910 57762 125916 57764
rect 60292 57702 125916 57762
rect 60292 57700 60298 57702
rect 125910 57700 125916 57702
rect 125980 57700 125986 57764
rect 183134 57762 183140 57764
rect 183094 57702 183140 57762
rect 183204 57760 183251 57764
rect 183246 57704 183251 57760
rect 183134 57700 183140 57702
rect 183204 57700 183251 57704
rect 214414 57700 214420 57764
rect 214484 57762 214490 57764
rect 288198 57762 288204 57764
rect 214484 57702 288204 57762
rect 214484 57700 214490 57702
rect 288198 57700 288204 57702
rect 288268 57700 288274 57764
rect 374494 57700 374500 57764
rect 374564 57762 374570 57764
rect 451230 57762 451290 57838
rect 460933 57836 460980 57840
rect 461044 57838 461090 57898
rect 465901 57896 465948 57900
rect 466012 57898 466018 57900
rect 465901 57840 465906 57896
rect 461044 57836 461050 57838
rect 465901 57836 465948 57840
rect 466012 57838 466058 57898
rect 470869 57896 470916 57900
rect 470980 57898 470986 57900
rect 470869 57840 470874 57896
rect 466012 57836 466018 57838
rect 470869 57836 470916 57840
rect 470980 57838 471026 57898
rect 478413 57896 478460 57900
rect 478524 57898 478530 57900
rect 478413 57840 478418 57896
rect 470980 57836 470986 57838
rect 478413 57836 478460 57840
rect 478524 57838 478570 57898
rect 485957 57896 486004 57900
rect 486068 57898 486074 57900
rect 503294 57898 503300 57900
rect 485957 57840 485962 57896
rect 478524 57836 478530 57838
rect 485957 57836 486004 57840
rect 486068 57838 486114 57898
rect 503254 57838 503300 57898
rect 503364 57896 503411 57900
rect 503406 57840 503411 57896
rect 486068 57836 486074 57838
rect 503294 57836 503300 57838
rect 503364 57836 503411 57840
rect 460933 57835 460999 57836
rect 465901 57835 465967 57836
rect 470869 57835 470935 57836
rect 478413 57835 478479 57836
rect 485957 57835 486023 57836
rect 503345 57835 503411 57836
rect 374564 57702 451290 57762
rect 374564 57700 374570 57702
rect 183185 57699 183251 57700
rect 54886 57564 54892 57628
rect 54956 57626 54962 57628
rect 115841 57626 115907 57629
rect 54956 57624 115907 57626
rect 54956 57568 115846 57624
rect 115902 57568 115907 57624
rect 54956 57566 115907 57568
rect 54956 57564 54962 57566
rect 115841 57563 115907 57566
rect 116117 57626 116183 57629
rect 116894 57626 116900 57628
rect 116117 57624 116900 57626
rect 116117 57568 116122 57624
rect 116178 57568 116900 57624
rect 116117 57566 116900 57568
rect 116117 57563 116183 57566
rect 116894 57564 116900 57566
rect 116964 57564 116970 57628
rect 122833 57626 122899 57629
rect 123518 57626 123524 57628
rect 122833 57624 123524 57626
rect 122833 57568 122838 57624
rect 122894 57568 123524 57624
rect 122833 57566 123524 57568
rect 122833 57563 122899 57566
rect 123518 57564 123524 57566
rect 123588 57564 123594 57628
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 162853 57626 162919 57629
rect 163262 57626 163268 57628
rect 162853 57624 163268 57626
rect 162853 57568 162858 57624
rect 162914 57568 163268 57624
rect 162853 57566 163268 57568
rect 162853 57563 162919 57566
rect 163262 57564 163268 57566
rect 163332 57564 163338 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 202270 57564 202276 57628
rect 202340 57626 202346 57628
rect 268929 57626 268995 57629
rect 202340 57624 268995 57626
rect 202340 57568 268934 57624
rect 268990 57568 268995 57624
rect 202340 57566 268995 57568
rect 202340 57564 202346 57566
rect 268929 57563 268995 57566
rect 269113 57626 269179 57629
rect 269798 57626 269804 57628
rect 269113 57624 269804 57626
rect 269113 57568 269118 57624
rect 269174 57568 269804 57624
rect 269113 57566 269804 57568
rect 269113 57563 269179 57566
rect 269798 57564 269804 57566
rect 269868 57564 269874 57628
rect 273345 57626 273411 57629
rect 274398 57626 274404 57628
rect 273345 57624 274404 57626
rect 273345 57568 273350 57624
rect 273406 57568 274404 57624
rect 273345 57566 274404 57568
rect 273345 57563 273411 57566
rect 274398 57564 274404 57566
rect 274468 57564 274474 57628
rect 277393 57626 277459 57629
rect 278078 57626 278084 57628
rect 277393 57624 278084 57626
rect 277393 57568 277398 57624
rect 277454 57568 278084 57624
rect 277393 57566 278084 57568
rect 277393 57563 277459 57566
rect 278078 57564 278084 57566
rect 278148 57564 278154 57628
rect 370446 57564 370452 57628
rect 370516 57626 370522 57628
rect 433149 57626 433215 57629
rect 433425 57628 433491 57629
rect 433374 57626 433380 57628
rect 370516 57624 433215 57626
rect 370516 57568 433154 57624
rect 433210 57568 433215 57624
rect 370516 57566 433215 57568
rect 433334 57566 433380 57626
rect 433444 57624 433491 57628
rect 433486 57568 433491 57624
rect 370516 57564 370522 57566
rect 433149 57563 433215 57566
rect 433374 57564 433380 57566
rect 433444 57564 433491 57568
rect 433425 57563 433491 57564
rect 434713 57626 434779 57629
rect 435766 57626 435772 57628
rect 434713 57624 435772 57626
rect 434713 57568 434718 57624
rect 434774 57568 435772 57624
rect 434713 57566 435772 57568
rect 434713 57563 434779 57566
rect 435766 57564 435772 57566
rect 435836 57564 435842 57628
rect 437473 57626 437539 57629
rect 438342 57626 438348 57628
rect 437473 57624 438348 57626
rect 437473 57568 437478 57624
rect 437534 57568 438348 57624
rect 437473 57566 438348 57568
rect 437473 57563 437539 57566
rect 438342 57564 438348 57566
rect 438412 57564 438418 57628
rect 57830 57428 57836 57492
rect 57900 57490 57906 57492
rect 117998 57490 118004 57492
rect 57900 57430 118004 57490
rect 57900 57428 57906 57430
rect 117998 57428 118004 57430
rect 118068 57428 118074 57492
rect 216070 57428 216076 57492
rect 216140 57490 216146 57492
rect 283782 57490 283788 57492
rect 216140 57430 283788 57490
rect 216140 57428 216146 57430
rect 283782 57428 283788 57430
rect 283852 57428 283858 57492
rect 379094 57428 379100 57492
rect 379164 57490 379170 57492
rect 448278 57490 448284 57492
rect 379164 57430 448284 57490
rect 379164 57428 379170 57430
rect 448278 57428 448284 57430
rect 448348 57428 448354 57492
rect 58566 57292 58572 57356
rect 58636 57354 58642 57356
rect 58636 57294 98746 57354
rect 58636 57292 58642 57294
rect 58934 57156 58940 57220
rect 59004 57218 59010 57220
rect 98494 57218 98500 57220
rect 59004 57158 98500 57218
rect 59004 57156 59010 57158
rect 98494 57156 98500 57158
rect 98564 57156 98570 57220
rect 98686 57218 98746 57294
rect 113030 57292 113036 57356
rect 113100 57354 113106 57356
rect 113265 57354 113331 57357
rect 113100 57352 113331 57354
rect 113100 57296 113270 57352
rect 113326 57296 113331 57352
rect 113100 57294 113331 57296
rect 113100 57292 113106 57294
rect 113265 57291 113331 57294
rect 115841 57354 115907 57357
rect 266353 57356 266419 57357
rect 118366 57354 118372 57356
rect 115841 57352 118372 57354
rect 115841 57296 115846 57352
rect 115902 57296 118372 57352
rect 115841 57294 118372 57296
rect 115841 57291 115907 57294
rect 118366 57292 118372 57294
rect 118436 57292 118442 57356
rect 203190 57292 203196 57356
rect 203260 57354 203266 57356
rect 255998 57354 256004 57356
rect 203260 57294 256004 57354
rect 203260 57292 203266 57294
rect 255998 57292 256004 57294
rect 256068 57292 256074 57356
rect 266302 57354 266308 57356
rect 266262 57294 266308 57354
rect 266372 57352 266419 57356
rect 266414 57296 266419 57352
rect 266302 57292 266308 57294
rect 266372 57292 266419 57296
rect 371918 57292 371924 57356
rect 371988 57354 371994 57356
rect 433558 57354 433564 57356
rect 371988 57294 433564 57354
rect 371988 57292 371994 57294
rect 433558 57292 433564 57294
rect 433628 57292 433634 57356
rect 266353 57291 266419 57292
rect 430941 57220 431007 57221
rect 103830 57218 103836 57220
rect 98686 57158 103836 57218
rect 103830 57156 103836 57158
rect 103900 57156 103906 57220
rect 113214 57156 113220 57220
rect 113284 57218 113290 57220
rect 114318 57218 114324 57220
rect 113284 57158 114324 57218
rect 113284 57156 113290 57158
rect 114318 57156 114324 57158
rect 114388 57156 114394 57220
rect 213126 57156 213132 57220
rect 213196 57218 213202 57220
rect 265934 57218 265940 57220
rect 213196 57158 265940 57218
rect 213196 57156 213202 57158
rect 265934 57156 265940 57158
rect 266004 57156 266010 57220
rect 378910 57156 378916 57220
rect 378980 57218 378986 57220
rect 418470 57218 418476 57220
rect 378980 57158 418476 57218
rect 378980 57156 378986 57158
rect 418470 57156 418476 57158
rect 418540 57156 418546 57220
rect 430941 57216 430988 57220
rect 431052 57218 431058 57220
rect 433149 57218 433215 57221
rect 440918 57218 440924 57220
rect 430941 57160 430946 57216
rect 430941 57156 430988 57160
rect 431052 57158 431098 57218
rect 433149 57216 440924 57218
rect 433149 57160 433154 57216
rect 433210 57160 440924 57216
rect 433149 57158 440924 57160
rect 431052 57156 431058 57158
rect 430941 57155 431007 57156
rect 433149 57155 433215 57158
rect 440918 57156 440924 57158
rect 440988 57156 440994 57220
rect 58750 57020 58756 57084
rect 58820 57082 58826 57084
rect 96286 57082 96292 57084
rect 58820 57022 96292 57082
rect 58820 57020 58826 57022
rect 96286 57020 96292 57022
rect 96356 57020 96362 57084
rect 215886 57020 215892 57084
rect 215956 57082 215962 57084
rect 260966 57082 260972 57084
rect 215956 57022 260972 57082
rect 215956 57020 215962 57022
rect 260966 57020 260972 57022
rect 261036 57020 261042 57084
rect 378726 57020 378732 57084
rect 378796 57082 378802 57084
rect 413502 57082 413508 57084
rect 378796 57022 413508 57082
rect 378796 57020 378802 57022
rect 413502 57020 413508 57022
rect 413572 57020 413578 57084
rect 411253 56948 411319 56949
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 412541 56946 412607 56949
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 412541 56944 412650 56946
rect 412541 56888 412546 56944
rect 412602 56888 412650 56944
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 412541 56883 412650 56888
rect 412590 56813 412650 56883
rect 412590 56808 412699 56813
rect 443494 56810 443500 56812
rect 412590 56752 412638 56808
rect 412694 56752 412699 56808
rect 412590 56750 412699 56752
rect 412633 56747 412699 56750
rect 431910 56750 443500 56810
rect 55070 56612 55076 56676
rect 55140 56674 55146 56676
rect 128670 56674 128676 56676
rect 55140 56614 128676 56674
rect 55140 56612 55146 56614
rect 128670 56612 128676 56614
rect 128740 56612 128746 56676
rect 155902 56612 155908 56676
rect 155972 56612 155978 56676
rect 158478 56612 158484 56676
rect 158548 56612 158554 56676
rect 210550 56612 210556 56676
rect 210620 56674 210626 56676
rect 293350 56674 293356 56676
rect 210620 56614 293356 56674
rect 210620 56612 210626 56614
rect 293350 56612 293356 56614
rect 293420 56612 293426 56676
rect 358118 56612 358124 56676
rect 358188 56674 358194 56676
rect 431910 56674 431970 56750
rect 443494 56748 443500 56750
rect 443564 56748 443570 56812
rect 358188 56614 431970 56674
rect 358188 56612 358194 56614
rect 439078 56612 439084 56676
rect 439148 56612 439154 56676
rect 50838 56476 50844 56540
rect 50908 56538 50914 56540
rect 155910 56538 155970 56612
rect 50908 56478 155970 56538
rect 50908 56476 50914 56478
rect 53598 56340 53604 56404
rect 53668 56402 53674 56404
rect 158486 56402 158546 56612
rect 219934 56476 219940 56540
rect 220004 56538 220010 56540
rect 421046 56538 421052 56540
rect 220004 56478 421052 56538
rect 220004 56476 220010 56478
rect 421046 56476 421052 56478
rect 421116 56476 421122 56540
rect 439086 56538 439146 56612
rect 431910 56478 439146 56538
rect 53668 56342 158546 56402
rect 53668 56340 53674 56342
rect 198590 56340 198596 56404
rect 198660 56402 198666 56404
rect 268326 56402 268332 56404
rect 198660 56342 268332 56402
rect 198660 56340 198666 56342
rect 268326 56340 268332 56342
rect 268396 56340 268402 56404
rect 377438 56340 377444 56404
rect 377508 56402 377514 56404
rect 431910 56402 431970 56478
rect 377508 56342 431970 56402
rect 377508 56340 377514 56342
rect 51758 56204 51764 56268
rect 51828 56266 51834 56268
rect 153285 56266 153351 56269
rect 51828 56264 153351 56266
rect 51828 56208 153290 56264
rect 153346 56208 153351 56264
rect 51828 56206 153351 56208
rect 51828 56204 51834 56206
rect 153285 56203 153351 56206
rect 377806 56204 377812 56268
rect 377876 56266 377882 56268
rect 425278 56266 425284 56268
rect 377876 56206 425284 56266
rect 377876 56204 377882 56206
rect 425278 56204 425284 56206
rect 425348 56204 425354 56268
rect 57462 56068 57468 56132
rect 57532 56130 57538 56132
rect 119061 56130 119127 56133
rect 57532 56128 119127 56130
rect 57532 56072 119066 56128
rect 119122 56072 119127 56128
rect 57532 56070 119127 56072
rect 57532 56068 57538 56070
rect 119061 56067 119127 56070
rect 48630 55116 48636 55180
rect 48700 55178 48706 55180
rect 165613 55178 165679 55181
rect 48700 55176 165679 55178
rect 48700 55120 165618 55176
rect 165674 55120 165679 55176
rect 48700 55118 165679 55120
rect 48700 55116 48706 55118
rect 165613 55115 165679 55118
rect 214465 55178 214531 55181
rect 269113 55178 269179 55181
rect 214465 55176 269179 55178
rect 214465 55120 214470 55176
rect 214526 55120 269118 55176
rect 269174 55120 269179 55176
rect 214465 55118 269179 55120
rect 214465 55115 214531 55118
rect 269113 55115 269179 55118
rect 50654 54980 50660 55044
rect 50724 55042 50730 55044
rect 162853 55042 162919 55045
rect 50724 55040 162919 55042
rect 50724 54984 162858 55040
rect 162914 54984 162919 55040
rect 50724 54982 162919 54984
rect 50724 54980 50730 54982
rect 162853 54979 162919 54982
rect 55438 54844 55444 54908
rect 55508 54906 55514 54908
rect 160093 54906 160159 54909
rect 55508 54904 160159 54906
rect 55508 54848 160098 54904
rect 160154 54848 160159 54904
rect 55508 54846 160159 54848
rect 55508 54844 55514 54846
rect 160093 54843 160159 54846
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 140037 4042 140103 4045
rect 210366 4042 210372 4044
rect 140037 4040 210372 4042
rect 140037 3984 140042 4040
rect 140098 3984 210372 4040
rect 140037 3982 210372 3984
rect 140037 3979 140103 3982
rect 210366 3980 210372 3982
rect 210436 3980 210442 4044
rect 129365 3906 129431 3909
rect 202086 3906 202092 3908
rect 129365 3904 202092 3906
rect 129365 3848 129370 3904
rect 129426 3848 202092 3904
rect 129365 3846 202092 3848
rect 129365 3843 129431 3846
rect 202086 3844 202092 3846
rect 202156 3844 202162 3908
rect 147121 3770 147187 3773
rect 360694 3770 360700 3772
rect 147121 3768 360700 3770
rect 147121 3712 147126 3768
rect 147182 3712 360700 3768
rect 147121 3710 360700 3712
rect 147121 3707 147187 3710
rect 360694 3708 360700 3710
rect 360764 3708 360770 3772
rect 150617 3634 150683 3637
rect 364926 3634 364932 3636
rect 150617 3632 364932 3634
rect 150617 3576 150622 3632
rect 150678 3576 364932 3632
rect 150617 3574 364932 3576
rect 150617 3571 150683 3574
rect 364926 3572 364932 3574
rect 364996 3572 365002 3636
rect 136449 3498 136515 3501
rect 365110 3498 365116 3500
rect 136449 3496 365116 3498
rect 136449 3440 136454 3496
rect 136510 3440 365116 3496
rect 136449 3438 365116 3440
rect 136449 3435 136515 3438
rect 365110 3436 365116 3438
rect 365180 3436 365186 3500
rect 132953 3362 133019 3365
rect 367686 3362 367692 3364
rect 132953 3360 367692 3362
rect 132953 3304 132958 3360
rect 133014 3304 367692 3360
rect 132953 3302 367692 3304
rect 132953 3299 133019 3302
rect 367686 3300 367692 3302
rect 367756 3300 367762 3364
rect 143533 3226 143599 3229
rect 206134 3226 206140 3228
rect 143533 3224 206140 3226
rect 143533 3168 143538 3224
rect 143594 3168 206140 3224
rect 143533 3166 206140 3168
rect 143533 3163 143599 3166
rect 206134 3164 206140 3166
rect 206204 3164 206210 3228
rect 365713 3226 365779 3229
rect 366950 3226 366956 3228
rect 365713 3224 366956 3226
rect 365713 3168 365718 3224
rect 365774 3168 366956 3224
rect 365713 3166 366956 3168
rect 365713 3163 365779 3166
rect 366950 3164 366956 3166
rect 367020 3164 367026 3228
<< via3 >>
rect 54340 639372 54404 639436
rect 476068 634884 476132 634948
rect 488580 634884 488644 634948
rect 506612 634884 506676 634948
rect 436140 611356 436204 611420
rect 436324 606596 436388 606660
rect 436508 586468 436572 586532
rect 324820 549476 324884 549540
rect 324820 529484 324884 529548
rect 436324 528396 436388 528460
rect 436508 528260 436572 528324
rect 436140 528124 436204 528188
rect 363460 523636 363524 523700
rect 360700 518060 360764 518124
rect 367692 489092 367756 489156
rect 476068 489092 476132 489156
rect 364932 487732 364996 487796
rect 365116 486508 365180 486572
rect 206140 486372 206204 486436
rect 488580 486372 488644 486436
rect 59308 485692 59372 485756
rect 55076 485556 55140 485620
rect 55628 485420 55692 485484
rect 199332 485692 199396 485756
rect 198044 485556 198108 485620
rect 357940 485556 358004 485620
rect 196572 485420 196636 485484
rect 213684 485420 213748 485484
rect 367876 485420 367940 485484
rect 51948 485284 52012 485348
rect 197860 485284 197924 485348
rect 201356 485284 201420 485348
rect 209636 485284 209700 485348
rect 211660 485284 211724 485348
rect 371740 485284 371804 485348
rect 53236 485148 53300 485212
rect 200804 485148 200868 485212
rect 202644 485148 202708 485212
rect 205220 485148 205284 485212
rect 375972 485148 376036 485212
rect 57836 485012 57900 485076
rect 200620 485012 200684 485076
rect 216996 485012 217060 485076
rect 219204 485012 219268 485076
rect 374684 485012 374748 485076
rect 59124 484876 59188 484940
rect 196756 484876 196820 484940
rect 198412 484876 198476 484940
rect 205404 484876 205468 484940
rect 198596 484740 198660 484804
rect 206692 484740 206756 484804
rect 212396 484740 212460 484804
rect 50292 484468 50356 484532
rect 50844 484528 50908 484532
rect 50844 484472 50894 484528
rect 50894 484472 50908 484528
rect 50844 484468 50908 484472
rect 217548 484468 217612 484532
rect 219940 484468 220004 484532
rect 213868 483788 213932 483852
rect 370452 483788 370516 483852
rect 214604 483652 214668 483716
rect 374500 483652 374564 483716
rect 46796 482700 46860 482764
rect 57100 482564 57164 482628
rect 359412 482428 359476 482492
rect 215340 482292 215404 482356
rect 375420 482292 375484 482356
rect 202460 480932 202524 480996
rect 214052 480796 214116 480860
rect 370084 480796 370148 480860
rect 57652 479844 57716 479908
rect 217180 479708 217244 479772
rect 359596 479708 359660 479772
rect 215892 479572 215956 479636
rect 378732 479572 378796 479636
rect 208348 479436 208412 479500
rect 210372 479436 210436 479500
rect 213316 478348 213380 478412
rect 210556 478212 210620 478276
rect 358124 478212 358188 478276
rect 213132 478076 213196 478140
rect 379468 478076 379532 478140
rect 57468 477260 57532 477324
rect 44772 477124 44836 477188
rect 44956 476988 45020 477052
rect 209820 476852 209884 476916
rect 214420 476716 214484 476780
rect 378180 476716 378244 476780
rect 359780 475628 359844 475692
rect 218652 475492 218716 475556
rect 360148 475492 360212 475556
rect 202092 475356 202156 475420
rect 207060 474132 207124 474196
rect 216076 473996 216140 474060
rect 378916 473996 378980 474060
rect 377260 472908 377324 472972
rect 216260 472772 216324 472836
rect 366956 472772 367020 472836
rect 506612 472772 506676 472836
rect 202276 472636 202340 472700
rect 371924 472636 371988 472700
rect 203196 472500 203260 472564
rect 379100 472500 379164 472564
rect 199516 471684 199580 471748
rect 204852 471548 204916 471612
rect 217364 471412 217428 471476
rect 377444 471276 377508 471340
rect 377628 471140 377692 471204
rect 47900 469780 47964 469844
rect 60228 469100 60292 469164
rect 48084 468964 48148 469028
rect 206324 468964 206388 469028
rect 46612 468828 46676 468892
rect 205036 468828 205100 468892
rect 55444 468692 55508 468756
rect 200988 468692 201052 468756
rect 53604 468556 53668 468620
rect 206508 468556 206572 468620
rect 50476 468420 50540 468484
rect 213500 468420 213564 468484
rect 377812 468420 377876 468484
rect 58940 468284 59004 468348
rect 48636 467876 48700 467940
rect 50660 467936 50724 467940
rect 50660 467880 50710 467936
rect 50710 467880 50724 467936
rect 50660 467876 50724 467880
rect 208900 467196 208964 467260
rect 218836 467060 218900 467124
rect 179644 466924 179708 466988
rect 178356 466516 178420 466580
rect 190868 466576 190932 466580
rect 190868 466520 190918 466576
rect 190918 466520 190932 466576
rect 190868 466516 190932 466520
rect 338436 466576 338500 466580
rect 338436 466520 338486 466576
rect 338486 466520 338500 466576
rect 338436 466516 338500 466520
rect 339724 466576 339788 466580
rect 339724 466520 339774 466576
rect 339774 466520 339788 466576
rect 339724 466516 339788 466520
rect 350948 466576 351012 466580
rect 350948 466520 350998 466576
rect 350998 466520 351012 466576
rect 350948 466516 351012 466520
rect 498516 466576 498580 466580
rect 498516 466520 498530 466576
rect 498530 466520 498580 466576
rect 498516 466516 498580 466520
rect 499804 466576 499868 466580
rect 499804 466520 499818 466576
rect 499818 466520 499868 466576
rect 499804 466516 499868 466520
rect 510844 466576 510908 466580
rect 510844 466520 510894 466576
rect 510894 466520 510908 466576
rect 510844 466516 510908 466520
rect 58572 466380 58636 466444
rect 54892 466244 54956 466308
rect 53420 466108 53484 466172
rect 198780 466108 198844 466172
rect 54708 465972 54772 466036
rect 51580 465836 51644 465900
rect 53052 465836 53116 465900
rect 207980 465836 208044 465900
rect 359964 465836 360028 465900
rect 52132 465700 52196 465764
rect 370636 465700 370700 465764
rect 58756 465564 58820 465628
rect 51764 465156 51828 465220
rect 199148 464340 199212 464404
rect 206692 415244 206756 415308
rect 53052 388452 53116 388516
rect 57468 388452 57532 388516
rect 377444 382332 377508 382396
rect 199148 381516 199212 381580
rect 248294 380836 248358 380900
rect 359780 380836 359844 380900
rect 428286 380836 428350 380900
rect 431142 380896 431206 380900
rect 431142 380840 431186 380896
rect 431186 380840 431206 380896
rect 431142 380836 431206 380840
rect 433590 380896 433654 380900
rect 433590 380840 433614 380896
rect 433614 380840 433654 380896
rect 433590 380836 433654 380840
rect 438486 380896 438550 380900
rect 438486 380840 438490 380896
rect 438490 380840 438546 380896
rect 438546 380840 438550 380896
rect 438486 380836 438550 380840
rect 111006 380760 111070 380764
rect 111006 380704 111026 380760
rect 111026 380704 111070 380760
rect 111006 380700 111070 380704
rect 113590 380760 113654 380764
rect 113590 380704 113602 380760
rect 113602 380704 113654 380760
rect 113590 380700 113654 380704
rect 116038 380760 116102 380764
rect 116038 380704 116086 380760
rect 116086 380704 116102 380760
rect 116038 380700 116102 380704
rect 118486 380700 118550 380764
rect 120934 380700 120998 380764
rect 123518 380760 123582 380764
rect 123518 380704 123538 380760
rect 123538 380704 123582 380760
rect 123518 380700 123582 380704
rect 125966 380760 126030 380764
rect 125966 380704 126022 380760
rect 126022 380704 126030 380760
rect 125966 380700 126030 380704
rect 130998 380760 131062 380764
rect 130998 380704 131026 380760
rect 131026 380704 131062 380760
rect 130998 380700 131062 380704
rect 133446 380700 133510 380764
rect 140926 380760 140990 380764
rect 140926 380704 140962 380760
rect 140962 380704 140990 380760
rect 140926 380700 140990 380704
rect 143510 380760 143574 380764
rect 143510 380704 143538 380760
rect 143538 380704 143574 380760
rect 143510 380700 143574 380704
rect 145958 380700 146022 380764
rect 155886 380700 155950 380764
rect 158470 380700 158534 380764
rect 160918 380760 160982 380764
rect 160918 380704 160926 380760
rect 160926 380704 160982 380760
rect 160918 380700 160982 380704
rect 163366 380760 163430 380764
rect 163366 380704 163410 380760
rect 163410 380704 163430 380760
rect 163366 380700 163430 380704
rect 165950 380760 166014 380764
rect 165950 380704 165986 380760
rect 165986 380704 166014 380760
rect 165950 380700 166014 380704
rect 202644 380700 202708 380764
rect 205220 380760 205284 380764
rect 205220 380704 205234 380760
rect 205234 380704 205284 380760
rect 205220 380700 205284 380704
rect 279166 380700 279230 380764
rect 410742 380760 410806 380764
rect 410742 380704 410762 380760
rect 410762 380704 410806 380760
rect 410742 380700 410806 380704
rect 421078 380760 421142 380764
rect 421078 380704 421102 380760
rect 421102 380704 421142 380760
rect 421078 380700 421142 380704
rect 436038 380760 436102 380764
rect 436038 380704 436062 380760
rect 436062 380704 436102 380760
rect 436038 380700 436102 380704
rect 440934 380760 440998 380764
rect 440934 380704 440938 380760
rect 440938 380704 440998 380760
rect 440934 380700 440998 380704
rect 443518 380700 443582 380764
rect 236054 380564 236118 380628
rect 237142 380624 237206 380628
rect 237142 380568 237158 380624
rect 237158 380568 237206 380624
rect 237142 380564 237206 380568
rect 243126 380624 243190 380628
rect 243126 380568 243138 380624
rect 243138 380568 243190 380624
rect 243126 380564 243190 380568
rect 245438 380564 245502 380628
rect 247614 380624 247678 380628
rect 247614 380568 247646 380624
rect 247646 380568 247678 380624
rect 247614 380564 247678 380568
rect 254550 380564 254614 380628
rect 255910 380624 255974 380628
rect 255910 380568 255926 380624
rect 255926 380568 255974 380624
rect 255910 380564 255974 380568
rect 256998 380624 257062 380628
rect 256998 380568 257030 380624
rect 257030 380568 257062 380624
rect 256998 380564 257062 380568
rect 258086 380624 258150 380628
rect 258086 380568 258134 380624
rect 258134 380568 258150 380624
rect 258086 380564 258150 380568
rect 259446 380624 259510 380628
rect 259446 380568 259458 380624
rect 259458 380568 259510 380624
rect 259446 380564 259510 380568
rect 260670 380564 260734 380628
rect 265294 380624 265358 380628
rect 265294 380568 265310 380624
rect 265310 380568 265358 380624
rect 265294 380564 265358 380568
rect 76052 380428 76116 380492
rect 217916 380428 217980 380492
rect 269782 380564 269846 380628
rect 271006 380624 271070 380628
rect 271006 380568 271014 380624
rect 271014 380568 271070 380624
rect 271006 380564 271070 380568
rect 405438 380624 405502 380628
rect 405438 380568 405462 380624
rect 405462 380568 405502 380624
rect 405438 380564 405502 380568
rect 413462 380624 413526 380628
rect 413462 380568 413466 380624
rect 413466 380568 413522 380624
rect 413522 380568 413526 380624
rect 413462 380564 413526 380568
rect 419446 380624 419510 380628
rect 419446 380568 419502 380624
rect 419502 380568 419510 380624
rect 419446 380564 419510 380568
rect 434406 380564 434470 380628
rect 485950 380624 486014 380628
rect 485950 380568 485962 380624
rect 485962 380568 486014 380624
rect 485950 380564 486014 380568
rect 426388 380488 426452 380492
rect 426388 380432 426438 380488
rect 426438 380432 426452 380488
rect 426388 380428 426452 380432
rect 119108 380292 119172 380356
rect 216996 380292 217060 380356
rect 323348 380292 323412 380356
rect 128308 380216 128372 380220
rect 128308 380160 128358 380216
rect 128358 380160 128372 380216
rect 128308 380156 128372 380160
rect 216628 380156 216692 380220
rect 217548 380156 217612 380220
rect 279188 380156 279252 380220
rect 359596 380156 359660 380220
rect 404124 380156 404188 380220
rect 50292 379476 50356 379540
rect 51948 379476 52012 379540
rect 208348 379476 208412 379540
rect 81756 379340 81820 379404
rect 81940 379340 82004 379404
rect 85436 379400 85500 379404
rect 85436 379344 85486 379400
rect 85486 379344 85500 379400
rect 85436 379340 85500 379344
rect 86540 379400 86604 379404
rect 86540 379344 86590 379400
rect 86590 379344 86604 379400
rect 86540 379340 86604 379344
rect 87644 379340 87708 379404
rect 88380 379400 88444 379404
rect 88380 379344 88394 379400
rect 88394 379344 88444 379400
rect 88380 379340 88444 379344
rect 88748 379400 88812 379404
rect 88748 379344 88798 379400
rect 88798 379344 88812 379400
rect 88748 379340 88812 379344
rect 90036 379400 90100 379404
rect 90036 379344 90086 379400
rect 90086 379344 90100 379400
rect 90036 379340 90100 379344
rect 90772 379340 90836 379404
rect 91324 379400 91388 379404
rect 91324 379344 91374 379400
rect 91374 379344 91388 379400
rect 91324 379340 91388 379344
rect 92428 379400 92492 379404
rect 92428 379344 92442 379400
rect 92442 379344 92492 379400
rect 92428 379340 92492 379344
rect 93348 379340 93412 379404
rect 96108 379400 96172 379404
rect 96108 379344 96122 379400
rect 96122 379344 96172 379400
rect 96108 379340 96172 379344
rect 98132 379340 98196 379404
rect 98500 379400 98564 379404
rect 98500 379344 98514 379400
rect 98514 379344 98564 379400
rect 98500 379340 98564 379344
rect 101076 379400 101140 379404
rect 101076 379344 101090 379400
rect 101090 379344 101140 379400
rect 101076 379340 101140 379344
rect 103284 379340 103348 379404
rect 105860 379340 105924 379404
rect 108252 379400 108316 379404
rect 108252 379344 108266 379400
rect 108266 379344 108316 379400
rect 108252 379340 108316 379344
rect 108804 379400 108868 379404
rect 108804 379344 108854 379400
rect 108854 379344 108868 379400
rect 108804 379340 108868 379344
rect 111196 379340 111260 379404
rect 112300 379400 112364 379404
rect 112300 379344 112350 379400
rect 112350 379344 112364 379400
rect 112300 379340 112364 379344
rect 113404 379400 113468 379404
rect 113404 379344 113454 379400
rect 113454 379344 113468 379400
rect 113404 379340 113468 379344
rect 114508 379400 114572 379404
rect 114508 379344 114522 379400
rect 114522 379344 114572 379400
rect 114508 379340 114572 379344
rect 115796 379400 115860 379404
rect 115796 379344 115846 379400
rect 115846 379344 115860 379400
rect 115796 379340 115860 379344
rect 135852 379400 135916 379404
rect 135852 379344 135902 379400
rect 135902 379344 135916 379400
rect 135852 379340 135916 379344
rect 138428 379400 138492 379404
rect 138428 379344 138478 379400
rect 138478 379344 138492 379400
rect 138428 379340 138492 379344
rect 150940 379400 151004 379404
rect 150940 379344 150990 379400
rect 150990 379344 151004 379400
rect 150940 379340 151004 379344
rect 153516 379340 153580 379404
rect 57100 379068 57164 379132
rect 80468 379264 80532 379268
rect 80468 379208 80482 379264
rect 80482 379208 80532 379264
rect 80468 379204 80532 379208
rect 93716 379204 93780 379268
rect 95924 379264 95988 379268
rect 95924 379208 95974 379264
rect 95974 379208 95988 379264
rect 95924 379204 95988 379208
rect 99420 379264 99484 379268
rect 99420 379208 99470 379264
rect 99470 379208 99484 379264
rect 99420 379204 99484 379208
rect 102916 379264 102980 379268
rect 102916 379208 102966 379264
rect 102966 379208 102980 379264
rect 102916 379204 102980 379208
rect 109724 379204 109788 379268
rect 246436 379340 246500 379404
rect 248644 379400 248708 379404
rect 248644 379344 248658 379400
rect 248658 379344 248708 379400
rect 248644 379340 248708 379344
rect 250116 379400 250180 379404
rect 250116 379344 250130 379400
rect 250130 379344 250180 379400
rect 250116 379340 250180 379344
rect 251220 379400 251284 379404
rect 251220 379344 251234 379400
rect 251234 379344 251284 379400
rect 251220 379340 251284 379344
rect 252324 379400 252388 379404
rect 252324 379344 252338 379400
rect 252338 379344 252388 379400
rect 252324 379340 252388 379344
rect 253428 379400 253492 379404
rect 253428 379344 253442 379400
rect 253442 379344 253492 379400
rect 253428 379340 253492 379344
rect 261708 379400 261772 379404
rect 261708 379344 261722 379400
rect 261722 379344 261772 379400
rect 261708 379340 261772 379344
rect 263916 379400 263980 379404
rect 263916 379344 263930 379400
rect 263930 379344 263980 379400
rect 263916 379340 263980 379344
rect 268700 379400 268764 379404
rect 268700 379344 268714 379400
rect 268714 379344 268764 379400
rect 268700 379340 268764 379344
rect 271092 379400 271156 379404
rect 271092 379344 271106 379400
rect 271106 379344 271156 379400
rect 271092 379340 271156 379344
rect 272196 379400 272260 379404
rect 272196 379344 272210 379400
rect 272210 379344 272260 379400
rect 272196 379340 272260 379344
rect 273300 379400 273364 379404
rect 273300 379344 273314 379400
rect 273314 379344 273364 379400
rect 273300 379340 273364 379344
rect 274404 379400 274468 379404
rect 274404 379344 274418 379400
rect 274418 379344 274468 379400
rect 274404 379340 274468 379344
rect 275692 379400 275756 379404
rect 275692 379344 275706 379400
rect 275706 379344 275756 379400
rect 275692 379340 275756 379344
rect 276060 379400 276124 379404
rect 276060 379344 276110 379400
rect 276110 379344 276124 379400
rect 276060 379340 276124 379344
rect 276980 379400 277044 379404
rect 276980 379344 277030 379400
rect 277030 379344 277044 379400
rect 276980 379340 277044 379344
rect 278452 379340 278516 379404
rect 285996 379400 286060 379404
rect 285996 379344 286010 379400
rect 286010 379344 286060 379400
rect 285996 379340 286060 379344
rect 288204 379340 288268 379404
rect 290964 379400 291028 379404
rect 290964 379344 290978 379400
rect 290978 379344 291028 379400
rect 290964 379340 291028 379344
rect 293356 379340 293420 379404
rect 295932 379340 295996 379404
rect 298508 379400 298572 379404
rect 298508 379344 298522 379400
rect 298522 379344 298572 379400
rect 298508 379340 298572 379344
rect 300900 379400 300964 379404
rect 300900 379344 300914 379400
rect 300914 379344 300964 379400
rect 300900 379340 300964 379344
rect 303476 379340 303540 379404
rect 305868 379400 305932 379404
rect 305868 379344 305882 379400
rect 305882 379344 305932 379400
rect 305868 379340 305932 379344
rect 308444 379340 308508 379404
rect 311020 379400 311084 379404
rect 311020 379344 311034 379400
rect 311034 379344 311084 379400
rect 311020 379340 311084 379344
rect 313412 379400 313476 379404
rect 313412 379344 313426 379400
rect 313426 379344 313476 379400
rect 313412 379340 313476 379344
rect 315804 379400 315868 379404
rect 315804 379344 315818 379400
rect 315818 379344 315868 379400
rect 315804 379340 315868 379344
rect 318380 379340 318444 379404
rect 396028 379400 396092 379404
rect 396028 379344 396078 379400
rect 396078 379344 396092 379400
rect 396028 379340 396092 379344
rect 397132 379400 397196 379404
rect 397132 379344 397146 379400
rect 397146 379344 397196 379400
rect 397132 379340 397196 379344
rect 278084 379204 278148 379268
rect 280844 379204 280908 379268
rect 283420 379264 283484 379268
rect 283420 379208 283434 379264
rect 283434 379208 283484 379264
rect 283420 379204 283484 379208
rect 325924 379264 325988 379268
rect 401732 379340 401796 379404
rect 406516 379340 406580 379404
rect 407620 379400 407684 379404
rect 407620 379344 407634 379400
rect 407634 379344 407684 379400
rect 407620 379340 407684 379344
rect 408356 379400 408420 379404
rect 408356 379344 408370 379400
rect 408370 379344 408420 379400
rect 408356 379340 408420 379344
rect 411300 379400 411364 379404
rect 411300 379344 411314 379400
rect 411314 379344 411364 379400
rect 411300 379340 411364 379344
rect 412404 379400 412468 379404
rect 412404 379344 412418 379400
rect 412418 379344 412468 379400
rect 412404 379340 412468 379344
rect 416084 379340 416148 379404
rect 426020 379400 426084 379404
rect 426020 379344 426034 379400
rect 426034 379344 426084 379400
rect 426020 379340 426084 379344
rect 435772 379340 435836 379404
rect 437980 379340 438044 379404
rect 445892 379400 445956 379404
rect 445892 379344 445906 379400
rect 445906 379344 445956 379400
rect 445892 379340 445956 379344
rect 448284 379340 448348 379404
rect 451044 379400 451108 379404
rect 451044 379344 451058 379400
rect 451058 379344 451108 379400
rect 451044 379340 451108 379344
rect 453436 379340 453500 379404
rect 455828 379340 455892 379404
rect 458404 379400 458468 379404
rect 458404 379344 458418 379400
rect 458418 379344 458468 379400
rect 458404 379340 458468 379344
rect 460980 379400 461044 379404
rect 460980 379344 460994 379400
rect 460994 379344 461044 379400
rect 460980 379340 461044 379344
rect 475884 379340 475948 379404
rect 325924 379208 325938 379264
rect 325938 379208 325988 379264
rect 325924 379204 325988 379208
rect 78260 379068 78324 379132
rect 77156 378992 77220 378996
rect 77156 378936 77206 378992
rect 77206 378936 77220 378992
rect 77156 378932 77220 378936
rect 94636 378992 94700 378996
rect 94636 378936 94686 378992
rect 94686 378936 94700 378992
rect 79548 378796 79612 378860
rect 83228 378856 83292 378860
rect 83228 378800 83278 378856
rect 83278 378800 83292 378856
rect 83228 378796 83292 378800
rect 94636 378932 94700 378936
rect 148548 378932 148612 378996
rect 183140 378932 183204 378996
rect 241836 379068 241900 379132
rect 398236 379204 398300 379268
rect 399524 379264 399588 379268
rect 399524 379208 399538 379264
rect 399538 379208 399588 379264
rect 399524 379204 399588 379208
rect 400444 379264 400508 379268
rect 400444 379208 400458 379264
rect 400458 379208 400508 379264
rect 400444 379204 400508 379208
rect 403020 379264 403084 379268
rect 403020 379208 403034 379264
rect 403034 379208 403084 379264
rect 403020 379204 403084 379208
rect 410012 379264 410076 379268
rect 410012 379208 410026 379264
rect 410026 379208 410076 379264
rect 410012 379204 410076 379208
rect 415900 379264 415964 379268
rect 415900 379208 415914 379264
rect 415914 379208 415964 379264
rect 415900 379204 415964 379208
rect 238156 378932 238220 378996
rect 417004 379204 417068 379268
rect 423444 379204 423508 379268
rect 463556 379264 463620 379268
rect 463556 379208 463570 379264
rect 463570 379208 463620 379264
rect 463556 379204 463620 379208
rect 473492 379264 473556 379268
rect 473492 379208 473506 379264
rect 473506 379208 473556 379264
rect 473492 379204 473556 379208
rect 503116 379264 503180 379268
rect 503116 379208 503130 379264
rect 503130 379208 503180 379264
rect 503116 379204 503180 379208
rect 503484 379264 503548 379268
rect 503484 379208 503534 379264
rect 503534 379208 503548 379264
rect 503484 379204 503548 379208
rect 465948 378932 466012 378996
rect 478460 378932 478524 378996
rect 239260 378796 239324 378860
rect 377628 378796 377692 378860
rect 427676 378796 427740 378860
rect 430988 378796 431052 378860
rect 470916 378796 470980 378860
rect 483428 378856 483492 378860
rect 483428 378800 483442 378856
rect 483442 378800 483492 378856
rect 483428 378796 483492 378800
rect 81940 378660 82004 378724
rect 209820 378660 209884 378724
rect 241468 378660 241532 378724
rect 377812 378660 377876 378724
rect 433380 378660 433444 378724
rect 436876 378660 436940 378724
rect 468524 378660 468588 378724
rect 97028 378524 97092 378588
rect 100708 378524 100772 378588
rect 118188 378524 118252 378588
rect 105308 378388 105372 378452
rect 183508 378388 183572 378452
rect 205404 378448 205468 378452
rect 205404 378392 205418 378448
rect 205418 378392 205468 378448
rect 205404 378388 205468 378392
rect 241836 378388 241900 378452
rect 253612 378584 253676 378588
rect 253612 378528 253626 378584
rect 253626 378528 253676 378584
rect 253612 378524 253676 378528
rect 256004 378584 256068 378588
rect 256004 378528 256018 378584
rect 256018 378528 256068 378584
rect 256004 378524 256068 378528
rect 258396 378584 258460 378588
rect 258396 378528 258410 378584
rect 258410 378528 258460 378584
rect 258396 378524 258460 378528
rect 260972 378584 261036 378588
rect 260972 378528 260986 378584
rect 260986 378528 261036 378584
rect 260972 378524 261036 378528
rect 263548 378584 263612 378588
rect 263548 378528 263598 378584
rect 263598 378528 263612 378584
rect 263548 378524 263612 378528
rect 265940 378584 266004 378588
rect 265940 378528 265954 378584
rect 265954 378528 266004 378584
rect 265940 378524 266004 378528
rect 268332 378524 268396 378588
rect 273484 378584 273548 378588
rect 273484 378528 273498 378584
rect 273498 378528 273548 378584
rect 273484 378524 273548 378528
rect 320956 378584 321020 378588
rect 320956 378528 320970 378584
rect 320970 378528 321020 378584
rect 320956 378524 321020 378528
rect 413508 378524 413572 378588
rect 414612 378584 414676 378588
rect 414612 378528 414626 378584
rect 414626 378528 414676 378584
rect 414612 378524 414676 378528
rect 418476 378584 418540 378588
rect 418476 378528 418490 378584
rect 418490 378528 418540 378584
rect 418476 378524 418540 378528
rect 343220 378448 343284 378452
rect 343220 378392 343234 378448
rect 343234 378392 343284 378448
rect 343220 378388 343284 378392
rect 240548 378252 240612 378316
rect 241468 378252 241532 378316
rect 244228 378312 244292 378316
rect 244228 378256 244278 378312
rect 244278 378256 244292 378312
rect 244228 378252 244292 378256
rect 250668 378312 250732 378316
rect 250668 378256 250682 378312
rect 250682 378256 250732 378312
rect 250668 378252 250732 378256
rect 262812 378312 262876 378316
rect 262812 378256 262826 378312
rect 262826 378256 262876 378312
rect 262812 378252 262876 378256
rect 266308 378312 266372 378316
rect 266308 378256 266358 378312
rect 266358 378256 266372 378312
rect 266308 378252 266372 378256
rect 267596 378312 267660 378316
rect 267596 378256 267610 378312
rect 267610 378256 267660 378312
rect 267596 378252 267660 378256
rect 343404 378252 343468 378316
rect 432276 378312 432340 378316
rect 432276 378256 432290 378312
rect 432290 378256 432340 378312
rect 432276 378252 432340 378256
rect 84332 378176 84396 378180
rect 84332 378120 84382 378176
rect 84382 378120 84396 378176
rect 84332 378116 84396 378120
rect 101812 378176 101876 378180
rect 101812 378120 101862 378176
rect 101862 378120 101876 378176
rect 101812 378116 101876 378120
rect 104020 378116 104084 378180
rect 106412 378176 106476 378180
rect 106412 378120 106462 378176
rect 106462 378120 106476 378176
rect 106412 378116 106476 378120
rect 107516 378176 107580 378180
rect 107516 378120 107566 378176
rect 107566 378120 107580 378176
rect 107516 378116 107580 378120
rect 117084 378116 117148 378180
rect 57468 377980 57532 378044
rect 377444 378176 377508 378180
rect 377444 378120 377458 378176
rect 377458 378120 377508 378176
rect 377444 378116 377508 378120
rect 408724 378176 408788 378180
rect 408724 378120 408738 378176
rect 408738 378120 408788 378176
rect 408724 378116 408788 378120
rect 418108 378176 418172 378180
rect 418108 378120 418158 378176
rect 418158 378120 418172 378176
rect 418108 378116 418172 378120
rect 420684 378176 420748 378180
rect 420684 378120 420698 378176
rect 420698 378120 420748 378176
rect 420684 378116 420748 378120
rect 421788 378116 421852 378180
rect 422892 378116 422956 378180
rect 423996 378176 424060 378180
rect 423996 378120 424010 378176
rect 424010 378120 424060 378176
rect 423996 378116 424060 378120
rect 425284 378116 425348 378180
rect 428596 378176 428660 378180
rect 428596 378120 428610 378176
rect 428610 378120 428660 378176
rect 428596 378116 428660 378120
rect 429700 378176 429764 378180
rect 429700 378120 429714 378176
rect 429714 378120 429764 378176
rect 429700 378116 429764 378120
rect 439084 378176 439148 378180
rect 439084 378120 439098 378176
rect 439098 378120 439148 378176
rect 439084 378116 439148 378120
rect 207060 377980 207124 378044
rect 211660 377980 211724 378044
rect 213684 377980 213748 378044
rect 214052 377980 214116 378044
rect 360148 377980 360212 378044
rect 480668 378116 480732 378180
rect 370084 377844 370148 377908
rect 213868 376620 213932 376684
rect 359964 376620 360028 376684
rect 216628 376484 216692 376548
rect 216996 375940 217060 376004
rect 215340 375396 215404 375460
rect 376708 374912 376772 374916
rect 376708 374856 376758 374912
rect 376758 374856 376772 374912
rect 376708 374852 376772 374856
rect 178540 358864 178604 358868
rect 178540 358808 178590 358864
rect 178590 358808 178604 358864
rect 178540 358804 178604 358808
rect 179644 358804 179708 358868
rect 190868 358864 190932 358868
rect 190868 358808 190918 358864
rect 190918 358808 190932 358864
rect 190868 358804 190932 358808
rect 338436 358864 338500 358868
rect 338436 358808 338486 358864
rect 338486 358808 338500 358864
rect 338436 358804 338500 358808
rect 339724 358804 339788 358868
rect 350948 358804 351012 358868
rect 498516 358804 498580 358868
rect 499804 358804 499868 358868
rect 510844 358864 510908 358868
rect 510844 358808 510894 358864
rect 510894 358808 510908 358864
rect 510844 358804 510908 358808
rect 377996 357308 378060 357372
rect 51580 282236 51644 282300
rect 113318 273864 113382 273868
rect 113318 273808 113362 273864
rect 113362 273808 113382 273864
rect 113318 273804 113382 273808
rect 426382 273864 426446 273868
rect 426382 273808 426438 273864
rect 426438 273808 426446 273864
rect 426382 273804 426446 273808
rect 133446 273728 133510 273732
rect 133446 273672 133474 273728
rect 133474 273672 133510 273728
rect 133446 273668 133510 273672
rect 135894 273592 135958 273596
rect 135894 273536 135902 273592
rect 135902 273536 135958 273592
rect 135894 273532 135958 273536
rect 138478 273592 138542 273596
rect 138478 273536 138534 273592
rect 138534 273536 138542 273592
rect 138478 273532 138542 273536
rect 140926 273532 140990 273596
rect 143510 273592 143574 273596
rect 143510 273536 143538 273592
rect 143538 273536 143574 273592
rect 143510 273532 143574 273536
rect 145958 273592 146022 273596
rect 145958 273536 145986 273592
rect 145986 273536 146022 273592
rect 145958 273532 146022 273536
rect 266382 273592 266446 273596
rect 266382 273536 266414 273592
rect 266414 273536 266446 273592
rect 266382 273532 266446 273536
rect 283518 273592 283582 273596
rect 283518 273536 283526 273592
rect 283526 273536 283582 273592
rect 283518 273532 283582 273536
rect 421078 273592 421142 273596
rect 421078 273536 421102 273592
rect 421102 273536 421142 273592
rect 421078 273532 421142 273536
rect 431142 273592 431206 273596
rect 431142 273536 431186 273592
rect 431186 273536 431206 273592
rect 431142 273532 431206 273536
rect 433318 273592 433382 273596
rect 433318 273536 433338 273592
rect 433338 273536 433382 273592
rect 433318 273532 433382 273536
rect 453446 273592 453510 273596
rect 453446 273536 453450 273592
rect 453450 273536 453510 273592
rect 453446 273532 453510 273536
rect 218836 273396 218900 273460
rect 273300 273456 273364 273460
rect 273300 273400 273314 273456
rect 273314 273400 273364 273456
rect 273300 273396 273364 273400
rect 430988 273456 431052 273460
rect 430988 273400 431002 273456
rect 431002 273400 431052 273456
rect 430988 273396 431052 273400
rect 57468 273260 57532 273324
rect 199516 273260 199580 273324
rect 250668 273260 250732 273324
rect 376892 273260 376956 273324
rect 377812 273260 377876 273324
rect 378180 273260 378244 273324
rect 76052 273184 76116 273188
rect 76052 273128 76066 273184
rect 76066 273128 76116 273184
rect 76052 273124 76116 273128
rect 77156 273184 77220 273188
rect 77156 273128 77170 273184
rect 77170 273128 77220 273184
rect 77156 273124 77220 273128
rect 83044 273184 83108 273188
rect 83044 273128 83058 273184
rect 83058 273128 83108 273184
rect 83044 273124 83108 273128
rect 90772 273184 90836 273188
rect 90772 273128 90786 273184
rect 90786 273128 90836 273184
rect 90772 273124 90836 273128
rect 93716 273184 93780 273188
rect 93716 273128 93730 273184
rect 93730 273128 93780 273184
rect 93716 273124 93780 273128
rect 95924 273184 95988 273188
rect 95924 273128 95938 273184
rect 95938 273128 95988 273184
rect 95924 273124 95988 273128
rect 101812 273124 101876 273188
rect 199332 273124 199396 273188
rect 318380 273124 318444 273188
rect 359412 273124 359476 273188
rect 422892 273184 422956 273188
rect 422892 273128 422906 273184
rect 422906 273128 422956 273184
rect 422892 273124 422956 273128
rect 423444 273184 423508 273188
rect 423444 273128 423458 273184
rect 423458 273128 423508 273184
rect 423444 273124 423508 273128
rect 426020 273184 426084 273188
rect 426020 273128 426034 273184
rect 426034 273128 426084 273184
rect 426020 273124 426084 273128
rect 102732 272988 102796 273052
rect 196756 272988 196820 273052
rect 311020 272988 311084 273052
rect 377812 272988 377876 273052
rect 425284 272988 425348 273052
rect 468524 273048 468588 273052
rect 468524 272992 468538 273048
rect 468538 272992 468588 273048
rect 468524 272988 468588 272992
rect 470916 273048 470980 273052
rect 470916 272992 470930 273048
rect 470930 272992 470980 273048
rect 470916 272988 470980 272992
rect 103836 272852 103900 272916
rect 217364 272852 217428 272916
rect 285996 272912 286060 272916
rect 285996 272856 286010 272912
rect 286010 272856 286060 272912
rect 96108 272776 96172 272780
rect 96108 272720 96122 272776
rect 96122 272720 96172 272776
rect 96108 272716 96172 272720
rect 98500 272776 98564 272780
rect 98500 272720 98514 272776
rect 98514 272720 98564 272776
rect 98500 272716 98564 272720
rect 285996 272852 286060 272856
rect 288204 272912 288268 272916
rect 288204 272856 288218 272912
rect 288218 272856 288268 272912
rect 288204 272852 288268 272856
rect 290964 272912 291028 272916
rect 290964 272856 290978 272912
rect 290978 272856 291028 272912
rect 290964 272852 291028 272856
rect 295932 272912 295996 272916
rect 295932 272856 295946 272912
rect 295946 272856 295996 272912
rect 295932 272852 295996 272856
rect 303476 272912 303540 272916
rect 303476 272856 303490 272912
rect 303490 272856 303540 272912
rect 303476 272852 303540 272856
rect 428228 272852 428292 272916
rect 473492 272912 473556 272916
rect 473492 272856 473506 272912
rect 473506 272856 473556 272912
rect 473492 272852 473556 272856
rect 475884 272912 475948 272916
rect 475884 272856 475898 272912
rect 475898 272856 475948 272912
rect 475884 272852 475948 272856
rect 293356 272716 293420 272780
rect 298508 272776 298572 272780
rect 298508 272720 298522 272776
rect 298522 272720 298572 272776
rect 298508 272716 298572 272720
rect 300900 272776 300964 272780
rect 300900 272720 300914 272776
rect 300914 272720 300964 272776
rect 300900 272716 300964 272720
rect 478460 272776 478524 272780
rect 478460 272720 478474 272776
rect 478474 272720 478524 272776
rect 478460 272716 478524 272720
rect 480852 272776 480916 272780
rect 480852 272720 480866 272776
rect 480866 272720 480916 272776
rect 480852 272716 480916 272720
rect 116900 272580 116964 272644
rect 305868 272640 305932 272644
rect 305868 272584 305882 272640
rect 305882 272584 305932 272640
rect 305868 272580 305932 272584
rect 320956 272640 321020 272644
rect 320956 272584 320970 272640
rect 320970 272584 321020 272640
rect 320956 272580 321020 272584
rect 377996 272580 378060 272644
rect 483244 272640 483308 272644
rect 483244 272584 483258 272640
rect 483258 272584 483308 272640
rect 483244 272580 483308 272584
rect 486004 272640 486068 272644
rect 486004 272584 486018 272640
rect 486018 272584 486068 272640
rect 486004 272580 486068 272584
rect 118004 272444 118068 272508
rect 423812 272504 423876 272508
rect 423812 272448 423826 272504
rect 423826 272448 423876 272504
rect 423812 272444 423876 272448
rect 87644 272368 87708 272372
rect 87644 272312 87658 272368
rect 87658 272312 87708 272368
rect 87644 272308 87708 272312
rect 94452 272368 94516 272372
rect 94452 272312 94466 272368
rect 94466 272312 94516 272368
rect 94452 272308 94516 272312
rect 99420 272232 99484 272236
rect 99420 272176 99434 272232
rect 99434 272176 99484 272232
rect 99420 272172 99484 272176
rect 265204 272232 265268 272236
rect 265204 272176 265218 272232
rect 265218 272176 265268 272232
rect 265204 272172 265268 272176
rect 401732 272232 401796 272236
rect 401732 272176 401746 272232
rect 401746 272176 401796 272232
rect 401732 272172 401796 272176
rect 415900 272232 415964 272236
rect 415900 272176 415914 272232
rect 415914 272176 415964 272232
rect 415900 272172 415964 272176
rect 416084 272232 416148 272236
rect 416084 272176 416098 272232
rect 416098 272176 416148 272232
rect 416084 272172 416148 272176
rect 455828 272232 455892 272236
rect 455828 272176 455842 272232
rect 455842 272176 455892 272232
rect 455828 272172 455892 272176
rect 53236 271824 53300 271828
rect 53236 271768 53286 271824
rect 53286 271768 53300 271824
rect 53236 271764 53300 271768
rect 83964 271764 84028 271828
rect 97028 271764 97092 271828
rect 100708 271824 100772 271828
rect 100708 271768 100758 271824
rect 100758 271768 100772 271824
rect 100708 271764 100772 271768
rect 106412 271764 106476 271828
rect 107516 271764 107580 271828
rect 112300 271824 112364 271828
rect 112300 271768 112350 271824
rect 112350 271768 112364 271824
rect 112300 271764 112364 271768
rect 123524 271764 123588 271828
rect 125916 271764 125980 271828
rect 128676 271764 128740 271828
rect 150940 271764 151004 271828
rect 154068 271764 154132 271828
rect 155908 271764 155972 271828
rect 263548 271824 263612 271828
rect 263548 271768 263598 271824
rect 263598 271768 263612 271824
rect 263548 271764 263612 271768
rect 265940 271764 266004 271828
rect 268332 271764 268396 271828
rect 270908 271764 270972 271828
rect 272564 271764 272628 271828
rect 276244 271764 276308 271828
rect 278452 271764 278516 271828
rect 279004 271764 279068 271828
rect 280844 271764 280908 271828
rect 308628 271764 308692 271828
rect 313412 271764 313476 271828
rect 79548 271628 79612 271692
rect 84700 271688 84764 271692
rect 84700 271632 84714 271688
rect 84714 271632 84764 271688
rect 84700 271628 84764 271632
rect 98132 271688 98196 271692
rect 98132 271632 98146 271688
rect 98146 271632 98196 271688
rect 98132 271628 98196 271632
rect 108252 271628 108316 271692
rect 115980 271688 116044 271692
rect 115980 271632 115994 271688
rect 115994 271632 116044 271688
rect 115980 271628 116044 271632
rect 118372 271628 118436 271692
rect 120764 271628 120828 271692
rect 158484 271628 158548 271692
rect 160876 271628 160940 271692
rect 163452 271628 163516 271692
rect 166028 271628 166092 271692
rect 198780 271628 198844 271692
rect 315068 271628 315132 271692
rect 428596 271764 428660 271828
rect 433564 271764 433628 271828
rect 436876 271764 436940 271828
rect 438532 271764 438596 271828
rect 443500 271764 443564 271828
rect 445892 271764 445956 271828
rect 448284 271764 448348 271828
rect 451044 271764 451108 271828
rect 458404 271764 458468 271828
rect 465948 271628 466012 271692
rect 503116 271628 503180 271692
rect 101076 271492 101140 271556
rect 115796 271552 115860 271556
rect 115796 271496 115846 271552
rect 115846 271496 115860 271552
rect 115796 271492 115860 271496
rect 105860 271356 105924 271420
rect 109540 271356 109604 271420
rect 114324 271356 114388 271420
rect 183140 271356 183204 271420
rect 217180 271492 217244 271556
rect 273484 271492 273548 271556
rect 276980 271492 277044 271556
rect 343404 271492 343468 271556
rect 460980 271492 461044 271556
rect 236500 271356 236564 271420
rect 343220 271356 343284 271420
rect 377260 271356 377324 271420
rect 408172 271356 408236 271420
rect 440924 271356 440988 271420
rect 81940 271220 82004 271284
rect 88380 271280 88444 271284
rect 88380 271224 88394 271280
rect 88394 271224 88444 271280
rect 88380 271220 88444 271224
rect 103836 271220 103900 271284
rect 111012 271220 111076 271284
rect 113220 271280 113284 271284
rect 113220 271224 113234 271280
rect 113234 271224 113284 271280
rect 113220 271220 113284 271224
rect 237052 271220 237116 271284
rect 258396 271220 258460 271284
rect 260972 271220 261036 271284
rect 271276 271220 271340 271284
rect 396028 271220 396092 271284
rect 435956 271220 436020 271284
rect 503484 271280 503548 271284
rect 503484 271224 503534 271280
rect 503534 271224 503548 271280
rect 503484 271220 503548 271224
rect 119108 271084 119172 271148
rect 183508 271144 183572 271148
rect 183508 271088 183522 271144
rect 183522 271088 183572 271144
rect 183508 271084 183572 271088
rect 248276 271084 248340 271148
rect 253612 271084 253676 271148
rect 256188 271084 256252 271148
rect 397132 271084 397196 271148
rect 410748 271084 410812 271148
rect 413692 271084 413756 271148
rect 418476 271084 418540 271148
rect 78260 270948 78324 271012
rect 130884 270948 130948 271012
rect 325556 270948 325620 271012
rect 462636 270948 462700 271012
rect 80468 270812 80532 270876
rect 88748 270812 88812 270876
rect 254532 270812 254596 270876
rect 268700 270812 268764 270876
rect 278084 270812 278148 270876
rect 406516 270812 406580 270876
rect 432276 270812 432340 270876
rect 434668 270812 434732 270876
rect 438348 270812 438412 270876
rect 439084 270812 439148 270876
rect 90036 270676 90100 270740
rect 93348 270676 93412 270740
rect 105308 270676 105372 270740
rect 148548 270676 148612 270740
rect 244228 270676 244292 270740
rect 252324 270676 252388 270740
rect 255820 270676 255884 270740
rect 260604 270676 260668 270740
rect 411300 270736 411364 270740
rect 411300 270680 411350 270736
rect 411350 270680 411364 270736
rect 411300 270676 411364 270680
rect 429700 270676 429764 270740
rect 86540 270540 86604 270604
rect 91324 270540 91388 270604
rect 108620 270540 108684 270604
rect 111196 270540 111260 270604
rect 238156 270540 238220 270604
rect 242940 270600 243004 270604
rect 242940 270544 242954 270600
rect 242954 270544 243004 270600
rect 242940 270540 243004 270544
rect 245332 270540 245396 270604
rect 246436 270540 246500 270604
rect 247724 270540 247788 270604
rect 248644 270540 248708 270604
rect 250116 270540 250180 270604
rect 251220 270600 251284 270604
rect 251220 270544 251234 270600
rect 251234 270544 251284 270600
rect 251220 270540 251284 270544
rect 253428 270540 253492 270604
rect 256924 270540 256988 270604
rect 258396 270540 258460 270604
rect 259500 270600 259564 270604
rect 259500 270544 259514 270600
rect 259514 270544 259564 270600
rect 259500 270540 259564 270544
rect 262076 270540 262140 270604
rect 262812 270540 262876 270604
rect 263916 270540 263980 270604
rect 267596 270540 267660 270604
rect 269804 270540 269868 270604
rect 274404 270540 274468 270604
rect 275324 270540 275388 270604
rect 397500 270600 397564 270604
rect 397500 270544 397514 270600
rect 397514 270544 397564 270600
rect 397500 270540 397564 270544
rect 399524 270540 399588 270604
rect 400444 270540 400508 270604
rect 403020 270600 403084 270604
rect 403020 270544 403034 270600
rect 403034 270544 403084 270600
rect 403020 270540 403084 270544
rect 404124 270540 404188 270604
rect 405044 270540 405108 270604
rect 407620 270540 407684 270604
rect 408724 270540 408788 270604
rect 410012 270540 410076 270604
rect 412404 270540 412468 270604
rect 413324 270540 413388 270604
rect 414428 270540 414492 270604
rect 417004 270540 417068 270604
rect 418108 270600 418172 270604
rect 418108 270544 418158 270600
rect 418158 270544 418172 270600
rect 418108 270540 418172 270544
rect 420684 270540 420748 270604
rect 421788 270540 421852 270604
rect 57652 270268 57716 270332
rect 91508 270404 91572 270468
rect 323348 270404 323412 270468
rect 239260 270268 239324 270332
rect 435772 270404 435836 270468
rect 217548 269996 217612 270060
rect 241652 269860 241716 269924
rect 419212 269860 419276 269924
rect 240548 269724 240612 269788
rect 427676 269724 427740 269788
rect 44956 268500 45020 268564
rect 44772 268364 44836 268428
rect 376892 267548 376956 267612
rect 377444 267548 377508 267612
rect 54340 253948 54404 254012
rect 190868 253676 190932 253740
rect 338436 253540 338500 253604
rect 499804 253268 499868 253332
rect 178540 253132 178604 253196
rect 179644 253132 179708 253196
rect 350948 253132 351012 253196
rect 339724 252996 339788 253060
rect 498516 252724 498580 252788
rect 510844 252648 510908 252652
rect 510844 252592 510894 252648
rect 510894 252592 510908 252648
rect 510844 252588 510908 252592
rect 57652 252452 57716 252516
rect 216996 252452 217060 252516
rect 377996 252452 378060 252516
rect 57836 166908 57900 166972
rect 198044 166908 198108 166972
rect 370636 166908 370700 166972
rect 47900 166772 47964 166836
rect 93716 166772 93780 166836
rect 98500 166832 98564 166836
rect 98500 166776 98514 166832
rect 98514 166776 98564 166832
rect 98500 166772 98564 166776
rect 101076 166832 101140 166836
rect 101076 166776 101090 166832
rect 101090 166776 101140 166832
rect 101076 166772 101140 166776
rect 105860 166832 105924 166836
rect 105860 166776 105874 166832
rect 105874 166776 105924 166832
rect 105860 166772 105924 166776
rect 108252 166832 108316 166836
rect 108252 166776 108266 166832
rect 108266 166776 108316 166832
rect 108252 166772 108316 166776
rect 138478 166832 138542 166836
rect 138478 166776 138534 166832
rect 138534 166776 138542 166832
rect 138478 166772 138542 166776
rect 140926 166772 140990 166836
rect 143510 166772 143574 166836
rect 145958 166832 146022 166836
rect 145958 166776 145986 166832
rect 145986 166776 146022 166832
rect 145958 166772 146022 166776
rect 205036 166772 205100 166836
rect 305958 166772 306022 166836
rect 313438 166772 313502 166836
rect 418476 166832 418540 166836
rect 418476 166776 418490 166832
rect 418490 166776 418540 166832
rect 418476 166772 418540 166776
rect 421052 166832 421116 166836
rect 421052 166776 421066 166832
rect 421066 166776 421116 166832
rect 421052 166772 421116 166776
rect 423444 166832 423508 166836
rect 423444 166776 423458 166832
rect 423458 166776 423508 166832
rect 423444 166772 423508 166776
rect 428228 166832 428292 166836
rect 428228 166776 428242 166832
rect 428242 166776 428292 166832
rect 428228 166772 428292 166776
rect 445892 166832 445956 166836
rect 445892 166776 445906 166832
rect 445906 166776 445956 166832
rect 445892 166772 445956 166776
rect 470990 166832 471054 166836
rect 470990 166776 471022 166832
rect 471022 166776 471054 166832
rect 470990 166772 471054 166776
rect 473438 166772 473502 166836
rect 475886 166832 475950 166836
rect 475886 166776 475898 166832
rect 475898 166776 475950 166832
rect 475886 166772 475950 166776
rect 478470 166832 478534 166836
rect 478470 166776 478474 166832
rect 478474 166776 478534 166832
rect 478470 166772 478534 166776
rect 480918 166832 480982 166836
rect 480918 166776 480958 166832
rect 480958 166776 480982 166832
rect 480918 166772 480982 166776
rect 163366 166696 163430 166700
rect 163366 166640 163374 166696
rect 163374 166640 163430 166696
rect 163366 166636 163430 166640
rect 165950 166636 166014 166700
rect 213500 166636 213564 166700
rect 298478 166636 298542 166700
rect 303510 166696 303574 166700
rect 303510 166640 303526 166696
rect 303526 166640 303574 166696
rect 303510 166636 303574 166640
rect 483366 166696 483430 166700
rect 483366 166640 483386 166696
rect 483386 166640 483430 166696
rect 483366 166636 483430 166640
rect 485950 166696 486014 166700
rect 485950 166640 485962 166696
rect 485962 166640 486014 166696
rect 485950 166636 486014 166640
rect 114406 166560 114470 166564
rect 114406 166504 114430 166560
rect 114430 166504 114470 166560
rect 114406 166500 114470 166504
rect 116990 166560 117054 166564
rect 116990 166504 117006 166560
rect 117006 166504 117054 166560
rect 116990 166500 117054 166504
rect 148548 166560 148612 166564
rect 148548 166504 148562 166560
rect 148562 166504 148612 166560
rect 148548 166500 148612 166504
rect 153332 166560 153396 166564
rect 153332 166504 153346 166560
rect 153346 166504 153396 166560
rect 153332 166500 153396 166504
rect 183222 166560 183286 166564
rect 183222 166504 183282 166560
rect 183282 166504 183286 166560
rect 183222 166500 183286 166504
rect 207980 166500 208044 166564
rect 196572 166364 196636 166428
rect 260972 166424 261036 166428
rect 260972 166368 260986 166424
rect 260986 166368 261036 166424
rect 96108 166288 96172 166292
rect 96108 166232 96122 166288
rect 96122 166232 96172 166288
rect 96108 166228 96172 166232
rect 260972 166364 261036 166368
rect 265940 166424 266004 166428
rect 265940 166368 265954 166424
rect 265954 166368 266004 166424
rect 265940 166364 266004 166368
rect 285966 166560 286030 166564
rect 285966 166504 286010 166560
rect 286010 166504 286030 166560
rect 285966 166500 286030 166504
rect 288278 166560 288342 166564
rect 288278 166504 288310 166560
rect 288310 166504 288342 166560
rect 288278 166500 288342 166504
rect 290998 166500 291062 166564
rect 293446 166560 293510 166564
rect 293446 166504 293462 166560
rect 293462 166504 293510 166560
rect 293446 166500 293510 166504
rect 295894 166560 295958 166564
rect 295894 166504 295946 166560
rect 295946 166504 295958 166560
rect 295894 166500 295958 166504
rect 503222 166560 503286 166564
rect 503222 166504 503258 166560
rect 503258 166504 503286 166560
rect 503222 166500 503286 166504
rect 270908 166228 270972 166292
rect 81756 165548 81820 165612
rect 85436 165548 85500 165612
rect 90772 165548 90836 165612
rect 92428 165548 92492 165612
rect 95740 165548 95804 165612
rect 99420 165608 99484 165612
rect 99420 165552 99434 165608
rect 99434 165552 99484 165608
rect 99420 165548 99484 165552
rect 103468 165608 103532 165612
rect 103468 165552 103518 165608
rect 103518 165552 103532 165608
rect 103468 165548 103532 165552
rect 109724 165548 109788 165612
rect 111012 165548 111076 165612
rect 111196 165608 111260 165612
rect 111196 165552 111210 165608
rect 111210 165552 111260 165608
rect 111196 165548 111260 165552
rect 112300 165548 112364 165612
rect 113588 165608 113652 165612
rect 113588 165552 113602 165608
rect 113602 165552 113652 165608
rect 113588 165548 113652 165552
rect 115980 165608 116044 165612
rect 115980 165552 115994 165608
rect 115994 165552 116044 165608
rect 115980 165548 116044 165552
rect 118004 165608 118068 165612
rect 118004 165552 118018 165608
rect 118018 165552 118068 165608
rect 118004 165548 118068 165552
rect 118372 165608 118436 165612
rect 118372 165552 118386 165608
rect 118386 165552 118436 165608
rect 118372 165548 118436 165552
rect 119108 165548 119172 165612
rect 120948 165608 121012 165612
rect 120948 165552 120962 165608
rect 120962 165552 121012 165608
rect 120948 165548 121012 165552
rect 123524 165608 123588 165612
rect 123524 165552 123538 165608
rect 123538 165552 123588 165608
rect 123524 165548 123588 165552
rect 125916 165608 125980 165612
rect 125916 165552 125930 165608
rect 125930 165552 125980 165608
rect 125916 165548 125980 165552
rect 128492 165548 128556 165612
rect 130884 165548 130948 165612
rect 133460 165548 133524 165612
rect 183324 165608 183388 165612
rect 183324 165552 183374 165608
rect 183374 165552 183388 165608
rect 183324 165548 183388 165552
rect 235948 165608 236012 165612
rect 235948 165552 235998 165608
rect 235998 165552 236012 165608
rect 235948 165548 236012 165552
rect 239628 165548 239692 165612
rect 243124 165548 243188 165612
rect 247540 165548 247604 165612
rect 248276 165548 248340 165612
rect 250668 165548 250732 165612
rect 253612 165548 253676 165612
rect 258396 165548 258460 165612
rect 261708 165548 261772 165612
rect 265204 165548 265268 165612
rect 268332 165548 268396 165612
rect 272196 165548 272260 165612
rect 273484 165608 273548 165612
rect 273484 165552 273498 165608
rect 273498 165552 273548 165608
rect 273484 165548 273548 165552
rect 275876 165608 275940 165612
rect 275876 165552 275926 165608
rect 275926 165552 275940 165608
rect 275876 165548 275940 165552
rect 276060 165548 276124 165612
rect 278452 165548 278516 165612
rect 279188 165548 279252 165612
rect 280844 165548 280908 165612
rect 283420 165608 283484 165612
rect 283420 165552 283434 165608
rect 283434 165552 283484 165608
rect 283420 165548 283484 165552
rect 300900 165608 300964 165612
rect 300900 165552 300914 165608
rect 300914 165552 300964 165608
rect 300900 165548 300964 165552
rect 323348 165608 323412 165612
rect 323348 165552 323362 165608
rect 323362 165552 323412 165608
rect 323348 165548 323412 165552
rect 343404 165608 343468 165612
rect 343404 165552 343454 165608
rect 343454 165552 343468 165608
rect 343404 165548 343468 165552
rect 398236 165548 398300 165612
rect 401732 165548 401796 165612
rect 405412 165548 405476 165612
rect 410748 165548 410812 165612
rect 415900 165548 415964 165612
rect 416084 165608 416148 165612
rect 416084 165552 416098 165608
rect 416098 165552 416148 165608
rect 416084 165548 416148 165552
rect 419396 165548 419460 165612
rect 423812 165608 423876 165612
rect 423812 165552 423826 165608
rect 423826 165552 423876 165608
rect 423812 165548 423876 165552
rect 434300 165548 434364 165612
rect 435956 165548 436020 165612
rect 436876 165548 436940 165612
rect 437796 165608 437860 165612
rect 437796 165552 437810 165608
rect 437810 165552 437860 165608
rect 437796 165548 437860 165552
rect 438532 165548 438596 165612
rect 439268 165548 439332 165612
rect 443500 165548 443564 165612
rect 448284 165548 448348 165612
rect 451044 165548 451108 165612
rect 453436 165548 453500 165612
rect 455828 165548 455892 165612
rect 458404 165608 458468 165612
rect 458404 165552 458418 165608
rect 458418 165552 458468 165608
rect 458404 165548 458468 165552
rect 503300 165608 503364 165612
rect 503300 165552 503350 165608
rect 503350 165552 503364 165608
rect 503300 165548 503364 165552
rect 158484 165412 158548 165476
rect 208900 165412 208964 165476
rect 325924 165412 325988 165476
rect 343220 165412 343284 165476
rect 468524 165412 468588 165476
rect 155908 165276 155972 165340
rect 204852 165276 204916 165340
rect 315804 165276 315868 165340
rect 150940 165140 151004 165204
rect 213316 165140 213380 165204
rect 311020 165140 311084 165204
rect 379652 165140 379716 165204
rect 463556 165276 463620 165340
rect 460980 165140 461044 165204
rect 136036 165004 136100 165068
rect 216260 165004 216324 165068
rect 308628 165004 308692 165068
rect 426020 165004 426084 165068
rect 440924 165004 440988 165068
rect 88380 164928 88444 164932
rect 88380 164872 88394 164928
rect 88394 164872 88444 164928
rect 88380 164868 88444 164872
rect 108620 164868 108684 164932
rect 206508 164868 206572 164932
rect 263732 164868 263796 164932
rect 408172 164868 408236 164932
rect 433564 164868 433628 164932
rect 107516 164732 107580 164796
rect 200988 164732 201052 164796
rect 256188 164732 256252 164796
rect 413692 164732 413756 164796
rect 421788 164732 421852 164796
rect 431172 164732 431236 164796
rect 50476 164596 50540 164660
rect 160876 164596 160940 164660
rect 267596 164596 267660 164660
rect 465948 164596 466012 164660
rect 100708 164520 100772 164524
rect 100708 164464 100758 164520
rect 100758 164464 100772 164520
rect 100708 164460 100772 164464
rect 113220 164460 113284 164524
rect 115796 164460 115860 164524
rect 244412 164520 244476 164524
rect 244412 164464 244426 164520
rect 244426 164464 244476 164520
rect 244412 164460 244476 164464
rect 252324 164460 252388 164524
rect 260604 164460 260668 164524
rect 266492 164460 266556 164524
rect 273300 164460 273364 164524
rect 77156 164324 77220 164388
rect 90036 164324 90100 164388
rect 202460 164324 202524 164388
rect 320956 164324 321020 164388
rect 397132 164324 397196 164388
rect 404124 164324 404188 164388
rect 412404 164324 412468 164388
rect 426388 164324 426452 164388
rect 429700 164324 429764 164388
rect 76052 164188 76116 164252
rect 78260 164188 78324 164252
rect 79548 164188 79612 164252
rect 80468 164188 80532 164252
rect 83044 164188 83108 164252
rect 84148 164188 84212 164252
rect 86540 164188 86604 164252
rect 87644 164188 87708 164252
rect 88748 164188 88812 164252
rect 91324 164188 91388 164252
rect 93348 164188 93412 164252
rect 94452 164188 94516 164252
rect 97028 164188 97092 164252
rect 98132 164188 98196 164252
rect 101812 164188 101876 164252
rect 102732 164188 102796 164252
rect 103836 164188 103900 164252
rect 105308 164188 105372 164252
rect 106412 164248 106476 164252
rect 106412 164192 106426 164248
rect 106426 164192 106476 164248
rect 106412 164188 106476 164192
rect 237052 164188 237116 164252
rect 238156 164188 238220 164252
rect 240548 164188 240612 164252
rect 241652 164188 241716 164252
rect 245332 164188 245396 164252
rect 246436 164188 246500 164252
rect 248644 164188 248708 164252
rect 250116 164188 250180 164252
rect 251220 164248 251284 164252
rect 251220 164192 251234 164248
rect 251234 164192 251284 164248
rect 251220 164188 251284 164192
rect 253428 164188 253492 164252
rect 254532 164188 254596 164252
rect 255820 164188 255884 164252
rect 256924 164188 256988 164252
rect 258396 164188 258460 164252
rect 259500 164248 259564 164252
rect 259500 164192 259514 164248
rect 259514 164192 259564 164248
rect 259500 164188 259564 164192
rect 262812 164188 262876 164252
rect 263916 164188 263980 164252
rect 268700 164188 268764 164252
rect 269804 164188 269868 164252
rect 271276 164188 271340 164252
rect 274404 164188 274468 164252
rect 276980 164188 277044 164252
rect 278084 164188 278148 164252
rect 57652 164052 57716 164116
rect 206324 164052 206388 164116
rect 318380 164188 318444 164252
rect 396028 164248 396092 164252
rect 396028 164192 396078 164248
rect 396078 164192 396092 164248
rect 396028 164188 396092 164192
rect 399524 164188 399588 164252
rect 400444 164188 400508 164252
rect 403020 164248 403084 164252
rect 403020 164192 403070 164248
rect 403070 164192 403084 164248
rect 403020 164188 403084 164192
rect 406516 164188 406580 164252
rect 407620 164188 407684 164252
rect 408724 164188 408788 164252
rect 410012 164188 410076 164252
rect 411300 164248 411364 164252
rect 411300 164192 411350 164248
rect 411350 164192 411364 164248
rect 411300 164188 411364 164192
rect 413324 164188 413388 164252
rect 414428 164188 414492 164252
rect 417004 164188 417068 164252
rect 418292 164188 418356 164252
rect 420684 164188 420748 164252
rect 422892 164188 422956 164252
rect 425284 164188 425348 164252
rect 427676 164248 427740 164252
rect 427676 164192 427726 164248
rect 427726 164192 427740 164248
rect 427676 164188 427740 164192
rect 428780 164188 428844 164252
rect 430988 164188 431052 164252
rect 432276 164188 432340 164252
rect 433380 164188 433444 164252
rect 435772 164188 435836 164252
rect 376892 164052 376956 164116
rect 217180 162692 217244 162756
rect 376892 162692 376956 162756
rect 363460 149092 363524 149156
rect 57652 147732 57716 147796
rect 377444 147732 377508 147796
rect 217548 146236 217612 146300
rect 377996 146236 378060 146300
rect 377628 145828 377692 145892
rect 377812 145556 377876 145620
rect 510844 145420 510908 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 190868 144876 190932 144940
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144876 499868 144940
rect 57468 140796 57532 140860
rect 375420 68852 375484 68916
rect 46796 67764 46860 67828
rect 214604 68036 214668 68100
rect 218652 60616 218716 60620
rect 218652 60560 218702 60616
rect 218702 60560 218716 60616
rect 218652 60556 218716 60560
rect 219204 60616 219268 60620
rect 219204 60560 219254 60616
rect 219254 60560 219268 60616
rect 219204 60556 219268 60560
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 94550 59800 94614 59804
rect 94550 59744 94558 59800
rect 94558 59744 94614 59800
rect 94550 59740 94614 59744
rect 101758 59800 101822 59804
rect 101758 59744 101770 59800
rect 101770 59744 101822 59800
rect 101758 59740 101822 59744
rect 102846 59740 102910 59804
rect 113590 59800 113654 59804
rect 113590 59744 113602 59800
rect 113602 59744 113654 59800
rect 113590 59740 113654 59744
rect 237142 59800 237206 59804
rect 237142 59744 237158 59800
rect 237158 59744 237206 59800
rect 237142 59740 237206 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 256998 59800 257062 59804
rect 256998 59744 257030 59800
rect 257030 59744 257062 59800
rect 256998 59740 257062 59744
rect 262846 59800 262910 59804
rect 262846 59744 262862 59800
rect 262862 59744 262910 59800
rect 262846 59740 262910 59744
rect 263934 59740 263998 59804
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 416998 59800 417062 59804
rect 416998 59744 417018 59800
rect 417018 59744 417062 59800
rect 416998 59740 417062 59744
rect 423526 59800 423590 59804
rect 423526 59744 423550 59800
rect 423550 59744 423590 59800
rect 423526 59740 423590 59744
rect 423934 59800 423998 59804
rect 423934 59744 423954 59800
rect 423954 59744 423998 59800
rect 423934 59740 423998 59744
rect 57652 59468 57716 59532
rect 105294 59604 105358 59668
rect 105974 59604 106038 59668
rect 107606 59664 107670 59668
rect 107606 59608 107622 59664
rect 107622 59608 107670 59664
rect 107606 59604 107670 59608
rect 258086 59664 258150 59668
rect 258086 59608 258134 59664
rect 258134 59608 258150 59664
rect 258086 59604 258150 59608
rect 260670 59664 260734 59668
rect 260670 59608 260710 59664
rect 260710 59608 260734 59664
rect 260670 59604 260734 59608
rect 261758 59664 261822 59668
rect 261758 59608 261814 59664
rect 261814 59608 261822 59664
rect 261758 59604 261822 59608
rect 308542 59664 308606 59668
rect 308542 59608 308550 59664
rect 308550 59608 308606 59664
rect 308542 59604 308606 59608
rect 315886 59664 315950 59668
rect 315886 59608 315910 59664
rect 315910 59608 315950 59664
rect 315886 59604 315950 59608
rect 403126 59604 403190 59668
rect 404214 59664 404278 59668
rect 404214 59608 404230 59664
rect 404230 59608 404278 59664
rect 404214 59604 404278 59608
rect 90036 59528 90100 59532
rect 90036 59472 90050 59528
rect 90050 59472 90100 59528
rect 90036 59468 90100 59472
rect 95924 59528 95988 59532
rect 95924 59472 95938 59528
rect 95938 59472 95988 59528
rect 95924 59468 95988 59472
rect 97028 59528 97092 59532
rect 97028 59472 97042 59528
rect 97042 59472 97092 59528
rect 97028 59468 97092 59472
rect 98132 59528 98196 59532
rect 98132 59472 98146 59528
rect 98146 59472 98196 59528
rect 98132 59468 98196 59472
rect 100708 59528 100772 59532
rect 413462 59604 413526 59668
rect 416046 59664 416110 59668
rect 416046 59608 416098 59664
rect 416098 59608 416110 59664
rect 416046 59604 416110 59608
rect 419446 59664 419510 59668
rect 419446 59608 419502 59664
rect 419502 59608 419510 59664
rect 419446 59604 419510 59608
rect 421758 59664 421822 59668
rect 421758 59608 421802 59664
rect 421802 59608 421822 59664
rect 421758 59604 421822 59608
rect 458478 59664 458542 59668
rect 458478 59608 458510 59664
rect 458510 59608 458542 59664
rect 458478 59604 458542 59608
rect 503222 59664 503286 59668
rect 503222 59608 503258 59664
rect 503258 59608 503286 59664
rect 503222 59604 503286 59608
rect 100708 59472 100758 59528
rect 100758 59472 100772 59528
rect 100708 59468 100772 59472
rect 410748 59528 410812 59532
rect 410748 59472 410762 59528
rect 410762 59472 410812 59528
rect 46612 59332 46676 59396
rect 410748 59468 410812 59472
rect 418108 59528 418172 59532
rect 418108 59472 418158 59528
rect 418158 59472 418172 59528
rect 418108 59468 418172 59472
rect 420684 59528 420748 59532
rect 420684 59472 420698 59528
rect 420698 59472 420748 59528
rect 420684 59468 420748 59472
rect 111012 59392 111076 59396
rect 111012 59336 111026 59392
rect 111026 59336 111076 59392
rect 111012 59332 111076 59336
rect 200804 59332 200868 59396
rect 263548 59332 263612 59396
rect 279188 59392 279252 59396
rect 279188 59336 279238 59392
rect 279238 59336 279252 59392
rect 279188 59332 279252 59336
rect 377628 59332 377692 59396
rect 422892 59332 422956 59396
rect 426020 59392 426084 59396
rect 426020 59336 426034 59392
rect 426034 59336 426084 59392
rect 426020 59332 426084 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 453436 59392 453500 59396
rect 453436 59336 453450 59392
rect 453450 59336 453500 59392
rect 453436 59332 453500 59336
rect 54708 59196 54772 59260
rect 143580 59196 143644 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 198412 59196 198476 59260
rect 280844 59196 280908 59260
rect 290964 59256 291028 59260
rect 290964 59200 290978 59256
rect 290978 59200 291028 59256
rect 290964 59196 291028 59200
rect 300900 59256 300964 59260
rect 300900 59200 300914 59256
rect 300914 59200 300964 59256
rect 300900 59196 300964 59200
rect 320956 59256 321020 59260
rect 320956 59200 320970 59256
rect 320970 59200 321020 59256
rect 320956 59196 321020 59200
rect 325924 59256 325988 59260
rect 325924 59200 325938 59256
rect 325938 59200 325988 59256
rect 325924 59196 325988 59200
rect 357940 59196 358004 59260
rect 480852 59196 480916 59260
rect 55628 59060 55692 59124
rect 140820 59060 140884 59124
rect 212396 59060 212460 59124
rect 285996 59060 286060 59124
rect 371740 59060 371804 59124
rect 483428 59060 483492 59124
rect 53420 58924 53484 58988
rect 138428 58924 138492 58988
rect 201356 58924 201420 58988
rect 273484 58924 273548 58988
rect 367876 58924 367940 58988
rect 468524 58924 468588 58988
rect 475884 58984 475948 58988
rect 475884 58928 475898 58984
rect 475898 58928 475948 58984
rect 475884 58924 475948 58928
rect 52132 58788 52196 58852
rect 135852 58788 135916 58852
rect 209636 58788 209700 58852
rect 276060 58788 276124 58852
rect 375972 58788 376036 58852
rect 473492 58788 473556 58852
rect 59308 58652 59372 58716
rect 120948 58652 121012 58716
rect 197860 58652 197924 58716
rect 253612 58652 253676 58716
rect 374684 58652 374748 58716
rect 463556 58652 463620 58716
rect 48084 58516 48148 58580
rect 108252 58516 108316 58580
rect 200620 58516 200684 58580
rect 250668 58516 250732 58580
rect 59124 58380 59188 58444
rect 101076 58380 101140 58444
rect 217364 58380 217428 58444
rect 259500 58380 259564 58444
rect 85436 58108 85500 58172
rect 92428 58108 92492 58172
rect 99420 58108 99484 58172
rect 113220 58108 113284 58172
rect 153332 58108 153396 58172
rect 235948 58108 236012 58172
rect 265204 58108 265268 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 398236 58108 398300 58172
rect 401732 58108 401796 58172
rect 405412 58108 405476 58172
rect 455828 58108 455892 58172
rect 83964 57972 84028 58036
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57836 79612 57900
rect 80468 57896 80532 57900
rect 80468 57840 80482 57896
rect 80482 57840 80532 57896
rect 80468 57836 80532 57840
rect 81940 57836 82004 57900
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88380 57896 88444 57900
rect 88380 57840 88394 57896
rect 88394 57840 88444 57896
rect 88380 57836 88444 57840
rect 88748 57896 88812 57900
rect 88748 57840 88762 57896
rect 88762 57840 88812 57896
rect 88748 57836 88812 57840
rect 90772 57896 90836 57900
rect 90772 57840 90786 57896
rect 90786 57840 90836 57896
rect 90772 57836 90836 57840
rect 91324 57836 91388 57900
rect 93348 57896 93412 57900
rect 93348 57840 93362 57896
rect 93362 57840 93412 57896
rect 93348 57836 93412 57840
rect 93716 57896 93780 57900
rect 93716 57840 93730 57896
rect 93730 57840 93780 57896
rect 93716 57836 93780 57840
rect 103836 57896 103900 57900
rect 103836 57840 103850 57896
rect 103850 57840 103900 57896
rect 103836 57836 103900 57840
rect 106412 57836 106476 57900
rect 108620 57836 108684 57900
rect 109540 57836 109604 57900
rect 111196 57896 111260 57900
rect 111196 57840 111210 57896
rect 111210 57840 111260 57896
rect 111196 57836 111260 57840
rect 112116 57896 112180 57900
rect 112116 57840 112130 57896
rect 112130 57840 112180 57896
rect 112116 57836 112180 57840
rect 115796 57896 115860 57900
rect 115796 57840 115810 57896
rect 115810 57840 115860 57896
rect 115796 57836 115860 57840
rect 115980 57896 116044 57900
rect 115980 57840 115994 57896
rect 115994 57840 116044 57896
rect 115980 57836 116044 57840
rect 119108 57896 119172 57900
rect 119108 57840 119122 57896
rect 119122 57840 119172 57896
rect 119108 57836 119172 57840
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 133460 57896 133524 57900
rect 133460 57840 133474 57896
rect 133474 57840 133524 57896
rect 133460 57836 133524 57840
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 183508 57896 183572 57900
rect 183508 57840 183522 57896
rect 183522 57840 183572 57896
rect 183508 57836 183572 57840
rect 238156 57836 238220 57900
rect 239260 57896 239324 57900
rect 239260 57840 239274 57896
rect 239274 57840 239324 57896
rect 239260 57836 239324 57840
rect 240548 57836 240612 57900
rect 241652 57896 241716 57900
rect 241652 57840 241666 57896
rect 241666 57840 241716 57896
rect 241652 57836 241716 57840
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 244228 57836 244292 57900
rect 245332 57896 245396 57900
rect 245332 57840 245346 57896
rect 245346 57840 245396 57896
rect 245332 57836 245396 57840
rect 246436 57836 246500 57900
rect 247724 57836 247788 57900
rect 248276 57896 248340 57900
rect 248276 57840 248290 57896
rect 248290 57840 248340 57896
rect 248276 57836 248340 57840
rect 248644 57896 248708 57900
rect 248644 57840 248658 57896
rect 248658 57840 248708 57896
rect 248644 57836 248708 57840
rect 250116 57836 250180 57900
rect 251220 57896 251284 57900
rect 251220 57840 251234 57896
rect 251234 57840 251284 57896
rect 251220 57836 251284 57840
rect 252324 57836 252388 57900
rect 253428 57896 253492 57900
rect 253428 57840 253442 57896
rect 253442 57840 253492 57896
rect 253428 57836 253492 57840
rect 254532 57836 254596 57900
rect 258396 57896 258460 57900
rect 258396 57840 258410 57896
rect 258410 57840 258460 57896
rect 258396 57836 258460 57840
rect 267596 57836 267660 57900
rect 268700 57836 268764 57900
rect 270908 57836 270972 57900
rect 271092 57896 271156 57900
rect 271092 57840 271106 57896
rect 271106 57840 271156 57896
rect 271092 57836 271156 57840
rect 273300 57896 273364 57900
rect 273300 57840 273314 57896
rect 273314 57840 273364 57896
rect 273300 57836 273364 57840
rect 276980 57896 277044 57900
rect 276980 57840 276994 57896
rect 276994 57840 277044 57896
rect 276980 57836 277044 57840
rect 278452 57836 278516 57900
rect 295932 57896 295996 57900
rect 295932 57840 295946 57896
rect 295946 57840 295996 57896
rect 295932 57836 295996 57840
rect 298508 57836 298572 57900
rect 303476 57896 303540 57900
rect 303476 57840 303490 57896
rect 303490 57840 303540 57896
rect 303476 57836 303540 57840
rect 305868 57896 305932 57900
rect 305868 57840 305882 57896
rect 305882 57840 305932 57896
rect 305868 57836 305932 57840
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 313412 57896 313476 57900
rect 313412 57840 313426 57896
rect 313426 57840 313476 57896
rect 313412 57836 313476 57840
rect 318380 57836 318444 57900
rect 323348 57896 323412 57900
rect 323348 57840 323362 57896
rect 323362 57840 323412 57896
rect 323348 57836 323412 57840
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57896 399588 57900
rect 399524 57840 399538 57896
rect 399538 57840 399588 57896
rect 399524 57836 399588 57840
rect 400444 57836 400508 57900
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 414612 57896 414676 57900
rect 414612 57840 414626 57896
rect 414626 57840 414676 57896
rect 414612 57836 414676 57840
rect 415532 57896 415596 57900
rect 415532 57840 415546 57896
rect 415546 57840 415596 57896
rect 415532 57836 415596 57840
rect 426388 57836 426452 57900
rect 427676 57896 427740 57900
rect 427676 57840 427690 57896
rect 427690 57840 427740 57896
rect 427676 57836 427740 57840
rect 428596 57836 428660 57900
rect 429700 57836 429764 57900
rect 431172 57836 431236 57900
rect 432276 57896 432340 57900
rect 432276 57840 432290 57896
rect 432290 57840 432340 57896
rect 432276 57836 432340 57840
rect 434668 57836 434732 57900
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 436876 57836 436940 57900
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 445892 57896 445956 57900
rect 445892 57840 445906 57896
rect 445906 57840 445956 57896
rect 445892 57836 445956 57840
rect 451044 57896 451108 57900
rect 451044 57840 451058 57896
rect 451058 57840 451108 57896
rect 451044 57836 451108 57840
rect 460980 57896 461044 57900
rect 460980 57840 460994 57896
rect 460994 57840 461044 57896
rect 60228 57700 60292 57764
rect 125916 57700 125980 57764
rect 183140 57760 183204 57764
rect 183140 57704 183190 57760
rect 183190 57704 183204 57760
rect 183140 57700 183204 57704
rect 214420 57700 214484 57764
rect 288204 57700 288268 57764
rect 374500 57700 374564 57764
rect 460980 57836 461044 57840
rect 465948 57896 466012 57900
rect 465948 57840 465962 57896
rect 465962 57840 466012 57896
rect 465948 57836 466012 57840
rect 470916 57896 470980 57900
rect 470916 57840 470930 57896
rect 470930 57840 470980 57896
rect 470916 57836 470980 57840
rect 478460 57896 478524 57900
rect 478460 57840 478474 57896
rect 478474 57840 478524 57896
rect 478460 57836 478524 57840
rect 486004 57896 486068 57900
rect 486004 57840 486018 57896
rect 486018 57840 486068 57896
rect 486004 57836 486068 57840
rect 503300 57896 503364 57900
rect 503300 57840 503350 57896
rect 503350 57840 503364 57896
rect 503300 57836 503364 57840
rect 54892 57564 54956 57628
rect 116900 57564 116964 57628
rect 123524 57564 123588 57628
rect 160876 57564 160940 57628
rect 163268 57564 163332 57628
rect 165844 57564 165908 57628
rect 202276 57564 202340 57628
rect 269804 57564 269868 57628
rect 274404 57564 274468 57628
rect 278084 57564 278148 57628
rect 370452 57564 370516 57628
rect 433380 57624 433444 57628
rect 433380 57568 433430 57624
rect 433430 57568 433444 57624
rect 433380 57564 433444 57568
rect 435772 57564 435836 57628
rect 438348 57564 438412 57628
rect 57836 57428 57900 57492
rect 118004 57428 118068 57492
rect 216076 57428 216140 57492
rect 283788 57428 283852 57492
rect 379100 57428 379164 57492
rect 448284 57428 448348 57492
rect 58572 57292 58636 57356
rect 58940 57156 59004 57220
rect 98500 57156 98564 57220
rect 113036 57292 113100 57356
rect 118372 57292 118436 57356
rect 203196 57292 203260 57356
rect 256004 57292 256068 57356
rect 266308 57352 266372 57356
rect 266308 57296 266358 57352
rect 266358 57296 266372 57352
rect 266308 57292 266372 57296
rect 371924 57292 371988 57356
rect 433564 57292 433628 57356
rect 103836 57156 103900 57220
rect 113220 57156 113284 57220
rect 114324 57156 114388 57220
rect 213132 57156 213196 57220
rect 265940 57156 266004 57220
rect 378916 57156 378980 57220
rect 418476 57156 418540 57220
rect 430988 57216 431052 57220
rect 430988 57160 431002 57216
rect 431002 57160 431052 57216
rect 430988 57156 431052 57160
rect 440924 57156 440988 57220
rect 58756 57020 58820 57084
rect 96292 57020 96356 57084
rect 215892 57020 215956 57084
rect 260972 57020 261036 57084
rect 378732 57020 378796 57084
rect 413508 57020 413572 57084
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 55076 56612 55140 56676
rect 128676 56612 128740 56676
rect 155908 56612 155972 56676
rect 158484 56612 158548 56676
rect 210556 56612 210620 56676
rect 293356 56612 293420 56676
rect 358124 56612 358188 56676
rect 443500 56748 443564 56812
rect 439084 56612 439148 56676
rect 50844 56476 50908 56540
rect 53604 56340 53668 56404
rect 219940 56476 220004 56540
rect 421052 56476 421116 56540
rect 198596 56340 198660 56404
rect 268332 56340 268396 56404
rect 377444 56340 377508 56404
rect 51764 56204 51828 56268
rect 377812 56204 377876 56268
rect 425284 56204 425348 56268
rect 57468 56068 57532 56132
rect 48636 55116 48700 55180
rect 50660 54980 50724 55044
rect 55444 54844 55508 54908
rect 210372 3980 210436 4044
rect 202092 3844 202156 3908
rect 360700 3708 360764 3772
rect 364932 3572 364996 3636
rect 365116 3436 365180 3500
rect 367692 3300 367756 3364
rect 206140 3164 206204 3228
rect 366956 3164 367020 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 54339 639436 54405 639437
rect 54339 639372 54340 639436
rect 54404 639372 54405 639436
rect 54339 639371 54405 639372
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 46795 482764 46861 482765
rect 46795 482700 46796 482764
rect 46860 482700 46861 482764
rect 46795 482699 46861 482700
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 44771 477188 44837 477189
rect 44771 477124 44772 477188
rect 44836 477124 44837 477188
rect 44771 477123 44837 477124
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 44774 268429 44834 477123
rect 44955 477052 45021 477053
rect 44955 476988 44956 477052
rect 45020 476988 45021 477052
rect 44955 476987 45021 476988
rect 44958 268565 45018 476987
rect 45234 442894 45854 478338
rect 46611 468892 46677 468893
rect 46611 468828 46612 468892
rect 46676 468828 46677 468892
rect 46611 468827 46677 468828
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 44955 268564 45021 268565
rect 44955 268500 44956 268564
rect 45020 268500 45021 268564
rect 44955 268499 45021 268500
rect 44771 268428 44837 268429
rect 44771 268364 44772 268428
rect 44836 268364 44837 268428
rect 44771 268363 44837 268364
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 46614 59397 46674 468827
rect 46798 67829 46858 482699
rect 48954 482614 49574 518058
rect 51947 485348 52013 485349
rect 51947 485284 51948 485348
rect 52012 485284 52013 485348
rect 51947 485283 52013 485284
rect 50291 484532 50357 484533
rect 50291 484468 50292 484532
rect 50356 484468 50357 484532
rect 50291 484467 50357 484468
rect 50843 484532 50909 484533
rect 50843 484468 50844 484532
rect 50908 484468 50909 484532
rect 50843 484467 50909 484468
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 47899 469844 47965 469845
rect 47899 469780 47900 469844
rect 47964 469780 47965 469844
rect 47899 469779 47965 469780
rect 47902 166837 47962 469779
rect 48083 469028 48149 469029
rect 48083 468964 48084 469028
rect 48148 468964 48149 469028
rect 48083 468963 48149 468964
rect 47899 166836 47965 166837
rect 47899 166772 47900 166836
rect 47964 166772 47965 166836
rect 47899 166771 47965 166772
rect 46795 67828 46861 67829
rect 46795 67764 46796 67828
rect 46860 67764 46861 67828
rect 46795 67763 46861 67764
rect 46611 59396 46677 59397
rect 46611 59332 46612 59396
rect 46676 59332 46677 59396
rect 46611 59331 46677 59332
rect 48086 58581 48146 468963
rect 48635 467940 48701 467941
rect 48635 467876 48636 467940
rect 48700 467876 48701 467940
rect 48635 467875 48701 467876
rect 48083 58580 48149 58581
rect 48083 58516 48084 58580
rect 48148 58516 48149 58580
rect 48083 58515 48149 58516
rect 48638 55181 48698 467875
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 50294 379541 50354 484467
rect 50475 468484 50541 468485
rect 50475 468420 50476 468484
rect 50540 468420 50541 468484
rect 50475 468419 50541 468420
rect 50291 379540 50357 379541
rect 50291 379476 50292 379540
rect 50356 379476 50357 379540
rect 50291 379475 50357 379476
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 50478 164661 50538 468419
rect 50659 467940 50725 467941
rect 50659 467876 50660 467940
rect 50724 467876 50725 467940
rect 50659 467875 50725 467876
rect 50475 164660 50541 164661
rect 50475 164596 50476 164660
rect 50540 164596 50541 164660
rect 50475 164595 50541 164596
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48635 55180 48701 55181
rect 48635 55116 48636 55180
rect 48700 55116 48701 55180
rect 48635 55115 48701 55116
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50662 55045 50722 467875
rect 50846 56541 50906 484467
rect 51579 465900 51645 465901
rect 51579 465836 51580 465900
rect 51644 465836 51645 465900
rect 51579 465835 51645 465836
rect 51582 282301 51642 465835
rect 51763 465220 51829 465221
rect 51763 465156 51764 465220
rect 51828 465156 51829 465220
rect 51763 465155 51829 465156
rect 51579 282300 51645 282301
rect 51579 282236 51580 282300
rect 51644 282236 51645 282300
rect 51579 282235 51645 282236
rect 50843 56540 50909 56541
rect 50843 56476 50844 56540
rect 50908 56476 50909 56540
rect 50843 56475 50909 56476
rect 51766 56269 51826 465155
rect 51950 379541 52010 485283
rect 53235 485212 53301 485213
rect 53235 485148 53236 485212
rect 53300 485148 53301 485212
rect 53235 485147 53301 485148
rect 53051 465900 53117 465901
rect 53051 465836 53052 465900
rect 53116 465836 53117 465900
rect 53051 465835 53117 465836
rect 52131 465764 52197 465765
rect 52131 465700 52132 465764
rect 52196 465700 52197 465764
rect 52131 465699 52197 465700
rect 51947 379540 52013 379541
rect 51947 379476 51948 379540
rect 52012 379476 52013 379540
rect 51947 379475 52013 379476
rect 52134 58853 52194 465699
rect 53054 388517 53114 465835
rect 53051 388516 53117 388517
rect 53051 388452 53052 388516
rect 53116 388452 53117 388516
rect 53051 388451 53117 388452
rect 53238 271829 53298 485147
rect 53603 468620 53669 468621
rect 53603 468556 53604 468620
rect 53668 468556 53669 468620
rect 53603 468555 53669 468556
rect 53419 466172 53485 466173
rect 53419 466108 53420 466172
rect 53484 466108 53485 466172
rect 53419 466107 53485 466108
rect 53235 271828 53301 271829
rect 53235 271764 53236 271828
rect 53300 271764 53301 271828
rect 53235 271763 53301 271764
rect 53422 58989 53482 466107
rect 53419 58988 53485 58989
rect 53419 58924 53420 58988
rect 53484 58924 53485 58988
rect 53419 58923 53485 58924
rect 52131 58852 52197 58853
rect 52131 58788 52132 58852
rect 52196 58788 52197 58852
rect 52131 58787 52197 58788
rect 53606 56405 53666 468555
rect 54342 254013 54402 639371
rect 55794 633454 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 640099 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 640099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 640099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 640099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 640099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 640099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 640099 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 640099 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 640099 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 640099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 640099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 640099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 640099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 640099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 640099 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 79568 633454 79888 633486
rect 79568 633218 79610 633454
rect 79846 633218 79888 633454
rect 79568 633134 79888 633218
rect 79568 632898 79610 633134
rect 79846 632898 79888 633134
rect 79568 632866 79888 632898
rect 110288 633454 110608 633486
rect 110288 633218 110330 633454
rect 110566 633218 110608 633454
rect 110288 633134 110608 633218
rect 110288 632898 110330 633134
rect 110566 632898 110608 633134
rect 110288 632866 110608 632898
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 565174 60134 573000
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 550000 60134 564618
rect 63234 568894 63854 573000
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 550000 63854 568338
rect 66954 572614 67574 573000
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 550000 67574 572058
rect 73794 562394 74414 573000
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 74414 562394
rect 73794 562074 74414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 74414 562074
rect 73794 550000 74414 561838
rect 77514 564234 78134 573000
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 78134 564234
rect 77514 563914 78134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 78134 563914
rect 77514 550000 78134 563678
rect 81234 550894 81854 573000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 550000 81854 550338
rect 84954 554614 85574 573000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 550000 85574 554058
rect 91794 561454 92414 573000
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 550000 92414 560898
rect 95514 565174 96134 573000
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 550000 96134 564618
rect 99234 568894 99854 573000
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 550000 99854 568338
rect 102954 572614 103574 573000
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 550000 103574 572058
rect 109794 562394 110414 573000
rect 109794 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 110414 562394
rect 109794 562074 110414 562158
rect 109794 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 110414 562074
rect 109794 550000 110414 561838
rect 113514 564234 114134 573000
rect 113514 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 114134 564234
rect 113514 563914 114134 563998
rect 113514 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 114134 563914
rect 113514 550000 114134 563678
rect 117234 550894 117854 573000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 550000 117854 550338
rect 120954 554614 121574 573000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 550000 121574 554058
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 550000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 550000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 550000 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 550000 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 640099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 640099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 640099 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 640099 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 640099 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 640099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 640099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 640099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 640099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 640099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 640099 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 640099 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 640099 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 640099 207854 640338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 640099 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 169568 633454 169888 633486
rect 169568 633218 169610 633454
rect 169846 633218 169888 633454
rect 169568 633134 169888 633218
rect 169568 632898 169610 633134
rect 169846 632898 169888 633134
rect 169568 632866 169888 632898
rect 200288 633454 200608 633486
rect 200288 633218 200330 633454
rect 200566 633218 200608 633454
rect 200288 633134 200608 633218
rect 200288 632898 200330 633134
rect 200566 632898 200608 633134
rect 200288 632866 200608 632898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 154208 615454 154528 615486
rect 154208 615218 154250 615454
rect 154486 615218 154528 615454
rect 154208 615134 154528 615218
rect 154208 614898 154250 615134
rect 154486 614898 154528 615134
rect 154208 614866 154528 614898
rect 184928 615454 185248 615486
rect 184928 615218 184970 615454
rect 185206 615218 185248 615454
rect 184928 615134 185248 615218
rect 184928 614898 184970 615134
rect 185206 614898 185248 615134
rect 184928 614866 185248 614898
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 169568 597454 169888 597486
rect 169568 597218 169610 597454
rect 169846 597218 169888 597454
rect 169568 597134 169888 597218
rect 169568 596898 169610 597134
rect 169846 596898 169888 597134
rect 169568 596866 169888 596898
rect 200288 597454 200608 597486
rect 200288 597218 200330 597454
rect 200566 597218 200608 597454
rect 200288 597134 200608 597218
rect 200288 596898 200330 597134
rect 200566 596898 200608 597134
rect 200288 596866 200608 596898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 562394 146414 578898
rect 154208 579454 154528 579486
rect 154208 579218 154250 579454
rect 154486 579218 154528 579454
rect 154208 579134 154528 579218
rect 154208 578898 154250 579134
rect 154486 578898 154528 579134
rect 154208 578866 154528 578898
rect 184928 579454 185248 579486
rect 184928 579218 184970 579454
rect 185206 579218 185248 579454
rect 184928 579134 185248 579218
rect 184928 578898 184970 579134
rect 185206 578898 185248 579134
rect 184928 578866 185248 578898
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 145794 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 146414 562394
rect 145794 562074 146414 562158
rect 145794 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 146414 562074
rect 145794 550000 146414 561838
rect 149514 564234 150134 573000
rect 149514 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 150134 564234
rect 149514 563914 150134 563998
rect 149514 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 150134 563914
rect 149514 550000 150134 563678
rect 153234 550894 153854 573000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 550000 153854 550338
rect 156954 554614 157574 573000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 550000 157574 554058
rect 163794 561454 164414 573000
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 550000 164414 560898
rect 167514 565174 168134 573000
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 550000 168134 564618
rect 171234 568894 171854 573000
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 550000 171854 568338
rect 174954 572614 175574 573000
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 550000 175574 572058
rect 181794 562394 182414 573000
rect 181794 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 182414 562394
rect 181794 562074 182414 562158
rect 181794 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 182414 562074
rect 181794 550000 182414 561838
rect 185514 564234 186134 573000
rect 185514 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 186134 564234
rect 185514 563914 186134 563998
rect 185514 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 186134 563914
rect 185514 550000 186134 563678
rect 189234 550894 189854 573000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 550000 189854 550338
rect 192954 554614 193574 573000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 550000 193574 554058
rect 199794 561454 200414 573000
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 550000 200414 560898
rect 203514 565174 204134 573000
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 550000 204134 564618
rect 207234 568894 207854 573000
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 550000 207854 568338
rect 210954 572614 211574 573000
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 550000 211574 572058
rect 217794 562394 218414 578898
rect 217794 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 218414 562394
rect 217794 562074 218414 562158
rect 217794 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 218414 562074
rect 217794 550000 218414 561838
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 564234 222134 582618
rect 221514 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 222134 564234
rect 221514 563914 222134 563998
rect 221514 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 222134 563914
rect 221514 550000 222134 563678
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 550000 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 550000 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 640099 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 640099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 640099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 640099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 640099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 640099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 640099 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 640099 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 640099 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 640099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 640099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 640099 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 640099 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 640099 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 640099 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 259568 633454 259888 633486
rect 259568 633218 259610 633454
rect 259846 633218 259888 633454
rect 259568 633134 259888 633218
rect 259568 632898 259610 633134
rect 259846 632898 259888 633134
rect 259568 632866 259888 632898
rect 290288 633454 290608 633486
rect 290288 633218 290330 633454
rect 290566 633218 290608 633454
rect 290288 633134 290608 633218
rect 290288 632898 290330 633134
rect 290566 632898 290608 633134
rect 290288 632866 290608 632898
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 244208 615454 244528 615486
rect 244208 615218 244250 615454
rect 244486 615218 244528 615454
rect 244208 615134 244528 615218
rect 244208 614898 244250 615134
rect 244486 614898 244528 615134
rect 244208 614866 244528 614898
rect 274928 615454 275248 615486
rect 274928 615218 274970 615454
rect 275206 615218 275248 615454
rect 274928 615134 275248 615218
rect 274928 614898 274970 615134
rect 275206 614898 275248 615134
rect 274928 614866 275248 614898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 259568 597454 259888 597486
rect 259568 597218 259610 597454
rect 259846 597218 259888 597454
rect 259568 597134 259888 597218
rect 259568 596898 259610 597134
rect 259846 596898 259888 597134
rect 259568 596866 259888 596898
rect 290288 597454 290608 597486
rect 290288 597218 290330 597454
rect 290566 597218 290608 597454
rect 290288 597134 290608 597218
rect 290288 596898 290330 597134
rect 290566 596898 290608 597134
rect 290288 596866 290608 596898
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 244208 579454 244528 579486
rect 244208 579218 244250 579454
rect 244486 579218 244528 579454
rect 244208 579134 244528 579218
rect 244208 578898 244250 579134
rect 244486 578898 244528 579134
rect 244208 578866 244528 578898
rect 274928 579454 275248 579486
rect 274928 579218 274970 579454
rect 275206 579218 275248 579454
rect 274928 579134 275248 579218
rect 274928 578898 274970 579134
rect 275206 578898 275248 579134
rect 274928 578866 275248 578898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 550000 236414 560898
rect 239514 565174 240134 573000
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 550000 240134 564618
rect 243234 568894 243854 573000
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 550000 243854 568338
rect 246954 572614 247574 573000
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 550000 247574 572058
rect 253794 562394 254414 573000
rect 253794 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 254414 562394
rect 253794 562074 254414 562158
rect 253794 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 254414 562074
rect 253794 550000 254414 561838
rect 257514 564234 258134 573000
rect 257514 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 258134 564234
rect 257514 563914 258134 563998
rect 257514 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 258134 563914
rect 257514 550000 258134 563678
rect 261234 550894 261854 573000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 550000 261854 550338
rect 264954 554614 265574 573000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 550000 265574 554058
rect 271794 561454 272414 573000
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 550000 272414 560898
rect 275514 565174 276134 573000
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 550000 276134 564618
rect 279234 568894 279854 573000
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 550000 279854 568338
rect 282954 572614 283574 573000
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 550000 283574 572058
rect 289794 562394 290414 573000
rect 289794 562158 289826 562394
rect 290062 562158 290146 562394
rect 290382 562158 290414 562394
rect 289794 562074 290414 562158
rect 289794 561838 289826 562074
rect 290062 561838 290146 562074
rect 290382 561838 290414 562074
rect 289794 550000 290414 561838
rect 293514 564234 294134 573000
rect 293514 563998 293546 564234
rect 293782 563998 293866 564234
rect 294102 563998 294134 564234
rect 293514 563914 294134 563998
rect 293514 563678 293546 563914
rect 293782 563678 293866 563914
rect 294102 563678 294134 563914
rect 293514 550000 294134 563678
rect 297234 550894 297854 573000
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 550000 297854 550338
rect 300954 554614 301574 573000
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 550000 301574 554058
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 64208 543454 64528 543486
rect 64208 543218 64250 543454
rect 64486 543218 64528 543454
rect 64208 543134 64528 543218
rect 64208 542898 64250 543134
rect 64486 542898 64528 543134
rect 64208 542866 64528 542898
rect 94928 543454 95248 543486
rect 94928 543218 94970 543454
rect 95206 543218 95248 543454
rect 94928 543134 95248 543218
rect 94928 542898 94970 543134
rect 95206 542898 95248 543134
rect 94928 542866 95248 542898
rect 125648 543454 125968 543486
rect 125648 543218 125690 543454
rect 125926 543218 125968 543454
rect 125648 543134 125968 543218
rect 125648 542898 125690 543134
rect 125926 542898 125968 543134
rect 125648 542866 125968 542898
rect 156368 543454 156688 543486
rect 156368 543218 156410 543454
rect 156646 543218 156688 543454
rect 156368 543134 156688 543218
rect 156368 542898 156410 543134
rect 156646 542898 156688 543134
rect 156368 542866 156688 542898
rect 187088 543454 187408 543486
rect 187088 543218 187130 543454
rect 187366 543218 187408 543454
rect 187088 543134 187408 543218
rect 187088 542898 187130 543134
rect 187366 542898 187408 543134
rect 187088 542866 187408 542898
rect 217808 543454 218128 543486
rect 217808 543218 217850 543454
rect 218086 543218 218128 543454
rect 217808 543134 218128 543218
rect 217808 542898 217850 543134
rect 218086 542898 218128 543134
rect 217808 542866 218128 542898
rect 248528 543454 248848 543486
rect 248528 543218 248570 543454
rect 248806 543218 248848 543454
rect 248528 543134 248848 543218
rect 248528 542898 248570 543134
rect 248806 542898 248848 543134
rect 248528 542866 248848 542898
rect 279248 543454 279568 543486
rect 279248 543218 279290 543454
rect 279526 543218 279568 543454
rect 279248 543134 279568 543218
rect 279248 542898 279290 543134
rect 279526 542898 279568 543134
rect 279248 542866 279568 542898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55075 485620 55141 485621
rect 55075 485556 55076 485620
rect 55140 485556 55141 485620
rect 55075 485555 55141 485556
rect 54891 466308 54957 466309
rect 54891 466244 54892 466308
rect 54956 466244 54957 466308
rect 54891 466243 54957 466244
rect 54707 466036 54773 466037
rect 54707 465972 54708 466036
rect 54772 465972 54773 466036
rect 54707 465971 54773 465972
rect 54339 254012 54405 254013
rect 54339 253948 54340 254012
rect 54404 253948 54405 254012
rect 54339 253947 54405 253948
rect 54710 59261 54770 465971
rect 54707 59260 54773 59261
rect 54707 59196 54708 59260
rect 54772 59196 54773 59260
rect 54707 59195 54773 59196
rect 54894 57629 54954 466243
rect 54891 57628 54957 57629
rect 54891 57564 54892 57628
rect 54956 57564 54957 57628
rect 54891 57563 54957 57564
rect 55078 56677 55138 485555
rect 55627 485484 55693 485485
rect 55627 485420 55628 485484
rect 55692 485420 55693 485484
rect 55627 485419 55693 485420
rect 55443 468756 55509 468757
rect 55443 468692 55444 468756
rect 55508 468692 55509 468756
rect 55443 468691 55509 468692
rect 55075 56676 55141 56677
rect 55075 56612 55076 56676
rect 55140 56612 55141 56676
rect 55075 56611 55141 56612
rect 53603 56404 53669 56405
rect 53603 56340 53604 56404
rect 53668 56340 53669 56404
rect 53603 56339 53669 56340
rect 51763 56268 51829 56269
rect 51763 56204 51764 56268
rect 51828 56204 51829 56268
rect 51763 56203 51829 56204
rect 50659 55044 50725 55045
rect 50659 54980 50660 55044
rect 50724 54980 50725 55044
rect 50659 54979 50725 54980
rect 55446 54909 55506 468691
rect 55630 59125 55690 485419
rect 55794 453454 56414 488898
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 206139 486436 206205 486437
rect 206139 486372 206140 486436
rect 206204 486372 206205 486436
rect 206139 486371 206205 486372
rect 59307 485756 59373 485757
rect 59307 485692 59308 485756
rect 59372 485692 59373 485756
rect 59307 485691 59373 485692
rect 57835 485076 57901 485077
rect 57835 485012 57836 485076
rect 57900 485012 57901 485076
rect 57835 485011 57901 485012
rect 57099 482628 57165 482629
rect 57099 482564 57100 482628
rect 57164 482564 57165 482628
rect 57099 482563 57165 482564
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57102 379133 57162 482563
rect 57651 479908 57717 479909
rect 57651 479844 57652 479908
rect 57716 479844 57717 479908
rect 57651 479843 57717 479844
rect 57467 477324 57533 477325
rect 57467 477260 57468 477324
rect 57532 477260 57533 477324
rect 57467 477259 57533 477260
rect 57470 388517 57530 477259
rect 57467 388516 57533 388517
rect 57467 388452 57468 388516
rect 57532 388452 57533 388516
rect 57467 388451 57533 388452
rect 57099 379132 57165 379133
rect 57099 379068 57100 379132
rect 57164 379068 57165 379132
rect 57099 379067 57165 379068
rect 57467 378044 57533 378045
rect 57467 377980 57468 378044
rect 57532 377980 57533 378044
rect 57467 377979 57533 377980
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 57470 273325 57530 377979
rect 57467 273324 57533 273325
rect 57467 273260 57468 273324
rect 57532 273260 57533 273324
rect 57467 273259 57533 273260
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57654 270333 57714 479843
rect 57651 270332 57717 270333
rect 57651 270268 57652 270332
rect 57716 270268 57717 270332
rect 57651 270267 57717 270268
rect 57651 252516 57717 252517
rect 57651 252452 57652 252516
rect 57716 252452 57717 252516
rect 57651 252451 57717 252452
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57654 164117 57714 252451
rect 57838 166973 57898 485011
rect 59123 484940 59189 484941
rect 59123 484876 59124 484940
rect 59188 484876 59189 484940
rect 59123 484875 59189 484876
rect 58939 468348 59005 468349
rect 58939 468284 58940 468348
rect 59004 468284 59005 468348
rect 58939 468283 59005 468284
rect 58571 466444 58637 466445
rect 58571 466380 58572 466444
rect 58636 466380 58637 466444
rect 58571 466379 58637 466380
rect 57835 166972 57901 166973
rect 57835 166908 57836 166972
rect 57900 166908 57901 166972
rect 57835 166907 57901 166908
rect 57651 164116 57717 164117
rect 57651 164052 57652 164116
rect 57716 164052 57717 164116
rect 57651 164051 57717 164052
rect 57654 161490 57714 164051
rect 57654 161430 57898 161490
rect 57651 147796 57717 147797
rect 57651 147732 57652 147796
rect 57716 147732 57717 147796
rect 57651 147731 57717 147732
rect 57467 140860 57533 140861
rect 57467 140796 57468 140860
rect 57532 140796 57533 140860
rect 57467 140795 57533 140796
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55627 59124 55693 59125
rect 55627 59060 55628 59124
rect 55692 59060 55693 59124
rect 55627 59059 55693 59060
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55443 54908 55509 54909
rect 55443 54844 55444 54908
rect 55508 54844 55509 54908
rect 55443 54843 55509 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57470 56133 57530 140795
rect 57654 59533 57714 147731
rect 57651 59532 57717 59533
rect 57651 59468 57652 59532
rect 57716 59468 57717 59532
rect 57651 59467 57717 59468
rect 57838 57493 57898 161430
rect 57835 57492 57901 57493
rect 57835 57428 57836 57492
rect 57900 57428 57901 57492
rect 57835 57427 57901 57428
rect 58574 57357 58634 466379
rect 58755 465628 58821 465629
rect 58755 465564 58756 465628
rect 58820 465564 58821 465628
rect 58755 465563 58821 465564
rect 58571 57356 58637 57357
rect 58571 57292 58572 57356
rect 58636 57292 58637 57356
rect 58571 57291 58637 57292
rect 58758 57085 58818 465563
rect 58942 57221 59002 468283
rect 59126 58445 59186 484875
rect 59310 58717 59370 485691
rect 59514 476114 60134 486000
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 60134 476114
rect 59514 475794 60134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 60134 475794
rect 59514 466308 60134 475558
rect 63234 477954 63854 486000
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 63854 477954
rect 63234 477634 63854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 63854 477634
rect 60227 469164 60293 469165
rect 60227 469100 60228 469164
rect 60292 469100 60293 469164
rect 60227 469099 60293 469100
rect 60230 464810 60290 469099
rect 63234 466308 63854 477398
rect 66954 481674 67574 486000
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 67574 481674
rect 66954 481354 67574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 67574 481354
rect 66954 466308 67574 481118
rect 73794 471454 74414 486000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 466308 74414 470898
rect 77514 475174 78134 486000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 466308 78134 474618
rect 81234 478894 81854 486000
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 466308 81854 478338
rect 84954 482614 85574 486000
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 466308 85574 482058
rect 91794 472394 92414 486000
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 92414 472394
rect 91794 472074 92414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 92414 472074
rect 91794 466308 92414 471838
rect 95514 476114 96134 486000
rect 95514 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 96134 476114
rect 95514 475794 96134 475878
rect 95514 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 96134 475794
rect 95514 466308 96134 475558
rect 99234 477954 99854 486000
rect 99234 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 99854 477954
rect 99234 477634 99854 477718
rect 99234 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 99854 477634
rect 99234 466308 99854 477398
rect 102954 481674 103574 486000
rect 102954 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 103574 481674
rect 102954 481354 103574 481438
rect 102954 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 103574 481354
rect 102954 466308 103574 481118
rect 109794 471454 110414 486000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 466308 110414 470898
rect 113514 475174 114134 486000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 466308 114134 474618
rect 117234 478894 117854 486000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 466308 117854 478338
rect 120954 482614 121574 486000
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 466308 121574 482058
rect 127794 472394 128414 486000
rect 127794 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 128414 472394
rect 127794 472074 128414 472158
rect 127794 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 128414 472074
rect 127794 466308 128414 471838
rect 131514 476114 132134 486000
rect 131514 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 132134 476114
rect 131514 475794 132134 475878
rect 131514 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 132134 475794
rect 131514 466308 132134 475558
rect 135234 477954 135854 486000
rect 135234 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 135854 477954
rect 135234 477634 135854 477718
rect 135234 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 135854 477634
rect 135234 466308 135854 477398
rect 138954 481674 139574 486000
rect 138954 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 139574 481674
rect 138954 481354 139574 481438
rect 138954 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 139574 481354
rect 138954 466308 139574 481118
rect 145794 471454 146414 486000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 466308 146414 470898
rect 149514 475174 150134 486000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 466308 150134 474618
rect 153234 478894 153854 486000
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 466308 153854 478338
rect 156954 482614 157574 486000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 466308 157574 482058
rect 163794 472394 164414 486000
rect 163794 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 164414 472394
rect 163794 472074 164414 472158
rect 163794 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 164414 472074
rect 163794 466308 164414 471838
rect 167514 476114 168134 486000
rect 167514 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 168134 476114
rect 167514 475794 168134 475878
rect 167514 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 168134 475794
rect 167514 466308 168134 475558
rect 171234 477954 171854 486000
rect 171234 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 171854 477954
rect 171234 477634 171854 477718
rect 171234 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 171854 477634
rect 171234 466308 171854 477398
rect 174954 481674 175574 486000
rect 174954 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 175574 481674
rect 174954 481354 175574 481438
rect 174954 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 175574 481354
rect 174954 466308 175574 481118
rect 181794 471454 182414 486000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 466988 179709 466989
rect 179643 466924 179644 466988
rect 179708 466924 179709 466988
rect 179643 466923 179709 466924
rect 178355 466580 178421 466581
rect 178355 466516 178356 466580
rect 178420 466516 178421 466580
rect 178355 466515 178421 466516
rect 59862 464750 60290 464810
rect 178358 464810 178418 466515
rect 179646 464810 179706 466923
rect 181794 466308 182414 470898
rect 185514 475174 186134 486000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 466308 186134 474618
rect 189234 478894 189854 486000
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 466308 189854 478338
rect 192954 482614 193574 486000
rect 199331 485756 199397 485757
rect 199331 485692 199332 485756
rect 199396 485692 199397 485756
rect 199331 485691 199397 485692
rect 198043 485620 198109 485621
rect 198043 485556 198044 485620
rect 198108 485556 198109 485620
rect 198043 485555 198109 485556
rect 196571 485484 196637 485485
rect 196571 485420 196572 485484
rect 196636 485420 196637 485484
rect 196571 485419 196637 485420
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190867 466580 190933 466581
rect 190867 466516 190868 466580
rect 190932 466516 190933 466580
rect 190867 466515 190933 466516
rect 190870 464810 190930 466515
rect 192954 466308 193574 482058
rect 178358 464750 178524 464810
rect 179646 464750 179748 464810
rect 59862 379810 59922 464750
rect 178464 464202 178524 464750
rect 179688 464202 179748 464750
rect 190840 464750 190930 464810
rect 190840 464202 190900 464750
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 76056 380493 76116 381106
rect 76051 380492 76117 380493
rect 76051 380428 76052 380492
rect 76116 380428 76117 380492
rect 77144 380490 77204 381106
rect 78232 380490 78292 381106
rect 79592 380490 79652 381106
rect 80544 380490 80604 381106
rect 81768 380490 81828 381106
rect 77144 380430 77218 380490
rect 78232 380430 78322 380490
rect 76051 380427 76117 380428
rect 59862 379750 60290 379810
rect 59514 368114 60134 379000
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 60134 368114
rect 59514 367794 60134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 60134 367794
rect 59514 359308 60134 367558
rect 60230 358730 60290 379750
rect 63234 369954 63854 379000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 359308 63854 369398
rect 66954 373674 67574 379000
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 67574 373674
rect 66954 373354 67574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 67574 373354
rect 66954 359308 67574 373118
rect 73794 363454 74414 379000
rect 77158 378997 77218 380430
rect 78262 379133 78322 380430
rect 79550 380430 79652 380490
rect 80470 380430 80604 380490
rect 81758 380430 81828 380490
rect 83128 380490 83188 381106
rect 84216 380490 84276 381106
rect 85440 380490 85500 381106
rect 83128 380430 83290 380490
rect 84216 380430 84394 380490
rect 78259 379132 78325 379133
rect 78259 379068 78260 379132
rect 78324 379068 78325 379132
rect 78259 379067 78325 379068
rect 77155 378996 77221 378997
rect 77155 378932 77156 378996
rect 77220 378932 77221 378996
rect 77155 378931 77221 378932
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 359308 74414 362898
rect 77514 367174 78134 379000
rect 79550 378861 79610 380430
rect 80470 379269 80530 380430
rect 81758 379405 81818 380430
rect 81755 379404 81821 379405
rect 81755 379340 81756 379404
rect 81820 379340 81821 379404
rect 81755 379339 81821 379340
rect 81939 379404 82005 379405
rect 81939 379340 81940 379404
rect 82004 379340 82005 379404
rect 81939 379339 82005 379340
rect 80467 379268 80533 379269
rect 80467 379204 80468 379268
rect 80532 379204 80533 379268
rect 80467 379203 80533 379204
rect 79547 378860 79613 378861
rect 79547 378796 79548 378860
rect 79612 378796 79613 378860
rect 79547 378795 79613 378796
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 359308 78134 366618
rect 81234 370894 81854 379000
rect 81942 378725 82002 379339
rect 83230 378861 83290 380430
rect 83227 378860 83293 378861
rect 83227 378796 83228 378860
rect 83292 378796 83293 378860
rect 83227 378795 83293 378796
rect 81939 378724 82005 378725
rect 81939 378660 81940 378724
rect 82004 378660 82005 378724
rect 81939 378659 82005 378660
rect 84334 378181 84394 380430
rect 85438 380430 85500 380490
rect 86528 380490 86588 381106
rect 87616 380490 87676 381106
rect 88296 380490 88356 381106
rect 88704 380490 88764 381106
rect 90064 380490 90124 381106
rect 86528 380430 86602 380490
rect 87616 380430 87706 380490
rect 88296 380430 88442 380490
rect 88704 380430 88810 380490
rect 85438 379405 85498 380430
rect 86542 379405 86602 380430
rect 87646 379405 87706 380430
rect 88382 379405 88442 380430
rect 88750 379405 88810 380430
rect 90038 380430 90124 380490
rect 90744 380490 90804 381106
rect 91288 380490 91348 381106
rect 92376 380490 92436 381106
rect 93464 380490 93524 381106
rect 90744 380430 90834 380490
rect 91288 380430 91386 380490
rect 92376 380430 92490 380490
rect 90038 379405 90098 380430
rect 90774 379405 90834 380430
rect 91326 379405 91386 380430
rect 92430 379405 92490 380430
rect 93350 380430 93524 380490
rect 93600 380490 93660 381106
rect 94552 380490 94612 381106
rect 95912 380490 95972 381106
rect 96048 380490 96108 381106
rect 97000 380490 97060 381106
rect 98088 380490 98148 381106
rect 98496 380490 98556 381106
rect 99448 380490 99508 381106
rect 93600 380430 93778 380490
rect 94552 380430 94698 380490
rect 95912 380430 95986 380490
rect 96048 380430 96170 380490
rect 97000 380430 97090 380490
rect 98088 380430 98194 380490
rect 98496 380430 98562 380490
rect 93350 379405 93410 380430
rect 85435 379404 85501 379405
rect 85435 379340 85436 379404
rect 85500 379340 85501 379404
rect 85435 379339 85501 379340
rect 86539 379404 86605 379405
rect 86539 379340 86540 379404
rect 86604 379340 86605 379404
rect 86539 379339 86605 379340
rect 87643 379404 87709 379405
rect 87643 379340 87644 379404
rect 87708 379340 87709 379404
rect 87643 379339 87709 379340
rect 88379 379404 88445 379405
rect 88379 379340 88380 379404
rect 88444 379340 88445 379404
rect 88379 379339 88445 379340
rect 88747 379404 88813 379405
rect 88747 379340 88748 379404
rect 88812 379340 88813 379404
rect 88747 379339 88813 379340
rect 90035 379404 90101 379405
rect 90035 379340 90036 379404
rect 90100 379340 90101 379404
rect 90035 379339 90101 379340
rect 90771 379404 90837 379405
rect 90771 379340 90772 379404
rect 90836 379340 90837 379404
rect 90771 379339 90837 379340
rect 91323 379404 91389 379405
rect 91323 379340 91324 379404
rect 91388 379340 91389 379404
rect 91323 379339 91389 379340
rect 92427 379404 92493 379405
rect 92427 379340 92428 379404
rect 92492 379340 92493 379404
rect 92427 379339 92493 379340
rect 93347 379404 93413 379405
rect 93347 379340 93348 379404
rect 93412 379340 93413 379404
rect 93347 379339 93413 379340
rect 93718 379269 93778 380430
rect 93715 379268 93781 379269
rect 93715 379204 93716 379268
rect 93780 379204 93781 379268
rect 93715 379203 93781 379204
rect 84331 378180 84397 378181
rect 84331 378116 84332 378180
rect 84396 378116 84397 378180
rect 84331 378115 84397 378116
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 359308 81854 370338
rect 84954 374614 85574 379000
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 359308 85574 374058
rect 91794 364394 92414 379000
rect 94638 378997 94698 380430
rect 95926 379269 95986 380430
rect 96110 379405 96170 380430
rect 96107 379404 96173 379405
rect 96107 379340 96108 379404
rect 96172 379340 96173 379404
rect 96107 379339 96173 379340
rect 95923 379268 95989 379269
rect 95923 379204 95924 379268
rect 95988 379204 95989 379268
rect 95923 379203 95989 379204
rect 94635 378996 94701 378997
rect 94635 378932 94636 378996
rect 94700 378932 94701 378996
rect 94635 378931 94701 378932
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 359308 92414 363838
rect 95514 368114 96134 379000
rect 97030 378589 97090 380430
rect 98134 379405 98194 380430
rect 98502 379405 98562 380430
rect 99422 380430 99508 380490
rect 100672 380490 100732 381106
rect 101080 380490 101140 381106
rect 100672 380430 100770 380490
rect 98131 379404 98197 379405
rect 98131 379340 98132 379404
rect 98196 379340 98197 379404
rect 98131 379339 98197 379340
rect 98499 379404 98565 379405
rect 98499 379340 98500 379404
rect 98564 379340 98565 379404
rect 98499 379339 98565 379340
rect 99422 379269 99482 380430
rect 99419 379268 99485 379269
rect 99419 379204 99420 379268
rect 99484 379204 99485 379268
rect 99419 379203 99485 379204
rect 97027 378588 97093 378589
rect 97027 378524 97028 378588
rect 97092 378524 97093 378588
rect 97027 378523 97093 378524
rect 95514 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 96134 368114
rect 95514 367794 96134 367878
rect 95514 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 96134 367794
rect 95514 359308 96134 367558
rect 99234 369954 99854 379000
rect 100710 378589 100770 380430
rect 101078 380430 101140 380490
rect 101760 380490 101820 381106
rect 102848 380490 102908 381106
rect 103528 380490 103588 381106
rect 101760 380430 101874 380490
rect 102848 380430 102978 380490
rect 101078 379405 101138 380430
rect 101075 379404 101141 379405
rect 101075 379340 101076 379404
rect 101140 379340 101141 379404
rect 101075 379339 101141 379340
rect 100707 378588 100773 378589
rect 100707 378524 100708 378588
rect 100772 378524 100773 378588
rect 100707 378523 100773 378524
rect 101814 378181 101874 380430
rect 102918 379269 102978 380430
rect 103286 380430 103588 380490
rect 103936 380490 103996 381106
rect 105296 380490 105356 381106
rect 105976 380490 106036 381106
rect 103936 380430 104082 380490
rect 105296 380430 105370 380490
rect 103286 379405 103346 380430
rect 103283 379404 103349 379405
rect 103283 379340 103284 379404
rect 103348 379340 103349 379404
rect 103283 379339 103349 379340
rect 102915 379268 102981 379269
rect 102915 379204 102916 379268
rect 102980 379204 102981 379268
rect 102915 379203 102981 379204
rect 101811 378180 101877 378181
rect 101811 378116 101812 378180
rect 101876 378116 101877 378180
rect 101811 378115 101877 378116
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 359308 99854 369398
rect 102954 373674 103574 379000
rect 104022 378181 104082 380430
rect 105310 378453 105370 380430
rect 105862 380430 106036 380490
rect 106384 380490 106444 381106
rect 107608 380490 107668 381106
rect 108288 380490 108348 381106
rect 106384 380430 106474 380490
rect 105862 379405 105922 380430
rect 105859 379404 105925 379405
rect 105859 379340 105860 379404
rect 105924 379340 105925 379404
rect 105859 379339 105925 379340
rect 105307 378452 105373 378453
rect 105307 378388 105308 378452
rect 105372 378388 105373 378452
rect 105307 378387 105373 378388
rect 106414 378181 106474 380430
rect 107518 380430 107668 380490
rect 108254 380430 108348 380490
rect 108696 380490 108756 381106
rect 109784 380490 109844 381106
rect 111008 380765 111068 381106
rect 111005 380764 111071 380765
rect 111005 380700 111006 380764
rect 111070 380700 111071 380764
rect 111005 380699 111071 380700
rect 108696 380430 108866 380490
rect 107518 378181 107578 380430
rect 108254 379405 108314 380430
rect 108806 379405 108866 380430
rect 109726 380430 109844 380490
rect 111144 380490 111204 381106
rect 112232 380490 112292 381106
rect 113320 380490 113380 381106
rect 113592 380765 113652 381106
rect 113589 380764 113655 380765
rect 113589 380700 113590 380764
rect 113654 380700 113655 380764
rect 113589 380699 113655 380700
rect 114408 380490 114468 381106
rect 115768 380490 115828 381106
rect 116040 380765 116100 381106
rect 116037 380764 116103 380765
rect 116037 380700 116038 380764
rect 116102 380700 116103 380764
rect 116037 380699 116103 380700
rect 116992 380490 117052 381106
rect 118080 380490 118140 381106
rect 118488 380765 118548 381106
rect 118485 380764 118551 380765
rect 118485 380700 118486 380764
rect 118550 380700 118551 380764
rect 118485 380699 118551 380700
rect 119168 380490 119228 381106
rect 120936 380765 120996 381106
rect 123520 380765 123580 381106
rect 125968 380765 126028 381106
rect 120933 380764 120999 380765
rect 120933 380700 120934 380764
rect 120998 380700 120999 380764
rect 120933 380699 120999 380700
rect 123517 380764 123583 380765
rect 123517 380700 123518 380764
rect 123582 380700 123583 380764
rect 123517 380699 123583 380700
rect 125965 380764 126031 380765
rect 125965 380700 125966 380764
rect 126030 380700 126031 380764
rect 125965 380699 126031 380700
rect 111144 380430 111258 380490
rect 112232 380430 112362 380490
rect 113320 380430 113466 380490
rect 114408 380430 114570 380490
rect 115768 380430 115858 380490
rect 116992 380430 117146 380490
rect 118080 380430 118250 380490
rect 108251 379404 108317 379405
rect 108251 379340 108252 379404
rect 108316 379340 108317 379404
rect 108251 379339 108317 379340
rect 108803 379404 108869 379405
rect 108803 379340 108804 379404
rect 108868 379340 108869 379404
rect 108803 379339 108869 379340
rect 109726 379269 109786 380430
rect 111198 379405 111258 380430
rect 112302 379405 112362 380430
rect 113406 379405 113466 380430
rect 114510 379405 114570 380430
rect 115798 379405 115858 380430
rect 111195 379404 111261 379405
rect 111195 379340 111196 379404
rect 111260 379340 111261 379404
rect 111195 379339 111261 379340
rect 112299 379404 112365 379405
rect 112299 379340 112300 379404
rect 112364 379340 112365 379404
rect 112299 379339 112365 379340
rect 113403 379404 113469 379405
rect 113403 379340 113404 379404
rect 113468 379340 113469 379404
rect 113403 379339 113469 379340
rect 114507 379404 114573 379405
rect 114507 379340 114508 379404
rect 114572 379340 114573 379404
rect 114507 379339 114573 379340
rect 115795 379404 115861 379405
rect 115795 379340 115796 379404
rect 115860 379340 115861 379404
rect 115795 379339 115861 379340
rect 109723 379268 109789 379269
rect 109723 379204 109724 379268
rect 109788 379204 109789 379268
rect 109723 379203 109789 379204
rect 104019 378180 104085 378181
rect 104019 378116 104020 378180
rect 104084 378116 104085 378180
rect 104019 378115 104085 378116
rect 106411 378180 106477 378181
rect 106411 378116 106412 378180
rect 106476 378116 106477 378180
rect 106411 378115 106477 378116
rect 107515 378180 107581 378181
rect 107515 378116 107516 378180
rect 107580 378116 107581 378180
rect 107515 378115 107581 378116
rect 102954 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 103574 373674
rect 102954 373354 103574 373438
rect 102954 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 103574 373354
rect 102954 359308 103574 373118
rect 109794 363454 110414 379000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 359308 110414 362898
rect 113514 367174 114134 379000
rect 117086 378181 117146 380430
rect 117083 378180 117149 378181
rect 117083 378116 117084 378180
rect 117148 378116 117149 378180
rect 117083 378115 117149 378116
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 359308 114134 366618
rect 117234 370894 117854 379000
rect 118190 378589 118250 380430
rect 119110 380430 119228 380490
rect 128280 380490 128340 381106
rect 131000 380765 131060 381106
rect 133448 380765 133508 381106
rect 130997 380764 131063 380765
rect 130997 380700 130998 380764
rect 131062 380700 131063 380764
rect 130997 380699 131063 380700
rect 133445 380764 133511 380765
rect 133445 380700 133446 380764
rect 133510 380700 133511 380764
rect 133445 380699 133511 380700
rect 135896 380490 135956 381106
rect 138480 380490 138540 381106
rect 140928 380765 140988 381106
rect 143512 380765 143572 381106
rect 145960 380765 146020 381106
rect 140925 380764 140991 380765
rect 140925 380700 140926 380764
rect 140990 380700 140991 380764
rect 140925 380699 140991 380700
rect 143509 380764 143575 380765
rect 143509 380700 143510 380764
rect 143574 380700 143575 380764
rect 143509 380699 143575 380700
rect 145957 380764 146023 380765
rect 145957 380700 145958 380764
rect 146022 380700 146023 380764
rect 145957 380699 146023 380700
rect 128280 380430 128370 380490
rect 119110 380357 119170 380430
rect 119107 380356 119173 380357
rect 119107 380292 119108 380356
rect 119172 380292 119173 380356
rect 119107 380291 119173 380292
rect 128310 380221 128370 380430
rect 135854 380430 135956 380490
rect 138430 380430 138540 380490
rect 148544 380490 148604 381106
rect 150992 380490 151052 381106
rect 148544 380430 148610 380490
rect 128307 380220 128373 380221
rect 128307 380156 128308 380220
rect 128372 380156 128373 380220
rect 128307 380155 128373 380156
rect 135854 379405 135914 380430
rect 138430 379405 138490 380430
rect 135851 379404 135917 379405
rect 135851 379340 135852 379404
rect 135916 379340 135917 379404
rect 135851 379339 135917 379340
rect 138427 379404 138493 379405
rect 138427 379340 138428 379404
rect 138492 379340 138493 379404
rect 138427 379339 138493 379340
rect 118187 378588 118253 378589
rect 118187 378524 118188 378588
rect 118252 378524 118253 378588
rect 118187 378523 118253 378524
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 359308 117854 370338
rect 120954 374614 121574 379000
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 359308 121574 374058
rect 127794 364394 128414 379000
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 359308 128414 363838
rect 131514 368114 132134 379000
rect 131514 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 132134 368114
rect 131514 367794 132134 367878
rect 131514 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 132134 367794
rect 131514 359308 132134 367558
rect 135234 369954 135854 379000
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 359308 135854 369398
rect 138954 373674 139574 379000
rect 138954 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 139574 373674
rect 138954 373354 139574 373438
rect 138954 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 139574 373354
rect 138954 359308 139574 373118
rect 145794 363454 146414 379000
rect 148550 378997 148610 380430
rect 150942 380430 151052 380490
rect 153440 380490 153500 381106
rect 155888 380765 155948 381106
rect 158472 380765 158532 381106
rect 160920 380765 160980 381106
rect 163368 380765 163428 381106
rect 165952 380765 166012 381106
rect 155885 380764 155951 380765
rect 155885 380700 155886 380764
rect 155950 380700 155951 380764
rect 155885 380699 155951 380700
rect 158469 380764 158535 380765
rect 158469 380700 158470 380764
rect 158534 380700 158535 380764
rect 158469 380699 158535 380700
rect 160917 380764 160983 380765
rect 160917 380700 160918 380764
rect 160982 380700 160983 380764
rect 160917 380699 160983 380700
rect 163365 380764 163431 380765
rect 163365 380700 163366 380764
rect 163430 380700 163431 380764
rect 163365 380699 163431 380700
rect 165949 380764 166015 380765
rect 165949 380700 165950 380764
rect 166014 380700 166015 380764
rect 165949 380699 166015 380700
rect 183224 380490 183284 381106
rect 153440 380430 153578 380490
rect 150942 379405 151002 380430
rect 153518 379405 153578 380430
rect 183142 380430 183284 380490
rect 183360 380490 183420 381106
rect 183360 380430 183570 380490
rect 150939 379404 151005 379405
rect 150939 379340 150940 379404
rect 151004 379340 151005 379404
rect 150939 379339 151005 379340
rect 153515 379404 153581 379405
rect 153515 379340 153516 379404
rect 153580 379340 153581 379404
rect 153515 379339 153581 379340
rect 148547 378996 148613 378997
rect 148547 378932 148548 378996
rect 148612 378932 148613 378996
rect 148547 378931 148613 378932
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 359308 146414 362898
rect 149514 367174 150134 379000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 359308 150134 366618
rect 153234 370894 153854 379000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 359308 153854 370338
rect 156954 374614 157574 379000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 359308 157574 374058
rect 163794 364394 164414 379000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 359308 164414 363838
rect 167514 368114 168134 379000
rect 167514 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 168134 368114
rect 167514 367794 168134 367878
rect 167514 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 168134 367794
rect 167514 359308 168134 367558
rect 171234 369954 171854 379000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 359308 171854 369398
rect 174954 373674 175574 379000
rect 174954 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 175574 373674
rect 174954 373354 175574 373438
rect 174954 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 175574 373354
rect 174954 359308 175574 373118
rect 181794 363454 182414 379000
rect 183142 378997 183202 380430
rect 183139 378996 183205 378997
rect 183139 378932 183140 378996
rect 183204 378932 183205 378996
rect 183139 378931 183205 378932
rect 183510 378453 183570 380430
rect 183507 378452 183573 378453
rect 183507 378388 183508 378452
rect 183572 378388 183573 378452
rect 183507 378387 183573 378388
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 359308 182414 362898
rect 185514 367174 186134 379000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 359308 186134 366618
rect 189234 370894 189854 379000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 359308 189854 370338
rect 192954 374614 193574 379000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 359308 193574 374058
rect 178539 358868 178605 358869
rect 178539 358804 178540 358868
rect 178604 358804 178605 358868
rect 178539 358803 178605 358804
rect 179643 358868 179709 358869
rect 179643 358804 179644 358868
rect 179708 358804 179709 358868
rect 179643 358803 179709 358804
rect 190867 358868 190933 358869
rect 190867 358804 190868 358868
rect 190932 358804 190933 358868
rect 190867 358803 190933 358804
rect 59862 358670 60290 358730
rect 59862 272370 59922 358670
rect 178542 358050 178602 358803
rect 178464 357990 178602 358050
rect 179646 358050 179706 358803
rect 190870 358050 190930 358803
rect 179646 357990 179748 358050
rect 178464 357202 178524 357990
rect 179688 357202 179748 357990
rect 190840 357990 190930 358050
rect 190840 357202 190900 357990
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 76056 273730 76116 274040
rect 76054 273670 76116 273730
rect 77144 273730 77204 274040
rect 78232 273730 78292 274040
rect 79592 273730 79652 274040
rect 80544 273730 80604 274040
rect 77144 273670 77218 273730
rect 78232 273670 78322 273730
rect 76054 273189 76114 273670
rect 77158 273189 77218 273670
rect 76051 273188 76117 273189
rect 76051 273124 76052 273188
rect 76116 273124 76117 273188
rect 76051 273123 76117 273124
rect 77155 273188 77221 273189
rect 77155 273124 77156 273188
rect 77220 273124 77221 273188
rect 77155 273123 77221 273124
rect 59862 272310 60290 272370
rect 59514 260114 60134 272000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 252308 60134 259558
rect 60230 251970 60290 272310
rect 63234 261954 63854 272000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 252308 63854 261398
rect 66954 265674 67574 272000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 252308 67574 265118
rect 73794 255454 74414 272000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 252308 74414 254898
rect 77514 259174 78134 272000
rect 78262 271013 78322 273670
rect 79550 273670 79652 273730
rect 80470 273670 80604 273730
rect 81768 273730 81828 274040
rect 83128 273730 83188 274040
rect 84216 273730 84276 274040
rect 85440 273730 85500 274040
rect 81768 273670 82002 273730
rect 79550 271693 79610 273670
rect 79547 271692 79613 271693
rect 79547 271628 79548 271692
rect 79612 271628 79613 271692
rect 79547 271627 79613 271628
rect 78259 271012 78325 271013
rect 78259 270948 78260 271012
rect 78324 270948 78325 271012
rect 78259 270947 78325 270948
rect 80470 270877 80530 273670
rect 80467 270876 80533 270877
rect 80467 270812 80468 270876
rect 80532 270812 80533 270876
rect 80467 270811 80533 270812
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 252308 78134 258618
rect 81234 262894 81854 272000
rect 81942 271285 82002 273670
rect 83046 273670 83188 273730
rect 83966 273670 84276 273730
rect 84702 273670 85500 273730
rect 86528 273730 86588 274040
rect 87616 273730 87676 274040
rect 88296 273730 88356 274040
rect 88704 273730 88764 274040
rect 90064 273730 90124 274040
rect 86528 273670 86602 273730
rect 87616 273670 87706 273730
rect 88296 273670 88442 273730
rect 88704 273670 88810 273730
rect 83046 273189 83106 273670
rect 83043 273188 83109 273189
rect 83043 273124 83044 273188
rect 83108 273124 83109 273188
rect 83043 273123 83109 273124
rect 83966 271829 84026 273670
rect 83963 271828 84029 271829
rect 83963 271764 83964 271828
rect 84028 271764 84029 271828
rect 83963 271763 84029 271764
rect 84702 271693 84762 273670
rect 84699 271692 84765 271693
rect 84699 271628 84700 271692
rect 84764 271628 84765 271692
rect 84699 271627 84765 271628
rect 81939 271284 82005 271285
rect 81939 271220 81940 271284
rect 82004 271220 82005 271284
rect 81939 271219 82005 271220
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 252308 81854 262338
rect 84954 266614 85574 272000
rect 86542 270605 86602 273670
rect 87646 272373 87706 273670
rect 87643 272372 87709 272373
rect 87643 272308 87644 272372
rect 87708 272308 87709 272372
rect 87643 272307 87709 272308
rect 88382 271285 88442 273670
rect 88379 271284 88445 271285
rect 88379 271220 88380 271284
rect 88444 271220 88445 271284
rect 88379 271219 88445 271220
rect 88750 270877 88810 273670
rect 90038 273670 90124 273730
rect 90744 273730 90804 274040
rect 91288 273730 91348 274040
rect 92376 273730 92436 274040
rect 93464 273730 93524 274040
rect 90744 273670 90834 273730
rect 91288 273670 91386 273730
rect 88747 270876 88813 270877
rect 88747 270812 88748 270876
rect 88812 270812 88813 270876
rect 88747 270811 88813 270812
rect 90038 270741 90098 273670
rect 90774 273189 90834 273670
rect 90771 273188 90837 273189
rect 90771 273124 90772 273188
rect 90836 273124 90837 273188
rect 90771 273123 90837 273124
rect 90035 270740 90101 270741
rect 90035 270676 90036 270740
rect 90100 270676 90101 270740
rect 90035 270675 90101 270676
rect 91326 270605 91386 273670
rect 91510 273670 92436 273730
rect 93350 273670 93524 273730
rect 93600 273730 93660 274040
rect 94552 273730 94612 274040
rect 93600 273670 93778 273730
rect 86539 270604 86605 270605
rect 86539 270540 86540 270604
rect 86604 270540 86605 270604
rect 86539 270539 86605 270540
rect 91323 270604 91389 270605
rect 91323 270540 91324 270604
rect 91388 270540 91389 270604
rect 91323 270539 91389 270540
rect 91510 270469 91570 273670
rect 91507 270468 91573 270469
rect 91507 270404 91508 270468
rect 91572 270404 91573 270468
rect 91507 270403 91573 270404
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 252308 85574 266058
rect 91794 256394 92414 272000
rect 93350 270741 93410 273670
rect 93718 273189 93778 273670
rect 94454 273670 94612 273730
rect 95912 273730 95972 274040
rect 96048 273730 96108 274040
rect 97000 273730 97060 274040
rect 98088 273730 98148 274040
rect 98496 273730 98556 274040
rect 99448 273730 99508 274040
rect 95912 273670 95986 273730
rect 96048 273670 96170 273730
rect 97000 273670 97090 273730
rect 98088 273670 98194 273730
rect 98496 273670 98562 273730
rect 93715 273188 93781 273189
rect 93715 273124 93716 273188
rect 93780 273124 93781 273188
rect 93715 273123 93781 273124
rect 94454 272373 94514 273670
rect 95926 273189 95986 273670
rect 95923 273188 95989 273189
rect 95923 273124 95924 273188
rect 95988 273124 95989 273188
rect 95923 273123 95989 273124
rect 96110 272781 96170 273670
rect 96107 272780 96173 272781
rect 96107 272716 96108 272780
rect 96172 272716 96173 272780
rect 96107 272715 96173 272716
rect 94451 272372 94517 272373
rect 94451 272308 94452 272372
rect 94516 272308 94517 272372
rect 94451 272307 94517 272308
rect 93347 270740 93413 270741
rect 93347 270676 93348 270740
rect 93412 270676 93413 270740
rect 93347 270675 93413 270676
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 252308 92414 255838
rect 95514 260114 96134 272000
rect 97030 271829 97090 273670
rect 97027 271828 97093 271829
rect 97027 271764 97028 271828
rect 97092 271764 97093 271828
rect 97027 271763 97093 271764
rect 98134 271693 98194 273670
rect 98502 272781 98562 273670
rect 99422 273670 99508 273730
rect 100672 273730 100732 274040
rect 101080 273730 101140 274040
rect 100672 273670 100770 273730
rect 98499 272780 98565 272781
rect 98499 272716 98500 272780
rect 98564 272716 98565 272780
rect 98499 272715 98565 272716
rect 99422 272237 99482 273670
rect 99419 272236 99485 272237
rect 99419 272172 99420 272236
rect 99484 272172 99485 272236
rect 99419 272171 99485 272172
rect 98131 271692 98197 271693
rect 98131 271628 98132 271692
rect 98196 271628 98197 271692
rect 98131 271627 98197 271628
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 252308 96134 259558
rect 99234 261954 99854 272000
rect 100710 271829 100770 273670
rect 101078 273670 101140 273730
rect 101760 273730 101820 274040
rect 102848 273730 102908 274040
rect 101760 273670 101874 273730
rect 100707 271828 100773 271829
rect 100707 271764 100708 271828
rect 100772 271764 100773 271828
rect 100707 271763 100773 271764
rect 101078 271557 101138 273670
rect 101814 273189 101874 273670
rect 102734 273670 102908 273730
rect 103528 273730 103588 274040
rect 103936 273730 103996 274040
rect 103528 273670 103714 273730
rect 101811 273188 101877 273189
rect 101811 273124 101812 273188
rect 101876 273124 101877 273188
rect 101811 273123 101877 273124
rect 102734 273053 102794 273670
rect 102731 273052 102797 273053
rect 102731 272988 102732 273052
rect 102796 272988 102797 273052
rect 102731 272987 102797 272988
rect 101075 271556 101141 271557
rect 101075 271492 101076 271556
rect 101140 271492 101141 271556
rect 101075 271491 101141 271492
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 252308 99854 261398
rect 102954 265674 103574 272000
rect 103654 271282 103714 273670
rect 103838 273670 103996 273730
rect 105296 273730 105356 274040
rect 105976 273730 106036 274040
rect 105296 273670 105370 273730
rect 103838 272917 103898 273670
rect 103835 272916 103901 272917
rect 103835 272852 103836 272916
rect 103900 272852 103901 272916
rect 103835 272851 103901 272852
rect 103835 271284 103901 271285
rect 103835 271282 103836 271284
rect 103654 271222 103836 271282
rect 103835 271220 103836 271222
rect 103900 271220 103901 271284
rect 103835 271219 103901 271220
rect 105310 270741 105370 273670
rect 105862 273670 106036 273730
rect 106384 273730 106444 274040
rect 107608 273730 107668 274040
rect 108288 273730 108348 274040
rect 108696 273730 108756 274040
rect 109784 273730 109844 274040
rect 106384 273670 106474 273730
rect 105862 271421 105922 273670
rect 106414 271829 106474 273670
rect 107518 273670 107668 273730
rect 108254 273670 108348 273730
rect 108622 273670 108756 273730
rect 109542 273670 109844 273730
rect 111008 273730 111068 274040
rect 111144 273730 111204 274040
rect 112232 273730 112292 274040
rect 113320 273869 113380 274040
rect 113317 273868 113383 273869
rect 113317 273804 113318 273868
rect 113382 273804 113383 273868
rect 113317 273803 113383 273804
rect 113592 273730 113652 274040
rect 114408 273730 114468 274040
rect 111008 273670 111074 273730
rect 111144 273670 111258 273730
rect 112232 273670 112362 273730
rect 107518 271829 107578 273670
rect 106411 271828 106477 271829
rect 106411 271764 106412 271828
rect 106476 271764 106477 271828
rect 106411 271763 106477 271764
rect 107515 271828 107581 271829
rect 107515 271764 107516 271828
rect 107580 271764 107581 271828
rect 107515 271763 107581 271764
rect 108254 271693 108314 273670
rect 108251 271692 108317 271693
rect 108251 271628 108252 271692
rect 108316 271628 108317 271692
rect 108251 271627 108317 271628
rect 105859 271420 105925 271421
rect 105859 271356 105860 271420
rect 105924 271356 105925 271420
rect 105859 271355 105925 271356
rect 105307 270740 105373 270741
rect 105307 270676 105308 270740
rect 105372 270676 105373 270740
rect 105307 270675 105373 270676
rect 108622 270605 108682 273670
rect 109542 271421 109602 273670
rect 109539 271420 109605 271421
rect 109539 271356 109540 271420
rect 109604 271356 109605 271420
rect 109539 271355 109605 271356
rect 108619 270604 108685 270605
rect 108619 270540 108620 270604
rect 108684 270540 108685 270604
rect 108619 270539 108685 270540
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 252308 103574 265118
rect 109794 255454 110414 272000
rect 111014 271285 111074 273670
rect 111011 271284 111077 271285
rect 111011 271220 111012 271284
rect 111076 271220 111077 271284
rect 111011 271219 111077 271220
rect 111198 270605 111258 273670
rect 112302 271829 112362 273670
rect 113222 273670 113652 273730
rect 114326 273670 114468 273730
rect 115768 273730 115828 274040
rect 116040 273730 116100 274040
rect 116992 273730 117052 274040
rect 118080 273730 118140 274040
rect 118488 273730 118548 274040
rect 119168 273730 119228 274040
rect 120936 273730 120996 274040
rect 115768 273670 115858 273730
rect 112299 271828 112365 271829
rect 112299 271764 112300 271828
rect 112364 271764 112365 271828
rect 112299 271763 112365 271764
rect 113222 271285 113282 273670
rect 113219 271284 113285 271285
rect 113219 271220 113220 271284
rect 113284 271220 113285 271284
rect 113219 271219 113285 271220
rect 111195 270604 111261 270605
rect 111195 270540 111196 270604
rect 111260 270540 111261 270604
rect 111195 270539 111261 270540
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 252308 110414 254898
rect 113514 259174 114134 272000
rect 114326 271421 114386 273670
rect 115798 271557 115858 273670
rect 115982 273670 116100 273730
rect 116902 273670 117052 273730
rect 118006 273670 118140 273730
rect 118374 273670 118548 273730
rect 119110 273670 119228 273730
rect 120766 273670 120996 273730
rect 123520 273730 123580 274040
rect 125968 273730 126028 274040
rect 123520 273670 123586 273730
rect 115982 271693 116042 273670
rect 116902 272645 116962 273670
rect 116899 272644 116965 272645
rect 116899 272580 116900 272644
rect 116964 272580 116965 272644
rect 116899 272579 116965 272580
rect 118006 272509 118066 273670
rect 118003 272508 118069 272509
rect 118003 272444 118004 272508
rect 118068 272444 118069 272508
rect 118003 272443 118069 272444
rect 115979 271692 116045 271693
rect 115979 271628 115980 271692
rect 116044 271628 116045 271692
rect 115979 271627 116045 271628
rect 115795 271556 115861 271557
rect 115795 271492 115796 271556
rect 115860 271492 115861 271556
rect 115795 271491 115861 271492
rect 114323 271420 114389 271421
rect 114323 271356 114324 271420
rect 114388 271356 114389 271420
rect 114323 271355 114389 271356
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 252308 114134 258618
rect 117234 262894 117854 272000
rect 118374 271693 118434 273670
rect 118371 271692 118437 271693
rect 118371 271628 118372 271692
rect 118436 271628 118437 271692
rect 118371 271627 118437 271628
rect 119110 271149 119170 273670
rect 120766 271693 120826 273670
rect 120763 271692 120829 271693
rect 120763 271628 120764 271692
rect 120828 271628 120829 271692
rect 120763 271627 120829 271628
rect 119107 271148 119173 271149
rect 119107 271084 119108 271148
rect 119172 271084 119173 271148
rect 119107 271083 119173 271084
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 252308 117854 262338
rect 120954 266614 121574 272000
rect 123526 271829 123586 273670
rect 125918 273670 126028 273730
rect 128280 273730 128340 274040
rect 131000 273730 131060 274040
rect 133448 273733 133508 274040
rect 128280 273670 128738 273730
rect 125918 271829 125978 273670
rect 123523 271828 123589 271829
rect 123523 271764 123524 271828
rect 123588 271764 123589 271828
rect 123523 271763 123589 271764
rect 125915 271828 125981 271829
rect 125915 271764 125916 271828
rect 125980 271764 125981 271828
rect 125915 271763 125981 271764
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 252308 121574 266058
rect 127794 256394 128414 272000
rect 128678 271829 128738 273670
rect 130886 273670 131060 273730
rect 133445 273732 133511 273733
rect 128675 271828 128741 271829
rect 128675 271764 128676 271828
rect 128740 271764 128741 271828
rect 128675 271763 128741 271764
rect 130886 271013 130946 273670
rect 133445 273668 133446 273732
rect 133510 273668 133511 273732
rect 133445 273667 133511 273668
rect 135896 273597 135956 274040
rect 138480 273597 138540 274040
rect 140928 273597 140988 274040
rect 143512 273597 143572 274040
rect 145960 273597 146020 274040
rect 148544 273730 148604 274040
rect 150992 273730 151052 274040
rect 148544 273670 148610 273730
rect 135893 273596 135959 273597
rect 135893 273532 135894 273596
rect 135958 273532 135959 273596
rect 135893 273531 135959 273532
rect 138477 273596 138543 273597
rect 138477 273532 138478 273596
rect 138542 273532 138543 273596
rect 138477 273531 138543 273532
rect 140925 273596 140991 273597
rect 140925 273532 140926 273596
rect 140990 273532 140991 273596
rect 140925 273531 140991 273532
rect 143509 273596 143575 273597
rect 143509 273532 143510 273596
rect 143574 273532 143575 273596
rect 143509 273531 143575 273532
rect 145957 273596 146023 273597
rect 145957 273532 145958 273596
rect 146022 273532 146023 273596
rect 145957 273531 146023 273532
rect 130883 271012 130949 271013
rect 130883 270948 130884 271012
rect 130948 270948 130949 271012
rect 130883 270947 130949 270948
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 252308 128414 255838
rect 131514 260114 132134 272000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 252308 132134 259558
rect 135234 261954 135854 272000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 252308 135854 261398
rect 138954 265674 139574 272000
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 252308 139574 265118
rect 145794 255454 146414 272000
rect 148550 270741 148610 273670
rect 150942 273670 151052 273730
rect 153440 273730 153500 274040
rect 155888 273730 155948 274040
rect 158472 273730 158532 274040
rect 160920 273730 160980 274040
rect 153440 273670 154130 273730
rect 155888 273670 155970 273730
rect 158472 273670 158546 273730
rect 148547 270740 148613 270741
rect 148547 270676 148548 270740
rect 148612 270676 148613 270740
rect 148547 270675 148613 270676
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 252308 146414 254898
rect 149514 259174 150134 272000
rect 150942 271829 151002 273670
rect 150939 271828 151005 271829
rect 150939 271764 150940 271828
rect 151004 271764 151005 271828
rect 150939 271763 151005 271764
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 252308 150134 258618
rect 153234 262894 153854 272000
rect 154070 271829 154130 273670
rect 155910 271829 155970 273670
rect 154067 271828 154133 271829
rect 154067 271764 154068 271828
rect 154132 271764 154133 271828
rect 154067 271763 154133 271764
rect 155907 271828 155973 271829
rect 155907 271764 155908 271828
rect 155972 271764 155973 271828
rect 155907 271763 155973 271764
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 252308 153854 262338
rect 156954 266614 157574 272000
rect 158486 271693 158546 273670
rect 160878 273670 160980 273730
rect 163368 273730 163428 274040
rect 165952 273730 166012 274040
rect 183224 273730 183284 274040
rect 163368 273670 163514 273730
rect 165952 273670 166090 273730
rect 160878 271693 160938 273670
rect 163454 271693 163514 273670
rect 158483 271692 158549 271693
rect 158483 271628 158484 271692
rect 158548 271628 158549 271692
rect 158483 271627 158549 271628
rect 160875 271692 160941 271693
rect 160875 271628 160876 271692
rect 160940 271628 160941 271692
rect 160875 271627 160941 271628
rect 163451 271692 163517 271693
rect 163451 271628 163452 271692
rect 163516 271628 163517 271692
rect 163451 271627 163517 271628
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 252308 157574 266058
rect 163794 256394 164414 272000
rect 166030 271693 166090 273670
rect 183142 273670 183284 273730
rect 183360 273730 183420 274040
rect 183360 273670 183570 273730
rect 166027 271692 166093 271693
rect 166027 271628 166028 271692
rect 166092 271628 166093 271692
rect 166027 271627 166093 271628
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 252308 164414 255838
rect 167514 260114 168134 272000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 252308 168134 259558
rect 171234 261954 171854 272000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 252308 171854 261398
rect 174954 265674 175574 272000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 252308 175574 265118
rect 181794 255454 182414 272000
rect 183142 271421 183202 273670
rect 183139 271420 183205 271421
rect 183139 271356 183140 271420
rect 183204 271356 183205 271420
rect 183139 271355 183205 271356
rect 183510 271149 183570 273670
rect 183507 271148 183573 271149
rect 183507 271084 183508 271148
rect 183572 271084 183573 271148
rect 183507 271083 183573 271084
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 178539 253196 178605 253197
rect 178539 253132 178540 253196
rect 178604 253132 178605 253196
rect 178539 253131 178605 253132
rect 179643 253196 179709 253197
rect 179643 253132 179644 253196
rect 179708 253132 179709 253196
rect 179643 253131 179709 253132
rect 59862 251910 60290 251970
rect 59862 166290 59922 251910
rect 178542 250610 178602 253131
rect 178464 250550 178602 250610
rect 179646 250610 179706 253131
rect 181794 252308 182414 254898
rect 185514 259174 186134 272000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 252308 186134 258618
rect 189234 262894 189854 272000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252308 189854 262338
rect 192954 266614 193574 272000
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 190867 253740 190933 253741
rect 190867 253676 190868 253740
rect 190932 253676 190933 253740
rect 190867 253675 190933 253676
rect 190870 250610 190930 253675
rect 192954 252308 193574 266058
rect 179646 250550 179748 250610
rect 178464 250240 178524 250550
rect 179688 250240 179748 250550
rect 190840 250550 190930 250610
rect 190840 250240 190900 250550
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 166290 76116 167106
rect 59862 166230 60290 166290
rect 59514 152114 60134 165000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 60230 145210 60290 166230
rect 76054 166230 76116 166290
rect 77144 166290 77204 167106
rect 78232 166290 78292 167106
rect 79592 166290 79652 167106
rect 80544 167010 80604 167106
rect 81768 167010 81828 167106
rect 83128 167010 83188 167106
rect 84216 167010 84276 167106
rect 85440 167010 85500 167106
rect 77144 166230 77218 166290
rect 78232 166230 78322 166290
rect 63234 155834 63854 165000
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 63854 155834
rect 63234 155514 63854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 63854 155514
rect 63234 145308 63854 155278
rect 66954 157674 67574 165000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 165000
rect 76054 164253 76114 166230
rect 77158 164389 77218 166230
rect 77155 164388 77221 164389
rect 77155 164324 77156 164388
rect 77220 164324 77221 164388
rect 77155 164323 77221 164324
rect 76051 164252 76117 164253
rect 76051 164188 76052 164252
rect 76116 164188 76117 164252
rect 76051 164187 76117 164188
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 165000
rect 78262 164253 78322 166230
rect 79550 166230 79652 166290
rect 80470 166950 80604 167010
rect 81758 166950 81828 167010
rect 83046 166950 83188 167010
rect 84150 166950 84276 167010
rect 85438 166950 85500 167010
rect 86528 167010 86588 167106
rect 87616 167010 87676 167106
rect 88296 167010 88356 167106
rect 88704 167010 88764 167106
rect 90064 167010 90124 167106
rect 86528 166950 86602 167010
rect 87616 166950 87706 167010
rect 88296 166950 88442 167010
rect 88704 166950 88810 167010
rect 79550 164253 79610 166230
rect 80470 164253 80530 166950
rect 81758 165613 81818 166950
rect 81755 165612 81821 165613
rect 81755 165548 81756 165612
rect 81820 165548 81821 165612
rect 81755 165547 81821 165548
rect 78259 164252 78325 164253
rect 78259 164188 78260 164252
rect 78324 164188 78325 164252
rect 78259 164187 78325 164188
rect 79547 164252 79613 164253
rect 79547 164188 79548 164252
rect 79612 164188 79613 164252
rect 79547 164187 79613 164188
rect 80467 164252 80533 164253
rect 80467 164188 80468 164252
rect 80532 164188 80533 164252
rect 80467 164187 80533 164188
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 165000
rect 83046 164253 83106 166950
rect 84150 164253 84210 166950
rect 85438 165613 85498 166950
rect 85435 165612 85501 165613
rect 85435 165548 85436 165612
rect 85500 165548 85501 165612
rect 85435 165547 85501 165548
rect 83043 164252 83109 164253
rect 83043 164188 83044 164252
rect 83108 164188 83109 164252
rect 83043 164187 83109 164188
rect 84147 164252 84213 164253
rect 84147 164188 84148 164252
rect 84212 164188 84213 164252
rect 84147 164187 84213 164188
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 165000
rect 86542 164253 86602 166950
rect 87646 164253 87706 166950
rect 88382 164933 88442 166950
rect 88379 164932 88445 164933
rect 88379 164868 88380 164932
rect 88444 164868 88445 164932
rect 88379 164867 88445 164868
rect 88750 164253 88810 166950
rect 90038 166950 90124 167010
rect 90744 167010 90804 167106
rect 91288 167010 91348 167106
rect 92376 167010 92436 167106
rect 93464 167010 93524 167106
rect 90744 166950 90834 167010
rect 91288 166950 91386 167010
rect 92376 166950 92490 167010
rect 90038 164389 90098 166950
rect 90774 165613 90834 166950
rect 90771 165612 90837 165613
rect 90771 165548 90772 165612
rect 90836 165548 90837 165612
rect 90771 165547 90837 165548
rect 90035 164388 90101 164389
rect 90035 164324 90036 164388
rect 90100 164324 90101 164388
rect 90035 164323 90101 164324
rect 91326 164253 91386 166950
rect 92430 165613 92490 166950
rect 93350 166950 93524 167010
rect 93600 167010 93660 167106
rect 94552 167010 94612 167106
rect 95912 167010 95972 167106
rect 93600 166950 93778 167010
rect 92427 165612 92493 165613
rect 92427 165548 92428 165612
rect 92492 165548 92493 165612
rect 92427 165547 92493 165548
rect 86539 164252 86605 164253
rect 86539 164188 86540 164252
rect 86604 164188 86605 164252
rect 86539 164187 86605 164188
rect 87643 164252 87709 164253
rect 87643 164188 87644 164252
rect 87708 164188 87709 164252
rect 87643 164187 87709 164188
rect 88747 164252 88813 164253
rect 88747 164188 88748 164252
rect 88812 164188 88813 164252
rect 88747 164187 88813 164188
rect 91323 164252 91389 164253
rect 91323 164188 91324 164252
rect 91388 164188 91389 164252
rect 91323 164187 91389 164188
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 165000
rect 93350 164253 93410 166950
rect 93718 166837 93778 166950
rect 94454 166950 94612 167010
rect 95742 166950 95972 167010
rect 96048 167010 96108 167106
rect 97000 167010 97060 167106
rect 98088 167010 98148 167106
rect 98496 167010 98556 167106
rect 99448 167010 99508 167106
rect 96048 166950 96170 167010
rect 97000 166950 97090 167010
rect 98088 166950 98194 167010
rect 98496 166950 98562 167010
rect 93715 166836 93781 166837
rect 93715 166772 93716 166836
rect 93780 166772 93781 166836
rect 93715 166771 93781 166772
rect 94454 164253 94514 166950
rect 95742 165613 95802 166950
rect 96110 166293 96170 166950
rect 96107 166292 96173 166293
rect 96107 166228 96108 166292
rect 96172 166228 96173 166292
rect 96107 166227 96173 166228
rect 95739 165612 95805 165613
rect 95739 165548 95740 165612
rect 95804 165548 95805 165612
rect 95739 165547 95805 165548
rect 93347 164252 93413 164253
rect 93347 164188 93348 164252
rect 93412 164188 93413 164252
rect 93347 164187 93413 164188
rect 94451 164252 94517 164253
rect 94451 164188 94452 164252
rect 94516 164188 94517 164252
rect 94451 164187 94517 164188
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 165000
rect 97030 164253 97090 166950
rect 98134 164253 98194 166950
rect 98502 166837 98562 166950
rect 99422 166950 99508 167010
rect 100672 167010 100732 167106
rect 101080 167010 101140 167106
rect 100672 166950 100770 167010
rect 98499 166836 98565 166837
rect 98499 166772 98500 166836
rect 98564 166772 98565 166836
rect 98499 166771 98565 166772
rect 99422 165613 99482 166950
rect 99419 165612 99485 165613
rect 99419 165548 99420 165612
rect 99484 165548 99485 165612
rect 99419 165547 99485 165548
rect 97027 164252 97093 164253
rect 97027 164188 97028 164252
rect 97092 164188 97093 164252
rect 97027 164187 97093 164188
rect 98131 164252 98197 164253
rect 98131 164188 98132 164252
rect 98196 164188 98197 164252
rect 98131 164187 98197 164188
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 155834 99854 165000
rect 100710 164525 100770 166950
rect 101078 166950 101140 167010
rect 101760 167010 101820 167106
rect 102848 167010 102908 167106
rect 103528 167010 103588 167106
rect 103936 167010 103996 167106
rect 101760 166950 101874 167010
rect 101078 166837 101138 166950
rect 101075 166836 101141 166837
rect 101075 166772 101076 166836
rect 101140 166772 101141 166836
rect 101075 166771 101141 166772
rect 100707 164524 100773 164525
rect 100707 164460 100708 164524
rect 100772 164460 100773 164524
rect 100707 164459 100773 164460
rect 101814 164253 101874 166950
rect 102734 166950 102908 167010
rect 103470 166950 103588 167010
rect 103838 166950 103996 167010
rect 105296 167010 105356 167106
rect 105976 167010 106036 167106
rect 105296 166950 105370 167010
rect 102734 164253 102794 166950
rect 103470 165613 103530 166950
rect 103467 165612 103533 165613
rect 103467 165548 103468 165612
rect 103532 165548 103533 165612
rect 103467 165547 103533 165548
rect 101811 164252 101877 164253
rect 101811 164188 101812 164252
rect 101876 164188 101877 164252
rect 101811 164187 101877 164188
rect 102731 164252 102797 164253
rect 102731 164188 102732 164252
rect 102796 164188 102797 164252
rect 102731 164187 102797 164188
rect 99234 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 99854 155834
rect 99234 155514 99854 155598
rect 99234 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 99854 155514
rect 99234 145308 99854 155278
rect 102954 157674 103574 165000
rect 103838 164253 103898 166950
rect 105310 164253 105370 166950
rect 105862 166950 106036 167010
rect 106384 167010 106444 167106
rect 107608 167010 107668 167106
rect 108288 167010 108348 167106
rect 108696 167010 108756 167106
rect 106384 166950 106474 167010
rect 105862 166837 105922 166950
rect 105859 166836 105925 166837
rect 105859 166772 105860 166836
rect 105924 166772 105925 166836
rect 105859 166771 105925 166772
rect 106414 164253 106474 166950
rect 107518 166950 107668 167010
rect 108254 166950 108348 167010
rect 108622 166950 108756 167010
rect 107518 164797 107578 166950
rect 108254 166837 108314 166950
rect 108251 166836 108317 166837
rect 108251 166772 108252 166836
rect 108316 166772 108317 166836
rect 108251 166771 108317 166772
rect 108622 164933 108682 166950
rect 109784 166290 109844 167106
rect 109726 166230 109844 166290
rect 111008 166290 111068 167106
rect 111144 166290 111204 167106
rect 112232 166290 112292 167106
rect 113320 166290 113380 167106
rect 113592 166290 113652 167106
rect 114408 166565 114468 167106
rect 114405 166564 114471 166565
rect 114405 166500 114406 166564
rect 114470 166500 114471 166564
rect 114405 166499 114471 166500
rect 111008 166230 111074 166290
rect 111144 166230 111258 166290
rect 112232 166230 112362 166290
rect 109726 165613 109786 166230
rect 111014 165613 111074 166230
rect 111198 165613 111258 166230
rect 112302 165613 112362 166230
rect 113222 166230 113380 166290
rect 113590 166230 113652 166290
rect 115768 166290 115828 167106
rect 116040 166290 116100 167106
rect 116992 166565 117052 167106
rect 116989 166564 117055 166565
rect 116989 166500 116990 166564
rect 117054 166500 117055 166564
rect 116989 166499 117055 166500
rect 118080 166290 118140 167106
rect 118488 166290 118548 167106
rect 119168 166290 119228 167106
rect 115768 166230 115858 166290
rect 109723 165612 109789 165613
rect 109723 165548 109724 165612
rect 109788 165548 109789 165612
rect 109723 165547 109789 165548
rect 111011 165612 111077 165613
rect 111011 165548 111012 165612
rect 111076 165548 111077 165612
rect 111011 165547 111077 165548
rect 111195 165612 111261 165613
rect 111195 165548 111196 165612
rect 111260 165548 111261 165612
rect 111195 165547 111261 165548
rect 112299 165612 112365 165613
rect 112299 165548 112300 165612
rect 112364 165548 112365 165612
rect 112299 165547 112365 165548
rect 108619 164932 108685 164933
rect 108619 164868 108620 164932
rect 108684 164868 108685 164932
rect 108619 164867 108685 164868
rect 107515 164796 107581 164797
rect 107515 164732 107516 164796
rect 107580 164732 107581 164796
rect 107515 164731 107581 164732
rect 103835 164252 103901 164253
rect 103835 164188 103836 164252
rect 103900 164188 103901 164252
rect 103835 164187 103901 164188
rect 105307 164252 105373 164253
rect 105307 164188 105308 164252
rect 105372 164188 105373 164252
rect 105307 164187 105373 164188
rect 106411 164252 106477 164253
rect 106411 164188 106412 164252
rect 106476 164188 106477 164252
rect 106411 164187 106477 164188
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 165000
rect 113222 164525 113282 166230
rect 113590 165613 113650 166230
rect 113587 165612 113653 165613
rect 113587 165548 113588 165612
rect 113652 165548 113653 165612
rect 113587 165547 113653 165548
rect 113219 164524 113285 164525
rect 113219 164460 113220 164524
rect 113284 164460 113285 164524
rect 113219 164459 113285 164460
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 165000
rect 115798 164525 115858 166230
rect 115982 166230 116100 166290
rect 118006 166230 118140 166290
rect 118374 166230 118548 166290
rect 119110 166230 119228 166290
rect 120936 166290 120996 167106
rect 123520 166290 123580 167106
rect 125968 166290 126028 167106
rect 128280 167010 128340 167106
rect 131000 167010 131060 167106
rect 128280 166950 128554 167010
rect 128280 166910 128370 166950
rect 120936 166230 121010 166290
rect 123520 166230 123586 166290
rect 115982 165613 116042 166230
rect 118006 165613 118066 166230
rect 118374 165613 118434 166230
rect 119110 165613 119170 166230
rect 120950 165613 121010 166230
rect 123526 165613 123586 166230
rect 125918 166230 126028 166290
rect 125918 165613 125978 166230
rect 128494 165613 128554 166950
rect 130886 166950 131060 167010
rect 133448 167010 133508 167106
rect 135896 167010 135956 167106
rect 133448 166950 133522 167010
rect 135896 166950 136098 167010
rect 130886 165613 130946 166950
rect 133462 165613 133522 166950
rect 115979 165612 116045 165613
rect 115979 165548 115980 165612
rect 116044 165548 116045 165612
rect 115979 165547 116045 165548
rect 118003 165612 118069 165613
rect 118003 165548 118004 165612
rect 118068 165548 118069 165612
rect 118003 165547 118069 165548
rect 118371 165612 118437 165613
rect 118371 165548 118372 165612
rect 118436 165548 118437 165612
rect 118371 165547 118437 165548
rect 119107 165612 119173 165613
rect 119107 165548 119108 165612
rect 119172 165548 119173 165612
rect 119107 165547 119173 165548
rect 120947 165612 121013 165613
rect 120947 165548 120948 165612
rect 121012 165548 121013 165612
rect 120947 165547 121013 165548
rect 123523 165612 123589 165613
rect 123523 165548 123524 165612
rect 123588 165548 123589 165612
rect 123523 165547 123589 165548
rect 125915 165612 125981 165613
rect 125915 165548 125916 165612
rect 125980 165548 125981 165612
rect 125915 165547 125981 165548
rect 128491 165612 128557 165613
rect 128491 165548 128492 165612
rect 128556 165548 128557 165612
rect 128491 165547 128557 165548
rect 130883 165612 130949 165613
rect 130883 165548 130884 165612
rect 130948 165548 130949 165612
rect 130883 165547 130949 165548
rect 133459 165612 133525 165613
rect 133459 165548 133460 165612
rect 133524 165548 133525 165612
rect 133459 165547 133525 165548
rect 136038 165069 136098 166950
rect 138480 166837 138540 167106
rect 140928 166837 140988 167106
rect 143512 166837 143572 167106
rect 145960 166837 146020 167106
rect 148544 167010 148604 167106
rect 150992 167010 151052 167106
rect 153440 167010 153500 167106
rect 148544 166950 148610 167010
rect 138477 166836 138543 166837
rect 138477 166772 138478 166836
rect 138542 166772 138543 166836
rect 138477 166771 138543 166772
rect 140925 166836 140991 166837
rect 140925 166772 140926 166836
rect 140990 166772 140991 166836
rect 140925 166771 140991 166772
rect 143509 166836 143575 166837
rect 143509 166772 143510 166836
rect 143574 166772 143575 166836
rect 143509 166771 143575 166772
rect 145957 166836 146023 166837
rect 145957 166772 145958 166836
rect 146022 166772 146023 166836
rect 145957 166771 146023 166772
rect 148550 166565 148610 166950
rect 150942 166950 151052 167010
rect 153334 166950 153500 167010
rect 155888 167010 155948 167106
rect 155888 166950 155970 167010
rect 148547 166564 148613 166565
rect 148547 166500 148548 166564
rect 148612 166500 148613 166564
rect 148547 166499 148613 166500
rect 150942 165205 151002 166950
rect 153334 166565 153394 166950
rect 153331 166564 153397 166565
rect 153331 166500 153332 166564
rect 153396 166500 153397 166564
rect 153331 166499 153397 166500
rect 155910 165341 155970 166950
rect 158472 166290 158532 167106
rect 160920 166290 160980 167106
rect 163368 166701 163428 167106
rect 165952 166701 166012 167106
rect 163365 166700 163431 166701
rect 163365 166636 163366 166700
rect 163430 166636 163431 166700
rect 163365 166635 163431 166636
rect 165949 166700 166015 166701
rect 165949 166636 165950 166700
rect 166014 166636 166015 166700
rect 165949 166635 166015 166636
rect 183224 166565 183284 167106
rect 183221 166564 183287 166565
rect 183221 166500 183222 166564
rect 183286 166500 183287 166564
rect 183221 166499 183287 166500
rect 183360 166290 183420 167106
rect 196574 166429 196634 485419
rect 197859 485348 197925 485349
rect 197859 485284 197860 485348
rect 197924 485284 197925 485348
rect 197859 485283 197925 485284
rect 196755 484940 196821 484941
rect 196755 484876 196756 484940
rect 196820 484876 196821 484940
rect 196755 484875 196821 484876
rect 196758 273053 196818 484875
rect 196755 273052 196821 273053
rect 196755 272988 196756 273052
rect 196820 272988 196821 273052
rect 196755 272987 196821 272988
rect 196571 166428 196637 166429
rect 196571 166364 196572 166428
rect 196636 166364 196637 166428
rect 196571 166363 196637 166364
rect 158472 166230 158546 166290
rect 158486 165477 158546 166230
rect 160878 166230 160980 166290
rect 183326 166230 183420 166290
rect 158483 165476 158549 165477
rect 158483 165412 158484 165476
rect 158548 165412 158549 165476
rect 158483 165411 158549 165412
rect 155907 165340 155973 165341
rect 155907 165276 155908 165340
rect 155972 165276 155973 165340
rect 155907 165275 155973 165276
rect 150939 165204 151005 165205
rect 150939 165140 150940 165204
rect 151004 165140 151005 165204
rect 150939 165139 151005 165140
rect 136035 165068 136101 165069
rect 136035 165004 136036 165068
rect 136100 165004 136101 165068
rect 136035 165003 136101 165004
rect 115795 164524 115861 164525
rect 115795 164460 115796 164524
rect 115860 164460 115861 164524
rect 115795 164459 115861 164460
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 165000
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 165000
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 165000
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 165000
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 155834 135854 165000
rect 135234 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 135854 155834
rect 135234 155514 135854 155598
rect 135234 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 135854 155514
rect 135234 145308 135854 155278
rect 138954 157674 139574 165000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 165000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 165000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 165000
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 165000
rect 160878 164661 160938 166230
rect 183326 165613 183386 166230
rect 183323 165612 183389 165613
rect 183323 165548 183324 165612
rect 183388 165548 183389 165612
rect 183323 165547 183389 165548
rect 160875 164660 160941 164661
rect 160875 164596 160876 164660
rect 160940 164596 160941 164660
rect 160875 164595 160941 164596
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 165000
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 165000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 155834 171854 165000
rect 171234 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 171854 155834
rect 171234 155514 171854 155598
rect 171234 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 171854 155514
rect 171234 145308 171854 155278
rect 174954 157674 175574 165000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 165000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 165000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 165000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 165000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 145308 193574 158058
rect 59862 145150 60290 145210
rect 59862 59530 59922 145150
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 190867 144940 190933 144941
rect 190867 144876 190868 144940
rect 190932 144876 190933 144940
rect 190867 144875 190933 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 144875
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 59862 59470 60290 59530
rect 59307 58716 59373 58717
rect 59307 58652 59308 58716
rect 59372 58652 59373 58716
rect 59307 58651 59373 58652
rect 59123 58444 59189 58445
rect 59123 58380 59124 58444
rect 59188 58380 59189 58444
rect 59123 58379 59189 58380
rect 58939 57220 59005 57221
rect 58939 57156 58940 57220
rect 59004 57156 59005 57220
rect 58939 57155 59005 57156
rect 58755 57084 58821 57085
rect 58755 57020 58756 57084
rect 58820 57020 58821 57084
rect 58755 57019 58821 57020
rect 57467 56132 57533 56133
rect 57467 56068 57468 56132
rect 57532 56068 57533 56132
rect 57467 56067 57533 56068
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 60230 57765 60290 59470
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59530 80604 60106
rect 78232 59470 78322 59530
rect 60227 57764 60293 57765
rect 60227 57700 60228 57764
rect 60292 57700 60293 57764
rect 60227 57699 60293 57700
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59470 80604 59530
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84216 59530 84276 60106
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 79550 57901 79610 59470
rect 80470 57901 80530 59470
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 83966 59470 84276 59530
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59533 90124 60106
rect 90035 59532 90124 59533
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 83966 58037 84026 59470
rect 85438 58173 85498 59470
rect 85435 58172 85501 58173
rect 85435 58108 85436 58172
rect 85500 58108 85501 58172
rect 85435 58107 85501 58108
rect 83963 58036 84029 58037
rect 83963 57972 83964 58036
rect 84028 57972 84029 58036
rect 83963 57971 84029 57972
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 88382 57901 88442 59470
rect 88750 57901 88810 59470
rect 90035 59468 90036 59532
rect 90100 59470 90124 59532
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 92376 59470 92490 59530
rect 90100 59468 90101 59470
rect 90035 59467 90101 59468
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92430 58173 92490 59470
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59805 94612 60106
rect 94549 59804 94615 59805
rect 94549 59740 94550 59804
rect 94614 59740 94615 59804
rect 94549 59739 94615 59740
rect 95912 59533 95972 60106
rect 96048 59666 96108 60106
rect 96048 59606 96354 59666
rect 95912 59532 95989 59533
rect 93600 59470 93778 59530
rect 95912 59470 95924 59532
rect 92427 58172 92493 58173
rect 92427 58108 92428 58172
rect 92492 58108 92493 58172
rect 92427 58107 92493 58108
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88379 57900 88445 57901
rect 88379 57836 88380 57900
rect 88444 57836 88445 57900
rect 88379 57835 88445 57836
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93718 57901 93778 59470
rect 95923 59468 95924 59470
rect 95988 59468 95989 59532
rect 95923 59467 95989 59468
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 93715 57900 93781 57901
rect 93715 57836 93716 57900
rect 93780 57836 93781 57900
rect 93715 57835 93781 57836
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 57085 96354 59606
rect 97000 59533 97060 60106
rect 98088 59533 98148 60106
rect 97000 59532 97093 59533
rect 97000 59470 97028 59532
rect 97027 59468 97028 59470
rect 97092 59468 97093 59532
rect 98088 59532 98197 59533
rect 98088 59470 98132 59532
rect 97027 59467 97093 59468
rect 98131 59468 98132 59470
rect 98196 59468 98197 59532
rect 98496 59530 98556 60106
rect 99448 59530 99508 60106
rect 100672 59666 100732 60106
rect 100672 59606 100770 59666
rect 100710 59533 100770 59606
rect 98496 59470 98562 59530
rect 98131 59467 98197 59468
rect 98502 57221 98562 59470
rect 99422 59470 99508 59530
rect 100707 59532 100773 59533
rect 99422 58173 99482 59470
rect 100707 59468 100708 59532
rect 100772 59468 100773 59532
rect 101080 59530 101140 60106
rect 101760 59805 101820 60106
rect 102848 59805 102908 60106
rect 101757 59804 101823 59805
rect 101757 59740 101758 59804
rect 101822 59740 101823 59804
rect 101757 59739 101823 59740
rect 102845 59804 102911 59805
rect 102845 59740 102846 59804
rect 102910 59740 102911 59804
rect 102845 59739 102911 59740
rect 100707 59467 100773 59468
rect 101078 59470 101140 59530
rect 103528 59530 103588 60106
rect 103936 59530 103996 60106
rect 105296 59669 105356 60106
rect 105976 59669 106036 60106
rect 105293 59668 105359 59669
rect 105293 59604 105294 59668
rect 105358 59604 105359 59668
rect 105293 59603 105359 59604
rect 105973 59668 106039 59669
rect 105973 59604 105974 59668
rect 106038 59604 106039 59668
rect 105973 59603 106039 59604
rect 103528 59470 103714 59530
rect 101078 58445 101138 59470
rect 101075 58444 101141 58445
rect 101075 58380 101076 58444
rect 101140 58380 101141 58444
rect 101075 58379 101141 58380
rect 99419 58172 99485 58173
rect 99419 58108 99420 58172
rect 99484 58108 99485 58172
rect 99419 58107 99485 58108
rect 98499 57220 98565 57221
rect 98499 57156 98500 57220
rect 98564 57156 98565 57220
rect 98499 57155 98565 57156
rect 96291 57084 96357 57085
rect 96291 57020 96292 57084
rect 96356 57020 96357 57084
rect 96291 57019 96357 57020
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103654 57218 103714 59470
rect 103838 59470 103996 59530
rect 106384 59530 106444 60106
rect 107608 59669 107668 60106
rect 107605 59668 107671 59669
rect 107605 59604 107606 59668
rect 107670 59604 107671 59668
rect 107605 59603 107671 59604
rect 108288 59530 108348 60106
rect 108696 59530 108756 60106
rect 109784 59530 109844 60106
rect 106384 59470 106474 59530
rect 103838 57901 103898 59470
rect 106414 57901 106474 59470
rect 108254 59470 108348 59530
rect 108622 59470 108756 59530
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59530 112292 60106
rect 113320 59530 113380 60106
rect 113592 59805 113652 60106
rect 113589 59804 113655 59805
rect 113589 59740 113590 59804
rect 113654 59740 113655 59804
rect 113589 59739 113655 59740
rect 114408 59530 114468 60106
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 108254 58581 108314 59470
rect 108251 58580 108317 58581
rect 108251 58516 108252 58580
rect 108316 58516 108317 58580
rect 108251 58515 108317 58516
rect 108622 57901 108682 59470
rect 109542 57901 109602 59470
rect 111014 59397 111074 59470
rect 111011 59396 111077 59397
rect 111011 59332 111012 59396
rect 111076 59332 111077 59396
rect 111011 59331 111077 59332
rect 103835 57900 103901 57901
rect 103835 57836 103836 57900
rect 103900 57836 103901 57900
rect 103835 57835 103901 57836
rect 106411 57900 106477 57901
rect 106411 57836 106412 57900
rect 106476 57836 106477 57900
rect 106411 57835 106477 57836
rect 108619 57900 108685 57901
rect 108619 57836 108620 57900
rect 108684 57836 108685 57900
rect 108619 57835 108685 57836
rect 109539 57900 109605 57901
rect 109539 57836 109540 57900
rect 109604 57836 109605 57900
rect 109539 57835 109605 57836
rect 103835 57220 103901 57221
rect 103835 57218 103836 57220
rect 103654 57158 103836 57218
rect 103835 57156 103836 57158
rect 103900 57156 103901 57220
rect 103835 57155 103901 57156
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 111198 57901 111258 59470
rect 112118 59470 112292 59530
rect 113222 59470 113380 59530
rect 114326 59470 114468 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59530 117052 60106
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 115768 59470 115858 59530
rect 112118 57901 112178 59470
rect 113222 58173 113282 59470
rect 113219 58172 113285 58173
rect 113219 58108 113220 58172
rect 113284 58108 113285 58172
rect 113219 58107 113285 58108
rect 113038 57930 113282 57990
rect 111195 57900 111261 57901
rect 111195 57836 111196 57900
rect 111260 57836 111261 57900
rect 111195 57835 111261 57836
rect 112115 57900 112181 57901
rect 112115 57836 112116 57900
rect 112180 57836 112181 57900
rect 112115 57835 112181 57836
rect 113038 57357 113098 57930
rect 113035 57356 113101 57357
rect 113035 57292 113036 57356
rect 113100 57292 113101 57356
rect 113035 57291 113101 57292
rect 113222 57221 113282 57930
rect 113219 57220 113285 57221
rect 113219 57156 113220 57220
rect 113284 57156 113285 57220
rect 113219 57155 113285 57156
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 114326 57221 114386 59470
rect 115798 57901 115858 59470
rect 115982 59470 116100 59530
rect 116902 59470 117052 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 120936 59530 120996 60106
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 120936 59470 121010 59530
rect 123520 59470 123586 59530
rect 115982 57901 116042 59470
rect 115795 57900 115861 57901
rect 115795 57836 115796 57900
rect 115860 57836 115861 57900
rect 115795 57835 115861 57836
rect 115979 57900 116045 57901
rect 115979 57836 115980 57900
rect 116044 57836 116045 57900
rect 115979 57835 116045 57836
rect 116902 57629 116962 59470
rect 116899 57628 116965 57629
rect 116899 57564 116900 57628
rect 116964 57564 116965 57628
rect 116899 57563 116965 57564
rect 114323 57220 114389 57221
rect 114323 57156 114324 57220
rect 114388 57156 114389 57220
rect 114323 57155 114389 57156
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57493 118066 59470
rect 118003 57492 118069 57493
rect 118003 57428 118004 57492
rect 118068 57428 118069 57492
rect 118003 57427 118069 57428
rect 118374 57357 118434 59470
rect 119110 57901 119170 59470
rect 120950 58717 121010 59470
rect 120947 58716 121013 58717
rect 120947 58652 120948 58716
rect 121012 58652 121013 58716
rect 120947 58651 121013 58652
rect 119107 57900 119173 57901
rect 119107 57836 119108 57900
rect 119172 57836 119173 57900
rect 119107 57835 119173 57836
rect 118371 57356 118437 57357
rect 118371 57292 118372 57356
rect 118436 57292 118437 57356
rect 118371 57291 118437 57292
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57629 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128738 59530
rect 125918 57765 125978 59470
rect 125915 57764 125981 57765
rect 125915 57700 125916 57764
rect 125980 57700 125981 57764
rect 125915 57699 125981 57700
rect 123523 57628 123589 57629
rect 123523 57564 123524 57628
rect 123588 57564 123589 57628
rect 123523 57563 123589 57564
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 128678 56677 128738 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 133448 59470 133522 59530
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 128675 56676 128741 56677
rect 128675 56612 128676 56676
rect 128740 56612 128741 56676
rect 128675 56611 128741 56612
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 57901 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 143512 59530 143572 60106
rect 145960 59530 146020 60106
rect 143512 59470 143642 59530
rect 135854 58853 135914 59470
rect 138430 58989 138490 59470
rect 140822 59125 140882 59470
rect 143582 59261 143642 59470
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 143579 59260 143645 59261
rect 143579 59196 143580 59260
rect 143644 59196 143645 59260
rect 143579 59195 143645 59196
rect 140819 59124 140885 59125
rect 140819 59060 140820 59124
rect 140884 59060 140885 59124
rect 140819 59059 140885 59060
rect 138427 58988 138493 58989
rect 138427 58924 138428 58988
rect 138492 58924 138493 58988
rect 138427 58923 138493 58924
rect 135851 58852 135917 58853
rect 135851 58788 135852 58852
rect 135916 58788 135917 58852
rect 135851 58787 135917 58788
rect 133459 57900 133525 57901
rect 133459 57836 133460 57900
rect 133524 57836 133525 57900
rect 133459 57835 133525 57836
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 56677 155970 59470
rect 155907 56676 155973 56677
rect 155907 56612 155908 56676
rect 155972 56612 155973 56676
rect 155907 56611 155973 56612
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 56677 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 160878 57629 160938 59470
rect 163270 57629 163330 59470
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163267 57628 163333 57629
rect 163267 57564 163268 57628
rect 163332 57564 163333 57628
rect 163267 57563 163333 57564
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 158483 56676 158549 56677
rect 158483 56612 158484 56676
rect 158548 56612 158549 56676
rect 158483 56611 158549 56612
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57765 183202 59470
rect 183510 57901 183570 59470
rect 197862 58717 197922 485283
rect 198046 166973 198106 485555
rect 198411 484940 198477 484941
rect 198411 484876 198412 484940
rect 198476 484876 198477 484940
rect 198411 484875 198477 484876
rect 198043 166972 198109 166973
rect 198043 166908 198044 166972
rect 198108 166908 198109 166972
rect 198043 166907 198109 166908
rect 198414 59261 198474 484875
rect 198595 484804 198661 484805
rect 198595 484740 198596 484804
rect 198660 484740 198661 484804
rect 198595 484739 198661 484740
rect 198411 59260 198477 59261
rect 198411 59196 198412 59260
rect 198476 59196 198477 59260
rect 198411 59195 198477 59196
rect 197859 58716 197925 58717
rect 197859 58652 197860 58716
rect 197924 58652 197925 58716
rect 197859 58651 197925 58652
rect 183507 57900 183573 57901
rect 183507 57836 183508 57900
rect 183572 57836 183573 57900
rect 183507 57835 183573 57836
rect 183139 57764 183205 57765
rect 183139 57700 183140 57764
rect 183204 57700 183205 57764
rect 183139 57699 183205 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 198598 56405 198658 484739
rect 198779 466172 198845 466173
rect 198779 466108 198780 466172
rect 198844 466108 198845 466172
rect 198779 466107 198845 466108
rect 198782 271693 198842 466107
rect 199147 464404 199213 464405
rect 199147 464340 199148 464404
rect 199212 464340 199213 464404
rect 199147 464339 199213 464340
rect 199150 381581 199210 464339
rect 199147 381580 199213 381581
rect 199147 381516 199148 381580
rect 199212 381516 199213 381580
rect 199147 381515 199213 381516
rect 199334 273189 199394 485691
rect 199794 472394 200414 486000
rect 201355 485348 201421 485349
rect 201355 485284 201356 485348
rect 201420 485284 201421 485348
rect 201355 485283 201421 485284
rect 200803 485212 200869 485213
rect 200803 485148 200804 485212
rect 200868 485148 200869 485212
rect 200803 485147 200869 485148
rect 200619 485076 200685 485077
rect 200619 485012 200620 485076
rect 200684 485012 200685 485076
rect 200619 485011 200685 485012
rect 199794 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 200414 472394
rect 199794 472074 200414 472158
rect 199794 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 200414 472074
rect 199515 471748 199581 471749
rect 199515 471684 199516 471748
rect 199580 471684 199581 471748
rect 199515 471683 199581 471684
rect 199518 273325 199578 471683
rect 199794 453454 200414 471838
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199515 273324 199581 273325
rect 199515 273260 199516 273324
rect 199580 273260 199581 273324
rect 199515 273259 199581 273260
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199331 273188 199397 273189
rect 199331 273124 199332 273188
rect 199396 273124 199397 273188
rect 199331 273123 199397 273124
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 198779 271692 198845 271693
rect 198779 271628 198780 271692
rect 198844 271628 198845 271692
rect 198779 271627 198845 271628
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 200622 58581 200682 485011
rect 200806 59397 200866 485147
rect 200987 468756 201053 468757
rect 200987 468692 200988 468756
rect 201052 468692 201053 468756
rect 200987 468691 201053 468692
rect 200990 164797 201050 468691
rect 200987 164796 201053 164797
rect 200987 164732 200988 164796
rect 201052 164732 201053 164796
rect 200987 164731 201053 164732
rect 200803 59396 200869 59397
rect 200803 59332 200804 59396
rect 200868 59332 200869 59396
rect 200803 59331 200869 59332
rect 201358 58989 201418 485283
rect 202643 485212 202709 485213
rect 202643 485148 202644 485212
rect 202708 485148 202709 485212
rect 202643 485147 202709 485148
rect 202459 480996 202525 480997
rect 202459 480932 202460 480996
rect 202524 480932 202525 480996
rect 202459 480931 202525 480932
rect 202091 475420 202157 475421
rect 202091 475356 202092 475420
rect 202156 475356 202157 475420
rect 202091 475355 202157 475356
rect 201355 58988 201421 58989
rect 201355 58924 201356 58988
rect 201420 58924 201421 58988
rect 201355 58923 201421 58924
rect 200619 58580 200685 58581
rect 200619 58516 200620 58580
rect 200684 58516 200685 58580
rect 200619 58515 200685 58516
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 198595 56404 198661 56405
rect 198595 56340 198596 56404
rect 198660 56340 198661 56404
rect 198595 56339 198661 56340
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 202094 3909 202154 475355
rect 202275 472700 202341 472701
rect 202275 472636 202276 472700
rect 202340 472636 202341 472700
rect 202275 472635 202341 472636
rect 202278 57629 202338 472635
rect 202462 164389 202522 480931
rect 202646 380765 202706 485147
rect 203514 476114 204134 486000
rect 205219 485212 205285 485213
rect 205219 485148 205220 485212
rect 205284 485148 205285 485212
rect 205219 485147 205285 485148
rect 203514 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 204134 476114
rect 203514 475794 204134 475878
rect 203514 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 204134 475794
rect 203195 472564 203261 472565
rect 203195 472500 203196 472564
rect 203260 472500 203261 472564
rect 203195 472499 203261 472500
rect 202643 380764 202709 380765
rect 202643 380700 202644 380764
rect 202708 380700 202709 380764
rect 202643 380699 202709 380700
rect 202459 164388 202525 164389
rect 202459 164324 202460 164388
rect 202524 164324 202525 164388
rect 202459 164323 202525 164324
rect 202275 57628 202341 57629
rect 202275 57564 202276 57628
rect 202340 57564 202341 57628
rect 202275 57563 202341 57564
rect 203198 57357 203258 472499
rect 203514 457174 204134 475558
rect 204851 471612 204917 471613
rect 204851 471548 204852 471612
rect 204916 471548 204917 471612
rect 204851 471547 204917 471548
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 368114 204134 384618
rect 203514 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 204134 368114
rect 203514 367794 204134 367878
rect 203514 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 204134 367794
rect 203514 349174 204134 367558
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 152114 204134 168618
rect 204854 165341 204914 471547
rect 205035 468892 205101 468893
rect 205035 468828 205036 468892
rect 205100 468828 205101 468892
rect 205035 468827 205101 468828
rect 205038 166837 205098 468827
rect 205222 380765 205282 485147
rect 205403 484940 205469 484941
rect 205403 484876 205404 484940
rect 205468 484876 205469 484940
rect 205403 484875 205469 484876
rect 205219 380764 205285 380765
rect 205219 380700 205220 380764
rect 205284 380700 205285 380764
rect 205219 380699 205285 380700
rect 205406 378453 205466 484875
rect 205403 378452 205469 378453
rect 205403 378388 205404 378452
rect 205468 378388 205469 378452
rect 205403 378387 205469 378388
rect 205035 166836 205101 166837
rect 205035 166772 205036 166836
rect 205100 166772 205101 166836
rect 205035 166771 205101 166772
rect 204851 165340 204917 165341
rect 204851 165276 204852 165340
rect 204916 165276 204917 165340
rect 204851 165275 204917 165276
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203195 57356 203261 57357
rect 203195 57292 203196 57356
rect 203260 57292 203261 57356
rect 203195 57291 203261 57292
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 202091 3908 202157 3909
rect 202091 3844 202092 3908
rect 202156 3844 202157 3908
rect 202091 3843 202157 3844
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 24618
rect 206142 3229 206202 486371
rect 206691 484804 206757 484805
rect 206691 484740 206692 484804
rect 206756 484740 206757 484804
rect 206691 484739 206757 484740
rect 206323 469028 206389 469029
rect 206323 468964 206324 469028
rect 206388 468964 206389 469028
rect 206323 468963 206389 468964
rect 206326 164117 206386 468963
rect 206507 468620 206573 468621
rect 206507 468556 206508 468620
rect 206572 468556 206573 468620
rect 206507 468555 206573 468556
rect 206510 164933 206570 468555
rect 206694 415309 206754 484739
rect 207234 477954 207854 486000
rect 209635 485348 209701 485349
rect 209635 485284 209636 485348
rect 209700 485284 209701 485348
rect 209635 485283 209701 485284
rect 208347 479500 208413 479501
rect 208347 479436 208348 479500
rect 208412 479436 208413 479500
rect 208347 479435 208413 479436
rect 207234 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 207854 477954
rect 207234 477634 207854 477718
rect 207234 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 207854 477634
rect 207059 474196 207125 474197
rect 207059 474132 207060 474196
rect 207124 474132 207125 474196
rect 207059 474131 207125 474132
rect 206691 415308 206757 415309
rect 206691 415244 206692 415308
rect 206756 415244 206757 415308
rect 206691 415243 206757 415244
rect 207062 378045 207122 474131
rect 207234 460894 207854 477398
rect 207979 465900 208045 465901
rect 207979 465836 207980 465900
rect 208044 465836 208045 465900
rect 207979 465835 208045 465836
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207059 378044 207125 378045
rect 207059 377980 207060 378044
rect 207124 377980 207125 378044
rect 207059 377979 207125 377980
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 206507 164932 206573 164933
rect 206507 164868 206508 164932
rect 206572 164868 206573 164932
rect 206507 164867 206573 164868
rect 206323 164116 206389 164117
rect 206323 164052 206324 164116
rect 206388 164052 206389 164116
rect 206323 164051 206389 164052
rect 207234 155834 207854 172338
rect 207982 166565 208042 465835
rect 208350 379541 208410 479435
rect 208899 467260 208965 467261
rect 208899 467196 208900 467260
rect 208964 467196 208965 467260
rect 208899 467195 208965 467196
rect 208347 379540 208413 379541
rect 208347 379476 208348 379540
rect 208412 379476 208413 379540
rect 208347 379475 208413 379476
rect 207979 166564 208045 166565
rect 207979 166500 207980 166564
rect 208044 166500 208045 166564
rect 207979 166499 208045 166500
rect 208902 165477 208962 467195
rect 208899 165476 208965 165477
rect 208899 165412 208900 165476
rect 208964 165412 208965 165476
rect 208899 165411 208965 165412
rect 207234 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 207854 155834
rect 207234 155514 207854 155598
rect 207234 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 207854 155514
rect 207234 136894 207854 155278
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 209638 58853 209698 485283
rect 210954 481674 211574 486000
rect 213683 485484 213749 485485
rect 213683 485420 213684 485484
rect 213748 485420 213749 485484
rect 213683 485419 213749 485420
rect 211659 485348 211725 485349
rect 211659 485284 211660 485348
rect 211724 485284 211725 485348
rect 211659 485283 211725 485284
rect 210954 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 211574 481674
rect 210954 481354 211574 481438
rect 210954 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 211574 481354
rect 210371 479500 210437 479501
rect 210371 479436 210372 479500
rect 210436 479436 210437 479500
rect 210371 479435 210437 479436
rect 209819 476916 209885 476917
rect 209819 476852 209820 476916
rect 209884 476852 209885 476916
rect 209819 476851 209885 476852
rect 209822 378725 209882 476851
rect 209819 378724 209885 378725
rect 209819 378660 209820 378724
rect 209884 378660 209885 378724
rect 209819 378659 209885 378660
rect 209635 58852 209701 58853
rect 209635 58788 209636 58852
rect 209700 58788 209701 58852
rect 209635 58787 209701 58788
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 206139 3228 206205 3229
rect 206139 3164 206140 3228
rect 206204 3164 206205 3228
rect 206139 3163 206205 3164
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 210374 4045 210434 479435
rect 210555 478276 210621 478277
rect 210555 478212 210556 478276
rect 210620 478212 210621 478276
rect 210555 478211 210621 478212
rect 210558 56677 210618 478211
rect 210954 464614 211574 481118
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 373674 211574 392058
rect 211662 378045 211722 485283
rect 212395 484804 212461 484805
rect 212395 484740 212396 484804
rect 212460 484740 212461 484804
rect 212395 484739 212461 484740
rect 211659 378044 211725 378045
rect 211659 377980 211660 378044
rect 211724 377980 211725 378044
rect 211659 377979 211725 377980
rect 210954 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 211574 373674
rect 210954 373354 211574 373438
rect 210954 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 211574 373354
rect 210954 356614 211574 373118
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 157674 211574 176058
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210555 56676 210621 56677
rect 210555 56612 210556 56676
rect 210620 56612 210621 56676
rect 210555 56611 210621 56612
rect 210954 32614 211574 68058
rect 212398 59125 212458 484739
rect 213315 478412 213381 478413
rect 213315 478348 213316 478412
rect 213380 478348 213381 478412
rect 213315 478347 213381 478348
rect 213131 478140 213197 478141
rect 213131 478076 213132 478140
rect 213196 478076 213197 478140
rect 213131 478075 213197 478076
rect 212395 59124 212461 59125
rect 212395 59060 212396 59124
rect 212460 59060 212461 59124
rect 212395 59059 212461 59060
rect 213134 57221 213194 478075
rect 213318 165205 213378 478347
rect 213499 468484 213565 468485
rect 213499 468420 213500 468484
rect 213564 468420 213565 468484
rect 213499 468419 213565 468420
rect 213502 166701 213562 468419
rect 213686 378045 213746 485419
rect 216995 485076 217061 485077
rect 216995 485012 216996 485076
rect 217060 485012 217061 485076
rect 216995 485011 217061 485012
rect 213867 483852 213933 483853
rect 213867 483788 213868 483852
rect 213932 483788 213933 483852
rect 213867 483787 213933 483788
rect 213683 378044 213749 378045
rect 213683 377980 213684 378044
rect 213748 377980 213749 378044
rect 213683 377979 213749 377980
rect 213870 376685 213930 483787
rect 214603 483716 214669 483717
rect 214603 483652 214604 483716
rect 214668 483652 214669 483716
rect 214603 483651 214669 483652
rect 214051 480860 214117 480861
rect 214051 480796 214052 480860
rect 214116 480796 214117 480860
rect 214051 480795 214117 480796
rect 214054 378045 214114 480795
rect 214419 476780 214485 476781
rect 214419 476716 214420 476780
rect 214484 476716 214485 476780
rect 214419 476715 214485 476716
rect 214051 378044 214117 378045
rect 214051 377980 214052 378044
rect 214116 377980 214117 378044
rect 214051 377979 214117 377980
rect 213867 376684 213933 376685
rect 213867 376620 213868 376684
rect 213932 376620 213933 376684
rect 213867 376619 213933 376620
rect 213499 166700 213565 166701
rect 213499 166636 213500 166700
rect 213564 166636 213565 166700
rect 213499 166635 213565 166636
rect 213315 165204 213381 165205
rect 213315 165140 213316 165204
rect 213380 165140 213381 165204
rect 213315 165139 213381 165140
rect 214422 57765 214482 476715
rect 214606 68101 214666 483651
rect 215339 482356 215405 482357
rect 215339 482292 215340 482356
rect 215404 482292 215405 482356
rect 215339 482291 215405 482292
rect 215342 375461 215402 482291
rect 215891 479636 215957 479637
rect 215891 479572 215892 479636
rect 215956 479572 215957 479636
rect 215891 479571 215957 479572
rect 215339 375460 215405 375461
rect 215339 375396 215340 375460
rect 215404 375396 215405 375460
rect 215339 375395 215405 375396
rect 214603 68100 214669 68101
rect 214603 68036 214604 68100
rect 214668 68036 214669 68100
rect 214603 68035 214669 68036
rect 214419 57764 214485 57765
rect 214419 57700 214420 57764
rect 214484 57700 214485 57764
rect 214419 57699 214485 57700
rect 213131 57220 213197 57221
rect 213131 57156 213132 57220
rect 213196 57156 213197 57220
rect 213131 57155 213197 57156
rect 215894 57085 215954 479571
rect 216075 474060 216141 474061
rect 216075 473996 216076 474060
rect 216140 473996 216141 474060
rect 216075 473995 216141 473996
rect 216078 57493 216138 473995
rect 216259 472836 216325 472837
rect 216259 472772 216260 472836
rect 216324 472772 216325 472836
rect 216259 472771 216325 472772
rect 216262 165069 216322 472771
rect 216998 380357 217058 485011
rect 217547 484532 217613 484533
rect 217547 484468 217548 484532
rect 217612 484468 217613 484532
rect 217547 484467 217613 484468
rect 217179 479772 217245 479773
rect 217179 479708 217180 479772
rect 217244 479708 217245 479772
rect 217179 479707 217245 479708
rect 216995 380356 217061 380357
rect 216995 380292 216996 380356
rect 217060 380292 217061 380356
rect 216995 380291 217061 380292
rect 216627 380220 216693 380221
rect 216627 380156 216628 380220
rect 216692 380156 216693 380220
rect 216627 380155 216693 380156
rect 216630 376549 216690 380155
rect 216627 376548 216693 376549
rect 216627 376484 216628 376548
rect 216692 376484 216693 376548
rect 216627 376483 216693 376484
rect 216995 376004 217061 376005
rect 216995 375940 216996 376004
rect 217060 375940 217061 376004
rect 216995 375939 217061 375940
rect 216998 252517 217058 375939
rect 217182 271557 217242 479707
rect 217363 471476 217429 471477
rect 217363 471412 217364 471476
rect 217428 471412 217429 471476
rect 217363 471411 217429 471412
rect 217366 272917 217426 471411
rect 217550 380490 217610 484467
rect 217794 471454 218414 486000
rect 219203 485076 219269 485077
rect 219203 485012 219204 485076
rect 219268 485012 219269 485076
rect 219203 485011 219269 485012
rect 218651 475556 218717 475557
rect 218651 475492 218652 475556
rect 218716 475492 218717 475556
rect 218651 475491 218717 475492
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 466308 218414 470898
rect 217915 380492 217981 380493
rect 217915 380490 217916 380492
rect 217550 380430 217916 380490
rect 217550 380221 217610 380430
rect 217915 380428 217916 380430
rect 217980 380428 217981 380492
rect 217915 380427 217981 380428
rect 217547 380220 217613 380221
rect 217547 380156 217548 380220
rect 217612 380156 217613 380220
rect 217547 380155 217613 380156
rect 217794 363454 218414 379000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 359308 218414 362898
rect 217363 272916 217429 272917
rect 217363 272852 217364 272916
rect 217428 272852 217429 272916
rect 217363 272851 217429 272852
rect 217179 271556 217245 271557
rect 217179 271492 217180 271556
rect 217244 271492 217245 271556
rect 217179 271491 217245 271492
rect 217547 270060 217613 270061
rect 217547 269996 217548 270060
rect 217612 269996 217613 270060
rect 217547 269995 217613 269996
rect 216995 252516 217061 252517
rect 216995 252452 216996 252516
rect 217060 252452 217061 252516
rect 216995 252451 217061 252452
rect 216998 248430 217058 252451
rect 216998 248370 217242 248430
rect 216259 165068 216325 165069
rect 216259 165004 216260 165068
rect 216324 165004 216325 165068
rect 216259 165003 216325 165004
rect 217182 162757 217242 248370
rect 217179 162756 217245 162757
rect 217179 162692 217180 162756
rect 217244 162692 217245 162756
rect 217179 162691 217245 162692
rect 217182 161490 217242 162691
rect 217182 161430 217426 161490
rect 217366 58445 217426 161430
rect 217550 146301 217610 269995
rect 217794 255454 218414 272000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 252308 218414 254898
rect 217794 147454 218414 165000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217547 146300 217613 146301
rect 217547 146236 217548 146300
rect 217612 146236 217613 146300
rect 217547 146235 217613 146236
rect 217794 145308 218414 146898
rect 218654 60621 218714 475491
rect 218835 467124 218901 467125
rect 218835 467060 218836 467124
rect 218900 467060 218901 467124
rect 218835 467059 218901 467060
rect 218838 273461 218898 467059
rect 218835 273460 218901 273461
rect 218835 273396 218836 273460
rect 218900 273396 218901 273460
rect 218835 273395 218901 273396
rect 219206 60621 219266 485011
rect 219939 484532 220005 484533
rect 219939 484468 219940 484532
rect 220004 484468 220005 484532
rect 219939 484467 220005 484468
rect 218651 60620 218717 60621
rect 218651 60556 218652 60620
rect 218716 60556 218717 60620
rect 218651 60555 218717 60556
rect 219203 60620 219269 60621
rect 219203 60556 219204 60620
rect 219268 60556 219269 60620
rect 219203 60555 219269 60556
rect 217363 58444 217429 58445
rect 217363 58380 217364 58444
rect 217428 58380 217429 58444
rect 217363 58379 217429 58380
rect 216075 57492 216141 57493
rect 216075 57428 216076 57492
rect 216140 57428 216141 57492
rect 216075 57427 216141 57428
rect 215891 57084 215957 57085
rect 215891 57020 215892 57084
rect 215956 57020 215957 57084
rect 215891 57019 215957 57020
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 210371 4044 210437 4045
rect 210371 3980 210372 4044
rect 210436 3980 210437 4044
rect 210371 3979 210437 3980
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219942 56541 220002 484467
rect 221514 475174 222134 486000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 466308 222134 474618
rect 225234 478894 225854 486000
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 466308 225854 478338
rect 228954 482614 229574 486000
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 466308 229574 482058
rect 235794 472394 236414 486000
rect 235794 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 236414 472394
rect 235794 472074 236414 472158
rect 235794 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 236414 472074
rect 235794 466308 236414 471838
rect 239514 476114 240134 486000
rect 239514 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 240134 476114
rect 239514 475794 240134 475878
rect 239514 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 240134 475794
rect 239514 466308 240134 475558
rect 243234 477954 243854 486000
rect 243234 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 243854 477954
rect 243234 477634 243854 477718
rect 243234 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 243854 477634
rect 243234 466308 243854 477398
rect 246954 481674 247574 486000
rect 246954 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 247574 481674
rect 246954 481354 247574 481438
rect 246954 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 247574 481354
rect 246954 466308 247574 481118
rect 253794 471454 254414 486000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 466308 254414 470898
rect 257514 475174 258134 486000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 466308 258134 474618
rect 261234 478894 261854 486000
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 466308 261854 478338
rect 264954 482614 265574 486000
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 466308 265574 482058
rect 271794 472394 272414 486000
rect 271794 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 271794 472074 272414 472158
rect 271794 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 271794 466308 272414 471838
rect 275514 476114 276134 486000
rect 275514 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 275514 475794 276134 475878
rect 275514 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 275514 466308 276134 475558
rect 279234 477954 279854 486000
rect 279234 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 279234 477634 279854 477718
rect 279234 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 279234 466308 279854 477398
rect 282954 481674 283574 486000
rect 282954 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 282954 481354 283574 481438
rect 282954 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 282954 466308 283574 481118
rect 289794 471454 290414 486000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 466308 290414 470898
rect 293514 475174 294134 486000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 466308 294134 474618
rect 297234 478894 297854 486000
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 466308 297854 478338
rect 300954 482614 301574 486000
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 466308 301574 482058
rect 307794 466308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 466308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 466308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 642033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 642033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 642033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 642033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 642033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 642033 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 642033 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 642033 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 642033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 642033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 642033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 642033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 642033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 642033 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 642033 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 642033 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 642033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 642033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 642033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 642033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 642033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 642033 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 642033 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 642033 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 642033 434414 650898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 344568 633454 344888 633486
rect 344568 633218 344610 633454
rect 344846 633218 344888 633454
rect 344568 633134 344888 633218
rect 344568 632898 344610 633134
rect 344846 632898 344888 633134
rect 344568 632866 344888 632898
rect 375288 633454 375608 633486
rect 375288 633218 375330 633454
rect 375566 633218 375608 633454
rect 375288 633134 375608 633218
rect 375288 632898 375330 633134
rect 375566 632898 375608 633134
rect 375288 632866 375608 632898
rect 406008 633454 406328 633486
rect 406008 633218 406050 633454
rect 406286 633218 406328 633454
rect 406008 633134 406328 633218
rect 406008 632898 406050 633134
rect 406286 632898 406328 633134
rect 406008 632866 406328 632898
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 329208 615454 329528 615486
rect 329208 615218 329250 615454
rect 329486 615218 329528 615454
rect 329208 615134 329528 615218
rect 329208 614898 329250 615134
rect 329486 614898 329528 615134
rect 329208 614866 329528 614898
rect 359928 615454 360248 615486
rect 359928 615218 359970 615454
rect 360206 615218 360248 615454
rect 359928 615134 360248 615218
rect 359928 614898 359970 615134
rect 360206 614898 360248 615134
rect 359928 614866 360248 614898
rect 390648 615454 390968 615486
rect 390648 615218 390690 615454
rect 390926 615218 390968 615454
rect 390648 615134 390968 615218
rect 390648 614898 390690 615134
rect 390926 614898 390968 615134
rect 390648 614866 390968 614898
rect 421368 615454 421688 615486
rect 421368 615218 421410 615454
rect 421646 615218 421688 615454
rect 421368 615134 421688 615218
rect 421368 614898 421410 615134
rect 421646 614898 421688 615134
rect 421368 614866 421688 614898
rect 436139 611420 436205 611421
rect 436139 611356 436140 611420
rect 436204 611356 436205 611420
rect 436139 611355 436205 611356
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 344568 597454 344888 597486
rect 344568 597218 344610 597454
rect 344846 597218 344888 597454
rect 344568 597134 344888 597218
rect 344568 596898 344610 597134
rect 344846 596898 344888 597134
rect 344568 596866 344888 596898
rect 375288 597454 375608 597486
rect 375288 597218 375330 597454
rect 375566 597218 375608 597454
rect 375288 597134 375608 597218
rect 375288 596898 375330 597134
rect 375566 596898 375608 597134
rect 375288 596866 375608 596898
rect 406008 597454 406328 597486
rect 406008 597218 406050 597454
rect 406286 597218 406328 597454
rect 406008 597134 406328 597218
rect 406008 596898 406050 597134
rect 406286 596898 406328 597134
rect 406008 596866 406328 596898
rect 329208 579454 329528 579486
rect 329208 579218 329250 579454
rect 329486 579218 329528 579454
rect 329208 579134 329528 579218
rect 329208 578898 329250 579134
rect 329486 578898 329528 579134
rect 329208 578866 329528 578898
rect 359928 579454 360248 579486
rect 359928 579218 359970 579454
rect 360206 579218 360248 579454
rect 359928 579134 360248 579218
rect 359928 578898 359970 579134
rect 360206 578898 360248 579134
rect 359928 578866 360248 578898
rect 390648 579454 390968 579486
rect 390648 579218 390690 579454
rect 390926 579218 390968 579454
rect 390648 579134 390968 579218
rect 390648 578898 390690 579134
rect 390926 578898 390968 579134
rect 390648 578866 390968 578898
rect 421368 579454 421688 579486
rect 421368 579218 421410 579454
rect 421646 579218 421688 579454
rect 421368 579134 421688 579218
rect 421368 578898 421410 579134
rect 421646 578898 421688 579134
rect 421368 578866 421688 578898
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 344568 561454 344888 561486
rect 344568 561218 344610 561454
rect 344846 561218 344888 561454
rect 344568 561134 344888 561218
rect 344568 560898 344610 561134
rect 344846 560898 344888 561134
rect 344568 560866 344888 560898
rect 375288 561454 375608 561486
rect 375288 561218 375330 561454
rect 375566 561218 375608 561454
rect 375288 561134 375608 561218
rect 375288 560898 375330 561134
rect 375566 560898 375608 561134
rect 375288 560866 375608 560898
rect 406008 561454 406328 561486
rect 406008 561218 406050 561454
rect 406286 561218 406328 561454
rect 406008 561134 406328 561218
rect 406008 560898 406050 561134
rect 406286 560898 406328 561134
rect 406008 560866 406328 560898
rect 324819 549540 324885 549541
rect 324819 549476 324820 549540
rect 324884 549476 324885 549540
rect 324819 549475 324885 549476
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 324822 529549 324882 549475
rect 329208 543454 329528 543486
rect 329208 543218 329250 543454
rect 329486 543218 329528 543454
rect 329208 543134 329528 543218
rect 329208 542898 329250 543134
rect 329486 542898 329528 543134
rect 329208 542866 329528 542898
rect 359928 543454 360248 543486
rect 359928 543218 359970 543454
rect 360206 543218 360248 543454
rect 359928 543134 360248 543218
rect 359928 542898 359970 543134
rect 360206 542898 360248 543134
rect 359928 542866 360248 542898
rect 390648 543454 390968 543486
rect 390648 543218 390690 543454
rect 390926 543218 390968 543454
rect 390648 543134 390968 543218
rect 390648 542898 390690 543134
rect 390926 542898 390968 543134
rect 390648 542866 390968 542898
rect 421368 543454 421688 543486
rect 421368 543218 421410 543454
rect 421646 543218 421688 543454
rect 421368 543134 421688 543218
rect 421368 542898 421410 543134
rect 421646 542898 421688 543134
rect 421368 542866 421688 542898
rect 324819 529548 324885 529549
rect 324819 529484 324820 529548
rect 324884 529484 324885 529548
rect 324819 529483 324885 529484
rect 436142 528189 436202 611355
rect 436323 606660 436389 606661
rect 436323 606596 436324 606660
rect 436388 606596 436389 606660
rect 436323 606595 436389 606596
rect 436326 528461 436386 606595
rect 436507 586532 436573 586533
rect 436507 586468 436508 586532
rect 436572 586468 436573 586532
rect 436507 586467 436573 586468
rect 436323 528460 436389 528461
rect 436323 528396 436324 528460
rect 436388 528396 436389 528460
rect 436323 528395 436389 528396
rect 436510 528325 436570 586467
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 436507 528324 436573 528325
rect 436507 528260 436508 528324
rect 436572 528260 436573 528324
rect 436507 528259 436573 528260
rect 436139 528188 436205 528189
rect 436139 528124 436140 528188
rect 436204 528124 436205 528188
rect 436139 528123 436205 528124
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 466308 319574 500058
rect 325794 507454 326414 527000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 466308 326414 470898
rect 329514 511174 330134 527000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 466308 330134 474618
rect 333234 514894 333854 527000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 466308 333854 478338
rect 336954 518614 337574 527000
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 466308 337574 482058
rect 343794 525454 344414 527000
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338435 466580 338501 466581
rect 338435 466516 338436 466580
rect 338500 466516 338501 466580
rect 338435 466515 338501 466516
rect 339723 466580 339789 466581
rect 339723 466516 339724 466580
rect 339788 466516 339789 466580
rect 339723 466515 339789 466516
rect 338438 464810 338498 466515
rect 339726 464810 339786 466515
rect 343794 466308 344414 488898
rect 347514 493174 348134 527000
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 466308 348134 492618
rect 351234 496894 351854 527000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 466580 351013 466581
rect 350947 466516 350948 466580
rect 351012 466516 351013 466580
rect 350947 466515 351013 466516
rect 350950 464810 351010 466515
rect 351234 466308 351854 496338
rect 354954 500614 355574 527000
rect 360699 518124 360765 518125
rect 360699 518060 360700 518124
rect 360764 518060 360765 518124
rect 360699 518059 360765 518060
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 466308 355574 500058
rect 357939 485620 358005 485621
rect 357939 485556 357940 485620
rect 358004 485556 358005 485620
rect 357939 485555 358005 485556
rect 338438 464750 338524 464810
rect 338464 464202 338524 464750
rect 339688 464750 339786 464810
rect 350840 464750 351010 464810
rect 339688 464202 339748 464750
rect 350840 464202 350900 464750
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 236056 380629 236116 381106
rect 237144 380629 237204 381106
rect 236053 380628 236119 380629
rect 236053 380564 236054 380628
rect 236118 380564 236119 380628
rect 236053 380563 236119 380564
rect 237141 380628 237207 380629
rect 237141 380564 237142 380628
rect 237206 380564 237207 380628
rect 237141 380563 237207 380564
rect 238232 380490 238292 381106
rect 239592 380490 239652 381106
rect 238158 380430 238292 380490
rect 239262 380430 239652 380490
rect 240544 380490 240604 381106
rect 241768 380490 241828 381106
rect 243128 380629 243188 381106
rect 243125 380628 243191 380629
rect 243125 380564 243126 380628
rect 243190 380564 243191 380628
rect 243125 380563 243191 380564
rect 244216 380490 244276 381106
rect 245440 380629 245500 381106
rect 245437 380628 245503 380629
rect 245437 380564 245438 380628
rect 245502 380564 245503 380628
rect 245437 380563 245503 380564
rect 246528 380490 246588 381106
rect 247616 380629 247676 381106
rect 248296 380901 248356 381106
rect 248293 380900 248359 380901
rect 248293 380836 248294 380900
rect 248358 380836 248359 380900
rect 248293 380835 248359 380836
rect 247613 380628 247679 380629
rect 247613 380564 247614 380628
rect 247678 380564 247679 380628
rect 247613 380563 247679 380564
rect 248704 380490 248764 381106
rect 240544 380430 240610 380490
rect 241768 380430 241898 380490
rect 244216 380430 244290 380490
rect 221514 367174 222134 379000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 359308 222134 366618
rect 225234 370894 225854 379000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 359308 225854 370338
rect 228954 374614 229574 379000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 359308 229574 374058
rect 235794 364394 236414 379000
rect 238158 378997 238218 380430
rect 238155 378996 238221 378997
rect 238155 378932 238156 378996
rect 238220 378932 238221 378996
rect 238155 378931 238221 378932
rect 239262 378861 239322 380430
rect 239259 378860 239325 378861
rect 239259 378796 239260 378860
rect 239324 378796 239325 378860
rect 239259 378795 239325 378796
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 359308 236414 363838
rect 239514 368114 240134 379000
rect 240550 378317 240610 380430
rect 241838 379133 241898 380430
rect 241835 379132 241901 379133
rect 241835 379068 241836 379132
rect 241900 379068 241901 379132
rect 241835 379067 241901 379068
rect 241467 378724 241533 378725
rect 241467 378660 241468 378724
rect 241532 378660 241533 378724
rect 241467 378659 241533 378660
rect 241470 378317 241530 378659
rect 241838 378453 241898 379067
rect 241835 378452 241901 378453
rect 241835 378388 241836 378452
rect 241900 378388 241901 378452
rect 241835 378387 241901 378388
rect 240547 378316 240613 378317
rect 240547 378252 240548 378316
rect 240612 378252 240613 378316
rect 240547 378251 240613 378252
rect 241467 378316 241533 378317
rect 241467 378252 241468 378316
rect 241532 378252 241533 378316
rect 241467 378251 241533 378252
rect 239514 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 240134 368114
rect 239514 367794 240134 367878
rect 239514 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 240134 367794
rect 239514 359308 240134 367558
rect 243234 369954 243854 379000
rect 244230 378317 244290 380430
rect 246438 380430 246588 380490
rect 248646 380430 248764 380490
rect 250064 380490 250124 381106
rect 250744 380898 250804 381106
rect 251288 380898 251348 381106
rect 250670 380838 250804 380898
rect 251222 380838 251348 380898
rect 250064 380430 250178 380490
rect 246438 379405 246498 380430
rect 248646 379405 248706 380430
rect 250118 379405 250178 380430
rect 246435 379404 246501 379405
rect 246435 379340 246436 379404
rect 246500 379340 246501 379404
rect 246435 379339 246501 379340
rect 248643 379404 248709 379405
rect 248643 379340 248644 379404
rect 248708 379340 248709 379404
rect 248643 379339 248709 379340
rect 250115 379404 250181 379405
rect 250115 379340 250116 379404
rect 250180 379340 250181 379404
rect 250115 379339 250181 379340
rect 244227 378316 244293 378317
rect 244227 378252 244228 378316
rect 244292 378252 244293 378316
rect 244227 378251 244293 378252
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 359308 243854 369398
rect 246954 373674 247574 379000
rect 250670 378317 250730 380838
rect 251222 379405 251282 380838
rect 252376 380490 252436 381106
rect 253464 380490 253524 381106
rect 252326 380430 252436 380490
rect 253430 380430 253524 380490
rect 253600 380490 253660 381106
rect 254552 380629 254612 381106
rect 255912 380629 255972 381106
rect 254549 380628 254615 380629
rect 254549 380564 254550 380628
rect 254614 380564 254615 380628
rect 254549 380563 254615 380564
rect 255909 380628 255975 380629
rect 255909 380564 255910 380628
rect 255974 380564 255975 380628
rect 255909 380563 255975 380564
rect 256048 380490 256108 381106
rect 257000 380629 257060 381106
rect 258088 380629 258148 381106
rect 256997 380628 257063 380629
rect 256997 380564 256998 380628
rect 257062 380564 257063 380628
rect 256997 380563 257063 380564
rect 258085 380628 258151 380629
rect 258085 380564 258086 380628
rect 258150 380564 258151 380628
rect 258085 380563 258151 380564
rect 258496 380490 258556 381106
rect 259448 380629 259508 381106
rect 260672 380629 260732 381106
rect 259445 380628 259511 380629
rect 259445 380564 259446 380628
rect 259510 380564 259511 380628
rect 259445 380563 259511 380564
rect 260669 380628 260735 380629
rect 260669 380564 260670 380628
rect 260734 380564 260735 380628
rect 260669 380563 260735 380564
rect 261080 380490 261140 381106
rect 261760 380490 261820 381106
rect 262848 380490 262908 381106
rect 253600 380430 253674 380490
rect 252326 379405 252386 380430
rect 253430 379405 253490 380430
rect 251219 379404 251285 379405
rect 251219 379340 251220 379404
rect 251284 379340 251285 379404
rect 251219 379339 251285 379340
rect 252323 379404 252389 379405
rect 252323 379340 252324 379404
rect 252388 379340 252389 379404
rect 252323 379339 252389 379340
rect 253427 379404 253493 379405
rect 253427 379340 253428 379404
rect 253492 379340 253493 379404
rect 253427 379339 253493 379340
rect 253614 378589 253674 380430
rect 256006 380430 256108 380490
rect 258398 380430 258556 380490
rect 260974 380430 261140 380490
rect 261710 380430 261820 380490
rect 262814 380430 262908 380490
rect 263528 380490 263588 381106
rect 263936 380490 263996 381106
rect 265296 380629 265356 381106
rect 265293 380628 265359 380629
rect 265293 380564 265294 380628
rect 265358 380564 265359 380628
rect 265293 380563 265359 380564
rect 265976 380490 266036 381106
rect 266384 380490 266444 381106
rect 267608 380490 267668 381106
rect 263528 380430 263610 380490
rect 253611 378588 253677 378589
rect 253611 378524 253612 378588
rect 253676 378524 253677 378588
rect 253611 378523 253677 378524
rect 250667 378316 250733 378317
rect 250667 378252 250668 378316
rect 250732 378252 250733 378316
rect 250667 378251 250733 378252
rect 246954 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 247574 373674
rect 246954 373354 247574 373438
rect 246954 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 247574 373354
rect 246954 359308 247574 373118
rect 253794 363454 254414 379000
rect 256006 378589 256066 380430
rect 256003 378588 256069 378589
rect 256003 378524 256004 378588
rect 256068 378524 256069 378588
rect 256003 378523 256069 378524
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 359308 254414 362898
rect 257514 367174 258134 379000
rect 258398 378589 258458 380430
rect 260974 378589 261034 380430
rect 261710 379405 261770 380430
rect 261707 379404 261773 379405
rect 261707 379340 261708 379404
rect 261772 379340 261773 379404
rect 261707 379339 261773 379340
rect 258395 378588 258461 378589
rect 258395 378524 258396 378588
rect 258460 378524 258461 378588
rect 258395 378523 258461 378524
rect 260971 378588 261037 378589
rect 260971 378524 260972 378588
rect 261036 378524 261037 378588
rect 260971 378523 261037 378524
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 359308 258134 366618
rect 261234 370894 261854 379000
rect 262814 378317 262874 380430
rect 263550 378589 263610 380430
rect 263918 380430 263996 380490
rect 265942 380430 266036 380490
rect 266310 380430 266444 380490
rect 267598 380430 267668 380490
rect 268288 380490 268348 381106
rect 268696 380490 268756 381106
rect 269784 380629 269844 381106
rect 271008 380629 271068 381106
rect 269781 380628 269847 380629
rect 269781 380564 269782 380628
rect 269846 380564 269847 380628
rect 269781 380563 269847 380564
rect 271005 380628 271071 380629
rect 271005 380564 271006 380628
rect 271070 380564 271071 380628
rect 271005 380563 271071 380564
rect 271144 380490 271204 381106
rect 272232 380490 272292 381106
rect 273320 380490 273380 381106
rect 273592 380490 273652 381106
rect 274408 380490 274468 381106
rect 275768 380490 275828 381106
rect 268288 380430 268394 380490
rect 268696 380430 268762 380490
rect 263918 379405 263978 380430
rect 263915 379404 263981 379405
rect 263915 379340 263916 379404
rect 263980 379340 263981 379404
rect 263915 379339 263981 379340
rect 263547 378588 263613 378589
rect 263547 378524 263548 378588
rect 263612 378524 263613 378588
rect 263547 378523 263613 378524
rect 262811 378316 262877 378317
rect 262811 378252 262812 378316
rect 262876 378252 262877 378316
rect 262811 378251 262877 378252
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 359308 261854 370338
rect 264954 374614 265574 379000
rect 265942 378589 266002 380430
rect 265939 378588 266005 378589
rect 265939 378524 265940 378588
rect 266004 378524 266005 378588
rect 265939 378523 266005 378524
rect 266310 378317 266370 380430
rect 267598 378317 267658 380430
rect 268334 378589 268394 380430
rect 268702 379405 268762 380430
rect 271094 380430 271204 380490
rect 272198 380430 272292 380490
rect 273302 380430 273380 380490
rect 273486 380430 273652 380490
rect 274406 380430 274468 380490
rect 275694 380430 275828 380490
rect 276040 380490 276100 381106
rect 276992 380490 277052 381106
rect 276040 380430 276122 380490
rect 271094 379405 271154 380430
rect 272198 379405 272258 380430
rect 273302 379405 273362 380430
rect 268699 379404 268765 379405
rect 268699 379340 268700 379404
rect 268764 379340 268765 379404
rect 268699 379339 268765 379340
rect 271091 379404 271157 379405
rect 271091 379340 271092 379404
rect 271156 379340 271157 379404
rect 271091 379339 271157 379340
rect 272195 379404 272261 379405
rect 272195 379340 272196 379404
rect 272260 379340 272261 379404
rect 272195 379339 272261 379340
rect 273299 379404 273365 379405
rect 273299 379340 273300 379404
rect 273364 379340 273365 379404
rect 273299 379339 273365 379340
rect 268331 378588 268397 378589
rect 268331 378524 268332 378588
rect 268396 378524 268397 378588
rect 268331 378523 268397 378524
rect 266307 378316 266373 378317
rect 266307 378252 266308 378316
rect 266372 378252 266373 378316
rect 266307 378251 266373 378252
rect 267595 378316 267661 378317
rect 267595 378252 267596 378316
rect 267660 378252 267661 378316
rect 267595 378251 267661 378252
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 359308 265574 374058
rect 271794 364394 272414 379000
rect 273486 378589 273546 380430
rect 274406 379405 274466 380430
rect 275694 379405 275754 380430
rect 276062 379405 276122 380430
rect 276982 380430 277052 380490
rect 278080 380490 278140 381106
rect 278488 380490 278548 381106
rect 279168 380765 279228 381106
rect 279165 380764 279231 380765
rect 279165 380700 279166 380764
rect 279230 380700 279231 380764
rect 279165 380699 279231 380700
rect 278080 380430 278146 380490
rect 276982 379405 277042 380430
rect 274403 379404 274469 379405
rect 274403 379340 274404 379404
rect 274468 379340 274469 379404
rect 274403 379339 274469 379340
rect 275691 379404 275757 379405
rect 275691 379340 275692 379404
rect 275756 379340 275757 379404
rect 275691 379339 275757 379340
rect 276059 379404 276125 379405
rect 276059 379340 276060 379404
rect 276124 379340 276125 379404
rect 276059 379339 276125 379340
rect 276979 379404 277045 379405
rect 276979 379340 276980 379404
rect 277044 379340 277045 379404
rect 276979 379339 277045 379340
rect 278086 379269 278146 380430
rect 278454 380430 278548 380490
rect 279168 380490 279228 380699
rect 280936 380490 280996 381106
rect 283520 380490 283580 381106
rect 279168 380430 279250 380490
rect 278454 379405 278514 380430
rect 279190 380221 279250 380430
rect 280846 380430 280996 380490
rect 283422 380430 283580 380490
rect 285968 380490 286028 381106
rect 288280 380490 288340 381106
rect 291000 380490 291060 381106
rect 293448 380490 293508 381106
rect 285968 380430 286058 380490
rect 279187 380220 279253 380221
rect 279187 380156 279188 380220
rect 279252 380156 279253 380220
rect 279187 380155 279253 380156
rect 278451 379404 278517 379405
rect 278451 379340 278452 379404
rect 278516 379340 278517 379404
rect 278451 379339 278517 379340
rect 280846 379269 280906 380430
rect 283422 379269 283482 380430
rect 285998 379405 286058 380430
rect 288206 380430 288340 380490
rect 290966 380430 291060 380490
rect 293358 380430 293508 380490
rect 295896 380490 295956 381106
rect 298480 380490 298540 381106
rect 300928 380490 300988 381106
rect 303512 380490 303572 381106
rect 305960 380490 306020 381106
rect 308544 380490 308604 381106
rect 295896 380430 295994 380490
rect 298480 380430 298570 380490
rect 288206 379405 288266 380430
rect 290966 379405 291026 380430
rect 293358 379405 293418 380430
rect 295934 379405 295994 380430
rect 298510 379405 298570 380430
rect 300902 380430 300988 380490
rect 303478 380430 303572 380490
rect 305870 380430 306020 380490
rect 308446 380430 308604 380490
rect 310992 380490 311052 381106
rect 313440 380490 313500 381106
rect 315888 380490 315948 381106
rect 318472 380490 318532 381106
rect 310992 380430 311082 380490
rect 300902 379405 300962 380430
rect 303478 379405 303538 380430
rect 305870 379405 305930 380430
rect 308446 379405 308506 380430
rect 311022 379405 311082 380430
rect 313414 380430 313500 380490
rect 315806 380430 315948 380490
rect 318382 380430 318532 380490
rect 320920 380490 320980 381106
rect 323368 380490 323428 381106
rect 325952 380490 326012 381106
rect 343224 380490 343284 381106
rect 320920 380430 321018 380490
rect 313414 379405 313474 380430
rect 315806 379405 315866 380430
rect 318382 379405 318442 380430
rect 285995 379404 286061 379405
rect 285995 379340 285996 379404
rect 286060 379340 286061 379404
rect 285995 379339 286061 379340
rect 288203 379404 288269 379405
rect 288203 379340 288204 379404
rect 288268 379340 288269 379404
rect 288203 379339 288269 379340
rect 290963 379404 291029 379405
rect 290963 379340 290964 379404
rect 291028 379340 291029 379404
rect 290963 379339 291029 379340
rect 293355 379404 293421 379405
rect 293355 379340 293356 379404
rect 293420 379340 293421 379404
rect 293355 379339 293421 379340
rect 295931 379404 295997 379405
rect 295931 379340 295932 379404
rect 295996 379340 295997 379404
rect 295931 379339 295997 379340
rect 298507 379404 298573 379405
rect 298507 379340 298508 379404
rect 298572 379340 298573 379404
rect 298507 379339 298573 379340
rect 300899 379404 300965 379405
rect 300899 379340 300900 379404
rect 300964 379340 300965 379404
rect 300899 379339 300965 379340
rect 303475 379404 303541 379405
rect 303475 379340 303476 379404
rect 303540 379340 303541 379404
rect 303475 379339 303541 379340
rect 305867 379404 305933 379405
rect 305867 379340 305868 379404
rect 305932 379340 305933 379404
rect 305867 379339 305933 379340
rect 308443 379404 308509 379405
rect 308443 379340 308444 379404
rect 308508 379340 308509 379404
rect 308443 379339 308509 379340
rect 311019 379404 311085 379405
rect 311019 379340 311020 379404
rect 311084 379340 311085 379404
rect 311019 379339 311085 379340
rect 313411 379404 313477 379405
rect 313411 379340 313412 379404
rect 313476 379340 313477 379404
rect 313411 379339 313477 379340
rect 315803 379404 315869 379405
rect 315803 379340 315804 379404
rect 315868 379340 315869 379404
rect 315803 379339 315869 379340
rect 318379 379404 318445 379405
rect 318379 379340 318380 379404
rect 318444 379340 318445 379404
rect 318379 379339 318445 379340
rect 278083 379268 278149 379269
rect 278083 379204 278084 379268
rect 278148 379204 278149 379268
rect 278083 379203 278149 379204
rect 280843 379268 280909 379269
rect 280843 379204 280844 379268
rect 280908 379204 280909 379268
rect 280843 379203 280909 379204
rect 283419 379268 283485 379269
rect 283419 379204 283420 379268
rect 283484 379204 283485 379268
rect 283419 379203 283485 379204
rect 273483 378588 273549 378589
rect 273483 378524 273484 378588
rect 273548 378524 273549 378588
rect 273483 378523 273549 378524
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 359308 272414 363838
rect 275514 368114 276134 379000
rect 275514 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 276134 368114
rect 275514 367794 276134 367878
rect 275514 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 276134 367794
rect 275514 359308 276134 367558
rect 279234 369954 279854 379000
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 359308 279854 369398
rect 282954 373674 283574 379000
rect 282954 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 283574 373674
rect 282954 373354 283574 373438
rect 282954 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 283574 373354
rect 282954 359308 283574 373118
rect 289794 363454 290414 379000
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 359308 290414 362898
rect 293514 367174 294134 379000
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 359308 294134 366618
rect 297234 370894 297854 379000
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 359308 297854 370338
rect 300954 374614 301574 379000
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 359308 301574 374058
rect 307794 364394 308414 379000
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 359308 308414 363838
rect 311514 368114 312134 379000
rect 311514 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 312134 368114
rect 311514 367794 312134 367878
rect 311514 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 312134 367794
rect 311514 359308 312134 367558
rect 315234 369954 315854 379000
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 359308 315854 369398
rect 318954 373674 319574 379000
rect 320958 378589 321018 380430
rect 323350 380430 323428 380490
rect 325926 380430 326012 380490
rect 343222 380430 343284 380490
rect 343360 380490 343420 381106
rect 343360 380430 343466 380490
rect 323350 380357 323410 380430
rect 323347 380356 323413 380357
rect 323347 380292 323348 380356
rect 323412 380292 323413 380356
rect 323347 380291 323413 380292
rect 325926 379269 325986 380430
rect 325923 379268 325989 379269
rect 325923 379204 325924 379268
rect 325988 379204 325989 379268
rect 325923 379203 325989 379204
rect 320955 378588 321021 378589
rect 320955 378524 320956 378588
rect 321020 378524 321021 378588
rect 320955 378523 321021 378524
rect 318954 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 319574 373674
rect 318954 373354 319574 373438
rect 318954 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 319574 373354
rect 318954 359308 319574 373118
rect 325794 363454 326414 379000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 359308 326414 362898
rect 329514 367174 330134 379000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 359308 330134 366618
rect 333234 370894 333854 379000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 359308 333854 370338
rect 336954 374614 337574 379000
rect 343222 378453 343282 380430
rect 343219 378452 343285 378453
rect 343219 378388 343220 378452
rect 343284 378388 343285 378452
rect 343219 378387 343285 378388
rect 343406 378317 343466 380430
rect 343403 378316 343469 378317
rect 343403 378252 343404 378316
rect 343468 378252 343469 378316
rect 343403 378251 343469 378252
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 359308 337574 374058
rect 343794 364394 344414 379000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 359308 344414 363838
rect 347514 368114 348134 379000
rect 347514 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 348134 368114
rect 347514 367794 348134 367878
rect 347514 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 348134 367794
rect 347514 359308 348134 367558
rect 351234 369954 351854 379000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 359308 351854 369398
rect 354954 373674 355574 379000
rect 354954 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 355574 373674
rect 354954 373354 355574 373438
rect 354954 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 355574 373354
rect 354954 359308 355574 373118
rect 338435 358868 338501 358869
rect 338435 358804 338436 358868
rect 338500 358804 338501 358868
rect 338435 358803 338501 358804
rect 339723 358868 339789 358869
rect 339723 358804 339724 358868
rect 339788 358804 339789 358868
rect 339723 358803 339789 358804
rect 350947 358868 351013 358869
rect 350947 358804 350948 358868
rect 351012 358804 351013 358868
rect 350947 358803 351013 358804
rect 338438 358050 338498 358803
rect 339726 358050 339786 358803
rect 350950 358050 351010 358803
rect 338438 357990 338524 358050
rect 338464 357202 338524 357990
rect 339688 357990 339786 358050
rect 350840 357990 351010 358050
rect 339688 357202 339748 357990
rect 350840 357202 350900 357990
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 236056 273730 236116 274040
rect 237144 273730 237204 274040
rect 238232 273730 238292 274040
rect 239592 273730 239652 274040
rect 236056 273670 236562 273730
rect 221514 259174 222134 272000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252308 222134 258618
rect 225234 262894 225854 272000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252308 225854 262338
rect 228954 266614 229574 272000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252308 229574 266058
rect 235794 256394 236414 272000
rect 236502 271421 236562 273670
rect 237054 273670 237204 273730
rect 238158 273670 238292 273730
rect 239262 273670 239652 273730
rect 240544 273730 240604 274040
rect 241768 273730 241828 274040
rect 243128 273730 243188 274040
rect 240544 273670 240610 273730
rect 236499 271420 236565 271421
rect 236499 271356 236500 271420
rect 236564 271356 236565 271420
rect 236499 271355 236565 271356
rect 237054 271285 237114 273670
rect 237051 271284 237117 271285
rect 237051 271220 237052 271284
rect 237116 271220 237117 271284
rect 237051 271219 237117 271220
rect 238158 270605 238218 273670
rect 238155 270604 238221 270605
rect 238155 270540 238156 270604
rect 238220 270540 238221 270604
rect 238155 270539 238221 270540
rect 239262 270333 239322 273670
rect 239259 270332 239325 270333
rect 239259 270268 239260 270332
rect 239324 270268 239325 270332
rect 239259 270267 239325 270268
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 252308 236414 255838
rect 239514 260114 240134 272000
rect 240550 269789 240610 273670
rect 241654 273670 241828 273730
rect 242942 273670 243188 273730
rect 244216 273730 244276 274040
rect 245440 273730 245500 274040
rect 246528 273730 246588 274040
rect 244216 273670 244290 273730
rect 241654 269925 241714 273670
rect 242942 270605 243002 273670
rect 242939 270604 243005 270605
rect 242939 270540 242940 270604
rect 243004 270540 243005 270604
rect 242939 270539 243005 270540
rect 241651 269924 241717 269925
rect 241651 269860 241652 269924
rect 241716 269860 241717 269924
rect 241651 269859 241717 269860
rect 240547 269788 240613 269789
rect 240547 269724 240548 269788
rect 240612 269724 240613 269788
rect 240547 269723 240613 269724
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 252308 240134 259558
rect 243234 261954 243854 272000
rect 244230 270741 244290 273670
rect 245334 273670 245500 273730
rect 246438 273670 246588 273730
rect 247616 273730 247676 274040
rect 248296 273730 248356 274040
rect 248704 273730 248764 274040
rect 247616 273670 247786 273730
rect 244227 270740 244293 270741
rect 244227 270676 244228 270740
rect 244292 270676 244293 270740
rect 244227 270675 244293 270676
rect 245334 270605 245394 273670
rect 246438 270605 246498 273670
rect 245331 270604 245397 270605
rect 245331 270540 245332 270604
rect 245396 270540 245397 270604
rect 245331 270539 245397 270540
rect 246435 270604 246501 270605
rect 246435 270540 246436 270604
rect 246500 270540 246501 270604
rect 246435 270539 246501 270540
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 252308 243854 261398
rect 246954 265674 247574 272000
rect 247726 270605 247786 273670
rect 248278 273670 248356 273730
rect 248646 273670 248764 273730
rect 250064 273730 250124 274040
rect 250744 273730 250804 274040
rect 251288 273730 251348 274040
rect 252376 273730 252436 274040
rect 253464 273730 253524 274040
rect 250064 273670 250178 273730
rect 248278 271149 248338 273670
rect 248275 271148 248341 271149
rect 248275 271084 248276 271148
rect 248340 271084 248341 271148
rect 248275 271083 248341 271084
rect 248646 270605 248706 273670
rect 250118 270605 250178 273670
rect 250670 273670 250804 273730
rect 251222 273670 251348 273730
rect 252326 273670 252436 273730
rect 253430 273670 253524 273730
rect 253600 273730 253660 274040
rect 254552 273730 254612 274040
rect 255912 273730 255972 274040
rect 253600 273670 253674 273730
rect 250670 273325 250730 273670
rect 250667 273324 250733 273325
rect 250667 273260 250668 273324
rect 250732 273260 250733 273324
rect 250667 273259 250733 273260
rect 251222 270605 251282 273670
rect 252326 270741 252386 273670
rect 252323 270740 252389 270741
rect 252323 270676 252324 270740
rect 252388 270676 252389 270740
rect 252323 270675 252389 270676
rect 253430 270605 253490 273670
rect 253614 271149 253674 273670
rect 254534 273670 254612 273730
rect 255822 273670 255972 273730
rect 256048 273730 256108 274040
rect 257000 273730 257060 274040
rect 256048 273670 256250 273730
rect 253611 271148 253677 271149
rect 253611 271084 253612 271148
rect 253676 271084 253677 271148
rect 253611 271083 253677 271084
rect 247723 270604 247789 270605
rect 247723 270540 247724 270604
rect 247788 270540 247789 270604
rect 247723 270539 247789 270540
rect 248643 270604 248709 270605
rect 248643 270540 248644 270604
rect 248708 270540 248709 270604
rect 248643 270539 248709 270540
rect 250115 270604 250181 270605
rect 250115 270540 250116 270604
rect 250180 270540 250181 270604
rect 250115 270539 250181 270540
rect 251219 270604 251285 270605
rect 251219 270540 251220 270604
rect 251284 270540 251285 270604
rect 251219 270539 251285 270540
rect 253427 270604 253493 270605
rect 253427 270540 253428 270604
rect 253492 270540 253493 270604
rect 253427 270539 253493 270540
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 252308 247574 265118
rect 253794 255454 254414 272000
rect 254534 270877 254594 273670
rect 254531 270876 254597 270877
rect 254531 270812 254532 270876
rect 254596 270812 254597 270876
rect 254531 270811 254597 270812
rect 255822 270741 255882 273670
rect 256190 271149 256250 273670
rect 256926 273670 257060 273730
rect 258088 273730 258148 274040
rect 258496 273730 258556 274040
rect 258088 273670 258274 273730
rect 256187 271148 256253 271149
rect 256187 271084 256188 271148
rect 256252 271084 256253 271148
rect 256187 271083 256253 271084
rect 255819 270740 255885 270741
rect 255819 270676 255820 270740
rect 255884 270676 255885 270740
rect 255819 270675 255885 270676
rect 256926 270605 256986 273670
rect 256923 270604 256989 270605
rect 256923 270540 256924 270604
rect 256988 270540 256989 270604
rect 256923 270539 256989 270540
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252308 254414 254898
rect 257514 259174 258134 272000
rect 258214 271010 258274 273670
rect 258398 273670 258556 273730
rect 259448 273730 259508 274040
rect 260672 273730 260732 274040
rect 261080 273730 261140 274040
rect 259448 273670 259562 273730
rect 258398 271285 258458 273670
rect 258395 271284 258461 271285
rect 258395 271220 258396 271284
rect 258460 271220 258461 271284
rect 258395 271219 258461 271220
rect 258214 270950 258458 271010
rect 258398 270605 258458 270950
rect 259502 270605 259562 273670
rect 260606 273670 260732 273730
rect 260974 273670 261140 273730
rect 261760 273730 261820 274040
rect 262848 273730 262908 274040
rect 261760 273670 262138 273730
rect 260606 270741 260666 273670
rect 260974 271285 261034 273670
rect 260971 271284 261037 271285
rect 260971 271220 260972 271284
rect 261036 271220 261037 271284
rect 260971 271219 261037 271220
rect 260603 270740 260669 270741
rect 260603 270676 260604 270740
rect 260668 270676 260669 270740
rect 260603 270675 260669 270676
rect 258395 270604 258461 270605
rect 258395 270540 258396 270604
rect 258460 270540 258461 270604
rect 258395 270539 258461 270540
rect 259499 270604 259565 270605
rect 259499 270540 259500 270604
rect 259564 270540 259565 270604
rect 259499 270539 259565 270540
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252308 258134 258618
rect 261234 262894 261854 272000
rect 262078 270605 262138 273670
rect 262814 273670 262908 273730
rect 263528 273730 263588 274040
rect 263936 273730 263996 274040
rect 265296 273730 265356 274040
rect 265976 273730 266036 274040
rect 263528 273670 263610 273730
rect 262814 270605 262874 273670
rect 263550 271829 263610 273670
rect 263918 273670 263996 273730
rect 265206 273670 265356 273730
rect 265942 273670 266036 273730
rect 263547 271828 263613 271829
rect 263547 271764 263548 271828
rect 263612 271764 263613 271828
rect 263547 271763 263613 271764
rect 263918 270605 263978 273670
rect 265206 272237 265266 273670
rect 265203 272236 265269 272237
rect 265203 272172 265204 272236
rect 265268 272172 265269 272236
rect 265203 272171 265269 272172
rect 262075 270604 262141 270605
rect 262075 270540 262076 270604
rect 262140 270540 262141 270604
rect 262075 270539 262141 270540
rect 262811 270604 262877 270605
rect 262811 270540 262812 270604
rect 262876 270540 262877 270604
rect 262811 270539 262877 270540
rect 263915 270604 263981 270605
rect 263915 270540 263916 270604
rect 263980 270540 263981 270604
rect 263915 270539 263981 270540
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252308 261854 262338
rect 264954 266614 265574 272000
rect 265942 271829 266002 273670
rect 266384 273597 266444 274040
rect 267608 273730 267668 274040
rect 267598 273670 267668 273730
rect 268288 273730 268348 274040
rect 268696 273730 268756 274040
rect 269784 273730 269844 274040
rect 271008 273730 271068 274040
rect 268288 273670 268394 273730
rect 268696 273670 268762 273730
rect 269784 273670 269866 273730
rect 266381 273596 266447 273597
rect 266381 273532 266382 273596
rect 266446 273532 266447 273596
rect 266381 273531 266447 273532
rect 265939 271828 266005 271829
rect 265939 271764 265940 271828
rect 266004 271764 266005 271828
rect 265939 271763 266005 271764
rect 267598 270605 267658 273670
rect 268334 271829 268394 273670
rect 268331 271828 268397 271829
rect 268331 271764 268332 271828
rect 268396 271764 268397 271828
rect 268331 271763 268397 271764
rect 268702 270877 268762 273670
rect 268699 270876 268765 270877
rect 268699 270812 268700 270876
rect 268764 270812 268765 270876
rect 268699 270811 268765 270812
rect 269806 270605 269866 273670
rect 270910 273670 271068 273730
rect 271144 273730 271204 274040
rect 272232 273730 272292 274040
rect 273320 273730 273380 274040
rect 273592 273730 273652 274040
rect 274408 273730 274468 274040
rect 275768 273730 275828 274040
rect 271144 273670 271338 273730
rect 272232 273670 272626 273730
rect 270910 271829 270970 273670
rect 270907 271828 270973 271829
rect 270907 271764 270908 271828
rect 270972 271764 270973 271828
rect 270907 271763 270973 271764
rect 271278 271285 271338 273670
rect 271275 271284 271341 271285
rect 271275 271220 271276 271284
rect 271340 271220 271341 271284
rect 271275 271219 271341 271220
rect 267595 270604 267661 270605
rect 267595 270540 267596 270604
rect 267660 270540 267661 270604
rect 267595 270539 267661 270540
rect 269803 270604 269869 270605
rect 269803 270540 269804 270604
rect 269868 270540 269869 270604
rect 269803 270539 269869 270540
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252308 265574 266058
rect 271794 256394 272414 272000
rect 272566 271829 272626 273670
rect 273302 273670 273380 273730
rect 273486 273670 273652 273730
rect 274406 273670 274468 273730
rect 275326 273670 275828 273730
rect 276040 273730 276100 274040
rect 276992 273730 277052 274040
rect 276040 273670 276306 273730
rect 273302 273461 273362 273670
rect 273299 273460 273365 273461
rect 273299 273396 273300 273460
rect 273364 273396 273365 273460
rect 273299 273395 273365 273396
rect 272563 271828 272629 271829
rect 272563 271764 272564 271828
rect 272628 271764 272629 271828
rect 272563 271763 272629 271764
rect 273486 271557 273546 273670
rect 273483 271556 273549 271557
rect 273483 271492 273484 271556
rect 273548 271492 273549 271556
rect 273483 271491 273549 271492
rect 274406 270605 274466 273670
rect 275326 270605 275386 273670
rect 274403 270604 274469 270605
rect 274403 270540 274404 270604
rect 274468 270540 274469 270604
rect 274403 270539 274469 270540
rect 275323 270604 275389 270605
rect 275323 270540 275324 270604
rect 275388 270540 275389 270604
rect 275323 270539 275389 270540
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 252308 272414 255838
rect 275514 260114 276134 272000
rect 276246 271829 276306 273670
rect 276982 273670 277052 273730
rect 278080 273730 278140 274040
rect 278488 273730 278548 274040
rect 279168 273730 279228 274040
rect 280936 273730 280996 274040
rect 278080 273670 278146 273730
rect 276243 271828 276309 271829
rect 276243 271764 276244 271828
rect 276308 271764 276309 271828
rect 276243 271763 276309 271764
rect 276982 271557 277042 273670
rect 276979 271556 277045 271557
rect 276979 271492 276980 271556
rect 277044 271492 277045 271556
rect 276979 271491 277045 271492
rect 278086 270877 278146 273670
rect 278454 273670 278548 273730
rect 279006 273670 279228 273730
rect 280846 273670 280996 273730
rect 278454 271829 278514 273670
rect 279006 271829 279066 273670
rect 278451 271828 278517 271829
rect 278451 271764 278452 271828
rect 278516 271764 278517 271828
rect 278451 271763 278517 271764
rect 279003 271828 279069 271829
rect 279003 271764 279004 271828
rect 279068 271764 279069 271828
rect 279003 271763 279069 271764
rect 278083 270876 278149 270877
rect 278083 270812 278084 270876
rect 278148 270812 278149 270876
rect 278083 270811 278149 270812
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 252308 276134 259558
rect 279234 261954 279854 272000
rect 280846 271829 280906 273670
rect 283520 273597 283580 274040
rect 285968 273730 286028 274040
rect 288280 273730 288340 274040
rect 291000 273730 291060 274040
rect 293448 273730 293508 274040
rect 285968 273670 286058 273730
rect 283517 273596 283583 273597
rect 283517 273532 283518 273596
rect 283582 273532 283583 273596
rect 283517 273531 283583 273532
rect 285998 272917 286058 273670
rect 288206 273670 288340 273730
rect 290966 273670 291060 273730
rect 293358 273670 293508 273730
rect 295896 273730 295956 274040
rect 298480 273730 298540 274040
rect 300928 273730 300988 274040
rect 303512 273730 303572 274040
rect 305960 273730 306020 274040
rect 295896 273670 295994 273730
rect 298480 273670 298570 273730
rect 288206 272917 288266 273670
rect 290966 272917 291026 273670
rect 285995 272916 286061 272917
rect 285995 272852 285996 272916
rect 286060 272852 286061 272916
rect 285995 272851 286061 272852
rect 288203 272916 288269 272917
rect 288203 272852 288204 272916
rect 288268 272852 288269 272916
rect 288203 272851 288269 272852
rect 290963 272916 291029 272917
rect 290963 272852 290964 272916
rect 291028 272852 291029 272916
rect 290963 272851 291029 272852
rect 293358 272781 293418 273670
rect 295934 272917 295994 273670
rect 295931 272916 295997 272917
rect 295931 272852 295932 272916
rect 295996 272852 295997 272916
rect 295931 272851 295997 272852
rect 298510 272781 298570 273670
rect 300902 273670 300988 273730
rect 303478 273670 303572 273730
rect 305870 273670 306020 273730
rect 308544 273730 308604 274040
rect 310992 273730 311052 274040
rect 313440 273730 313500 274040
rect 315888 273730 315948 274040
rect 318472 273730 318532 274040
rect 308544 273670 308690 273730
rect 310992 273670 311082 273730
rect 300902 272781 300962 273670
rect 303478 272917 303538 273670
rect 303475 272916 303541 272917
rect 303475 272852 303476 272916
rect 303540 272852 303541 272916
rect 303475 272851 303541 272852
rect 293355 272780 293421 272781
rect 293355 272716 293356 272780
rect 293420 272716 293421 272780
rect 293355 272715 293421 272716
rect 298507 272780 298573 272781
rect 298507 272716 298508 272780
rect 298572 272716 298573 272780
rect 298507 272715 298573 272716
rect 300899 272780 300965 272781
rect 300899 272716 300900 272780
rect 300964 272716 300965 272780
rect 300899 272715 300965 272716
rect 305870 272645 305930 273670
rect 305867 272644 305933 272645
rect 305867 272580 305868 272644
rect 305932 272580 305933 272644
rect 305867 272579 305933 272580
rect 280843 271828 280909 271829
rect 280843 271764 280844 271828
rect 280908 271764 280909 271828
rect 280843 271763 280909 271764
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 252308 279854 261398
rect 282954 265674 283574 272000
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 252308 283574 265118
rect 289794 255454 290414 272000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252308 290414 254898
rect 293514 259174 294134 272000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252308 294134 258618
rect 297234 262894 297854 272000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252308 297854 262338
rect 300954 266614 301574 272000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252308 301574 266058
rect 307794 256394 308414 272000
rect 308630 271829 308690 273670
rect 311022 273053 311082 273670
rect 313414 273670 313500 273730
rect 315070 273670 315948 273730
rect 318382 273670 318532 273730
rect 320920 273730 320980 274040
rect 323368 273730 323428 274040
rect 325952 273730 326012 274040
rect 343224 273730 343284 274040
rect 320920 273670 321018 273730
rect 311019 273052 311085 273053
rect 311019 272988 311020 273052
rect 311084 272988 311085 273052
rect 311019 272987 311085 272988
rect 308627 271828 308693 271829
rect 308627 271764 308628 271828
rect 308692 271764 308693 271828
rect 308627 271763 308693 271764
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 252308 308414 255838
rect 311514 260114 312134 272000
rect 313414 271829 313474 273670
rect 313411 271828 313477 271829
rect 313411 271764 313412 271828
rect 313476 271764 313477 271828
rect 313411 271763 313477 271764
rect 315070 271693 315130 273670
rect 318382 273189 318442 273670
rect 318379 273188 318445 273189
rect 318379 273124 318380 273188
rect 318444 273124 318445 273188
rect 318379 273123 318445 273124
rect 320958 272645 321018 273670
rect 323350 273670 323428 273730
rect 325742 273670 326012 273730
rect 343222 273670 343284 273730
rect 343360 273730 343420 274040
rect 343360 273670 343466 273730
rect 320955 272644 321021 272645
rect 320955 272580 320956 272644
rect 321020 272580 321021 272644
rect 320955 272579 321021 272580
rect 315067 271692 315133 271693
rect 315067 271628 315068 271692
rect 315132 271628 315133 271692
rect 315067 271627 315133 271628
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 252308 312134 259558
rect 315234 261954 315854 272000
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 252308 315854 261398
rect 318954 265674 319574 272000
rect 323350 270469 323410 273670
rect 325742 272370 325802 273670
rect 325558 272310 325802 272370
rect 325558 271013 325618 272310
rect 325555 271012 325621 271013
rect 325555 270948 325556 271012
rect 325620 270948 325621 271012
rect 325555 270947 325621 270948
rect 323347 270468 323413 270469
rect 323347 270404 323348 270468
rect 323412 270404 323413 270468
rect 323347 270403 323413 270404
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 252308 319574 265118
rect 325794 255454 326414 272000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252308 326414 254898
rect 329514 259174 330134 272000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252308 330134 258618
rect 333234 262894 333854 272000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252308 333854 262338
rect 336954 266614 337574 272000
rect 343222 271421 343282 273670
rect 343406 271557 343466 273670
rect 343403 271556 343469 271557
rect 343403 271492 343404 271556
rect 343468 271492 343469 271556
rect 343403 271491 343469 271492
rect 343219 271420 343285 271421
rect 343219 271356 343220 271420
rect 343284 271356 343285 271420
rect 343219 271355 343285 271356
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252308 337574 266058
rect 343794 256394 344414 272000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 338435 253604 338501 253605
rect 338435 253540 338436 253604
rect 338500 253540 338501 253604
rect 338435 253539 338501 253540
rect 338438 250610 338498 253539
rect 339723 253060 339789 253061
rect 339723 252996 339724 253060
rect 339788 252996 339789 253060
rect 339723 252995 339789 252996
rect 339726 250610 339786 252995
rect 343794 252308 344414 255838
rect 347514 260114 348134 272000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 252308 348134 259558
rect 351234 261954 351854 272000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 350947 253196 351013 253197
rect 350947 253132 350948 253196
rect 351012 253132 351013 253196
rect 350947 253131 351013 253132
rect 350950 250610 351010 253131
rect 351234 252308 351854 261398
rect 354954 265674 355574 272000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 252308 355574 265118
rect 338438 250550 338524 250610
rect 338464 250240 338524 250550
rect 339688 250550 339786 250610
rect 350840 250550 351010 250610
rect 339688 250240 339748 250550
rect 350840 250240 350900 250550
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 166290 236116 167106
rect 237144 166290 237204 167106
rect 238232 166290 238292 167106
rect 235950 166230 236116 166290
rect 237054 166230 237204 166290
rect 238158 166230 238292 166290
rect 239592 166290 239652 167106
rect 240544 166290 240604 167106
rect 241768 166290 241828 167106
rect 243128 166290 243188 167106
rect 244216 167010 244276 167106
rect 245440 167010 245500 167106
rect 246528 167010 246588 167106
rect 247616 167010 247676 167106
rect 248296 167010 248356 167106
rect 248704 167010 248764 167106
rect 244216 166950 244474 167010
rect 244216 166910 244290 166950
rect 239592 166230 239690 166290
rect 240544 166230 240610 166290
rect 235950 165613 236010 166230
rect 235947 165612 236013 165613
rect 235947 165548 235948 165612
rect 236012 165548 236013 165612
rect 235947 165547 236013 165548
rect 221514 151174 222134 165000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 165000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 165000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 165000
rect 237054 164253 237114 166230
rect 238158 164253 238218 166230
rect 239630 165613 239690 166230
rect 239627 165612 239693 165613
rect 239627 165548 239628 165612
rect 239692 165548 239693 165612
rect 239627 165547 239693 165548
rect 237051 164252 237117 164253
rect 237051 164188 237052 164252
rect 237116 164188 237117 164252
rect 237051 164187 237117 164188
rect 238155 164252 238221 164253
rect 238155 164188 238156 164252
rect 238220 164188 238221 164252
rect 238155 164187 238221 164188
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 165000
rect 240550 164253 240610 166230
rect 241654 166230 241828 166290
rect 243126 166230 243188 166290
rect 241654 164253 241714 166230
rect 243126 165613 243186 166230
rect 243123 165612 243189 165613
rect 243123 165548 243124 165612
rect 243188 165548 243189 165612
rect 243123 165547 243189 165548
rect 240547 164252 240613 164253
rect 240547 164188 240548 164252
rect 240612 164188 240613 164252
rect 240547 164187 240613 164188
rect 241651 164252 241717 164253
rect 241651 164188 241652 164252
rect 241716 164188 241717 164252
rect 241651 164187 241717 164188
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 155834 243854 165000
rect 244414 164525 244474 166950
rect 245334 166950 245500 167010
rect 246438 166950 246588 167010
rect 247542 166950 247676 167010
rect 248278 166950 248356 167010
rect 248646 166950 248764 167010
rect 250064 167010 250124 167106
rect 250744 167010 250804 167106
rect 251288 167010 251348 167106
rect 252376 167010 252436 167106
rect 253464 167010 253524 167106
rect 250064 166950 250178 167010
rect 244411 164524 244477 164525
rect 244411 164460 244412 164524
rect 244476 164460 244477 164524
rect 244411 164459 244477 164460
rect 245334 164253 245394 166950
rect 246438 164253 246498 166950
rect 247542 165613 247602 166950
rect 248278 165613 248338 166950
rect 247539 165612 247605 165613
rect 247539 165548 247540 165612
rect 247604 165548 247605 165612
rect 247539 165547 247605 165548
rect 248275 165612 248341 165613
rect 248275 165548 248276 165612
rect 248340 165548 248341 165612
rect 248275 165547 248341 165548
rect 245331 164252 245397 164253
rect 245331 164188 245332 164252
rect 245396 164188 245397 164252
rect 245331 164187 245397 164188
rect 246435 164252 246501 164253
rect 246435 164188 246436 164252
rect 246500 164188 246501 164252
rect 246435 164187 246501 164188
rect 243234 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 243854 155834
rect 243234 155514 243854 155598
rect 243234 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 243854 155514
rect 243234 145308 243854 155278
rect 246954 157674 247574 165000
rect 248646 164253 248706 166950
rect 250118 164253 250178 166950
rect 250670 166950 250804 167010
rect 251222 166950 251348 167010
rect 252326 166950 252436 167010
rect 253430 166950 253524 167010
rect 253600 167010 253660 167106
rect 254552 167010 254612 167106
rect 255912 167010 255972 167106
rect 253600 166950 253674 167010
rect 250670 165613 250730 166950
rect 250667 165612 250733 165613
rect 250667 165548 250668 165612
rect 250732 165548 250733 165612
rect 250667 165547 250733 165548
rect 251222 164253 251282 166950
rect 252326 164525 252386 166950
rect 252323 164524 252389 164525
rect 252323 164460 252324 164524
rect 252388 164460 252389 164524
rect 252323 164459 252389 164460
rect 253430 164253 253490 166950
rect 253614 165613 253674 166950
rect 254534 166950 254612 167010
rect 255822 166950 255972 167010
rect 256048 167010 256108 167106
rect 257000 167010 257060 167106
rect 256048 166950 256250 167010
rect 253611 165612 253677 165613
rect 253611 165548 253612 165612
rect 253676 165548 253677 165612
rect 253611 165547 253677 165548
rect 248643 164252 248709 164253
rect 248643 164188 248644 164252
rect 248708 164188 248709 164252
rect 248643 164187 248709 164188
rect 250115 164252 250181 164253
rect 250115 164188 250116 164252
rect 250180 164188 250181 164252
rect 250115 164187 250181 164188
rect 251219 164252 251285 164253
rect 251219 164188 251220 164252
rect 251284 164188 251285 164252
rect 251219 164187 251285 164188
rect 253427 164252 253493 164253
rect 253427 164188 253428 164252
rect 253492 164188 253493 164252
rect 253427 164187 253493 164188
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 165000
rect 254534 164253 254594 166950
rect 255822 164253 255882 166950
rect 256190 164797 256250 166950
rect 256926 166950 257060 167010
rect 258088 167010 258148 167106
rect 258496 167010 258556 167106
rect 258088 166950 258274 167010
rect 256187 164796 256253 164797
rect 256187 164732 256188 164796
rect 256252 164732 256253 164796
rect 256187 164731 256253 164732
rect 256926 164253 256986 166950
rect 254531 164252 254597 164253
rect 254531 164188 254532 164252
rect 254596 164188 254597 164252
rect 254531 164187 254597 164188
rect 255819 164252 255885 164253
rect 255819 164188 255820 164252
rect 255884 164188 255885 164252
rect 255819 164187 255885 164188
rect 256923 164252 256989 164253
rect 256923 164188 256924 164252
rect 256988 164188 256989 164252
rect 256923 164187 256989 164188
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 165000
rect 258214 164250 258274 166950
rect 258398 166950 258556 167010
rect 259448 167010 259508 167106
rect 260672 167010 260732 167106
rect 261080 167010 261140 167106
rect 261760 167010 261820 167106
rect 262848 167010 262908 167106
rect 259448 166950 259562 167010
rect 258398 165613 258458 166950
rect 258395 165612 258461 165613
rect 258395 165548 258396 165612
rect 258460 165548 258461 165612
rect 258395 165547 258461 165548
rect 259502 164253 259562 166950
rect 260606 166950 260732 167010
rect 260974 166950 261140 167010
rect 261710 166950 261820 167010
rect 262814 166950 262908 167010
rect 263528 167010 263588 167106
rect 263936 167010 263996 167106
rect 265296 167010 265356 167106
rect 265976 167010 266036 167106
rect 263528 166950 263794 167010
rect 260606 164525 260666 166950
rect 260974 166429 261034 166950
rect 260971 166428 261037 166429
rect 260971 166364 260972 166428
rect 261036 166364 261037 166428
rect 260971 166363 261037 166364
rect 261710 165613 261770 166950
rect 261707 165612 261773 165613
rect 261707 165548 261708 165612
rect 261772 165548 261773 165612
rect 261707 165547 261773 165548
rect 260603 164524 260669 164525
rect 260603 164460 260604 164524
rect 260668 164460 260669 164524
rect 260603 164459 260669 164460
rect 258395 164252 258461 164253
rect 258395 164250 258396 164252
rect 258214 164190 258396 164250
rect 258395 164188 258396 164190
rect 258460 164188 258461 164252
rect 258395 164187 258461 164188
rect 259499 164252 259565 164253
rect 259499 164188 259500 164252
rect 259564 164188 259565 164252
rect 259499 164187 259565 164188
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 165000
rect 262814 164253 262874 166950
rect 263734 164933 263794 166950
rect 263918 166950 263996 167010
rect 265206 166950 265356 167010
rect 265942 166950 266036 167010
rect 266384 167010 266444 167106
rect 267608 167010 267668 167106
rect 266384 166950 266554 167010
rect 263731 164932 263797 164933
rect 263731 164868 263732 164932
rect 263796 164868 263797 164932
rect 263731 164867 263797 164868
rect 263918 164253 263978 166950
rect 265206 165613 265266 166950
rect 265942 166429 266002 166950
rect 265939 166428 266005 166429
rect 265939 166364 265940 166428
rect 266004 166364 266005 166428
rect 265939 166363 266005 166364
rect 265203 165612 265269 165613
rect 265203 165548 265204 165612
rect 265268 165548 265269 165612
rect 265203 165547 265269 165548
rect 262811 164252 262877 164253
rect 262811 164188 262812 164252
rect 262876 164188 262877 164252
rect 262811 164187 262877 164188
rect 263915 164252 263981 164253
rect 263915 164188 263916 164252
rect 263980 164188 263981 164252
rect 263915 164187 263981 164188
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 165000
rect 266494 164525 266554 166950
rect 267598 166950 267668 167010
rect 268288 167010 268348 167106
rect 268696 167010 268756 167106
rect 269784 167010 269844 167106
rect 271008 167010 271068 167106
rect 268288 166950 268394 167010
rect 268696 166950 268762 167010
rect 269784 166950 269866 167010
rect 267598 164661 267658 166950
rect 268334 165613 268394 166950
rect 268331 165612 268397 165613
rect 268331 165548 268332 165612
rect 268396 165548 268397 165612
rect 268331 165547 268397 165548
rect 267595 164660 267661 164661
rect 267595 164596 267596 164660
rect 267660 164596 267661 164660
rect 267595 164595 267661 164596
rect 266491 164524 266557 164525
rect 266491 164460 266492 164524
rect 266556 164460 266557 164524
rect 266491 164459 266557 164460
rect 268702 164253 268762 166950
rect 269806 164253 269866 166950
rect 270910 166950 271068 167010
rect 271144 167010 271204 167106
rect 272232 167010 272292 167106
rect 273320 167010 273380 167106
rect 273592 167010 273652 167106
rect 274408 167010 274468 167106
rect 271144 166950 271338 167010
rect 270910 166293 270970 166950
rect 270907 166292 270973 166293
rect 270907 166228 270908 166292
rect 270972 166228 270973 166292
rect 270907 166227 270973 166228
rect 271278 164253 271338 166950
rect 272198 166950 272292 167010
rect 273302 166950 273380 167010
rect 273486 166950 273652 167010
rect 274406 166950 274468 167010
rect 275768 167010 275828 167106
rect 276040 167010 276100 167106
rect 276992 167010 277052 167106
rect 275768 166950 275938 167010
rect 276040 166950 276122 167010
rect 272198 165613 272258 166950
rect 272195 165612 272261 165613
rect 272195 165548 272196 165612
rect 272260 165548 272261 165612
rect 272195 165547 272261 165548
rect 268699 164252 268765 164253
rect 268699 164188 268700 164252
rect 268764 164188 268765 164252
rect 268699 164187 268765 164188
rect 269803 164252 269869 164253
rect 269803 164188 269804 164252
rect 269868 164188 269869 164252
rect 269803 164187 269869 164188
rect 271275 164252 271341 164253
rect 271275 164188 271276 164252
rect 271340 164188 271341 164252
rect 271275 164187 271341 164188
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 165000
rect 273302 164525 273362 166950
rect 273486 165613 273546 166950
rect 273483 165612 273549 165613
rect 273483 165548 273484 165612
rect 273548 165548 273549 165612
rect 273483 165547 273549 165548
rect 273299 164524 273365 164525
rect 273299 164460 273300 164524
rect 273364 164460 273365 164524
rect 273299 164459 273365 164460
rect 274406 164253 274466 166950
rect 275878 165613 275938 166950
rect 276062 165613 276122 166950
rect 276982 166950 277052 167010
rect 278080 167010 278140 167106
rect 278488 167010 278548 167106
rect 278080 166950 278146 167010
rect 275875 165612 275941 165613
rect 275875 165548 275876 165612
rect 275940 165548 275941 165612
rect 275875 165547 275941 165548
rect 276059 165612 276125 165613
rect 276059 165548 276060 165612
rect 276124 165548 276125 165612
rect 276059 165547 276125 165548
rect 274403 164252 274469 164253
rect 274403 164188 274404 164252
rect 274468 164188 274469 164252
rect 274403 164187 274469 164188
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 165000
rect 276982 164253 277042 166950
rect 278086 164253 278146 166950
rect 278454 166950 278548 167010
rect 279168 167010 279228 167106
rect 280936 167010 280996 167106
rect 279168 166950 279250 167010
rect 278454 165613 278514 166950
rect 279190 165613 279250 166950
rect 280846 166950 280996 167010
rect 280846 165613 280906 166950
rect 283520 166290 283580 167106
rect 285968 166565 286028 167106
rect 288280 166565 288340 167106
rect 291000 166565 291060 167106
rect 293448 166565 293508 167106
rect 295896 166565 295956 167106
rect 298480 166701 298540 167106
rect 298477 166700 298543 166701
rect 298477 166636 298478 166700
rect 298542 166636 298543 166700
rect 298477 166635 298543 166636
rect 285965 166564 286031 166565
rect 285965 166500 285966 166564
rect 286030 166500 286031 166564
rect 285965 166499 286031 166500
rect 288277 166564 288343 166565
rect 288277 166500 288278 166564
rect 288342 166500 288343 166564
rect 288277 166499 288343 166500
rect 290997 166564 291063 166565
rect 290997 166500 290998 166564
rect 291062 166500 291063 166564
rect 290997 166499 291063 166500
rect 293445 166564 293511 166565
rect 293445 166500 293446 166564
rect 293510 166500 293511 166564
rect 293445 166499 293511 166500
rect 295893 166564 295959 166565
rect 295893 166500 295894 166564
rect 295958 166500 295959 166564
rect 295893 166499 295959 166500
rect 300928 166290 300988 167106
rect 303512 166701 303572 167106
rect 305960 166837 306020 167106
rect 305957 166836 306023 166837
rect 305957 166772 305958 166836
rect 306022 166772 306023 166836
rect 308544 166834 308604 167106
rect 310992 166834 311052 167106
rect 313440 166837 313500 167106
rect 313437 166836 313503 166837
rect 308544 166774 308690 166834
rect 310992 166774 311082 166834
rect 305957 166771 306023 166772
rect 303509 166700 303575 166701
rect 303509 166636 303510 166700
rect 303574 166636 303575 166700
rect 303509 166635 303575 166636
rect 283422 166230 283580 166290
rect 300902 166230 300988 166290
rect 283422 165613 283482 166230
rect 300902 165613 300962 166230
rect 278451 165612 278517 165613
rect 278451 165548 278452 165612
rect 278516 165548 278517 165612
rect 278451 165547 278517 165548
rect 279187 165612 279253 165613
rect 279187 165548 279188 165612
rect 279252 165548 279253 165612
rect 279187 165547 279253 165548
rect 280843 165612 280909 165613
rect 280843 165548 280844 165612
rect 280908 165548 280909 165612
rect 280843 165547 280909 165548
rect 283419 165612 283485 165613
rect 283419 165548 283420 165612
rect 283484 165548 283485 165612
rect 283419 165547 283485 165548
rect 300899 165612 300965 165613
rect 300899 165548 300900 165612
rect 300964 165548 300965 165612
rect 300899 165547 300965 165548
rect 308630 165069 308690 166774
rect 311022 165205 311082 166774
rect 313437 166772 313438 166836
rect 313502 166772 313503 166836
rect 315888 166834 315948 167106
rect 318472 166834 318532 167106
rect 313437 166771 313503 166772
rect 315806 166774 315948 166834
rect 318382 166774 318532 166834
rect 320920 166834 320980 167106
rect 323368 166834 323428 167106
rect 320920 166774 321018 166834
rect 315806 165341 315866 166774
rect 315803 165340 315869 165341
rect 315803 165276 315804 165340
rect 315868 165276 315869 165340
rect 315803 165275 315869 165276
rect 311019 165204 311085 165205
rect 311019 165140 311020 165204
rect 311084 165140 311085 165204
rect 311019 165139 311085 165140
rect 308627 165068 308693 165069
rect 308627 165004 308628 165068
rect 308692 165004 308693 165068
rect 308627 165003 308693 165004
rect 276979 164252 277045 164253
rect 276979 164188 276980 164252
rect 277044 164188 277045 164252
rect 276979 164187 277045 164188
rect 278083 164252 278149 164253
rect 278083 164188 278084 164252
rect 278148 164188 278149 164252
rect 278083 164187 278149 164188
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 155834 279854 165000
rect 279234 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 279854 155834
rect 279234 155514 279854 155598
rect 279234 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 279854 155514
rect 279234 145308 279854 155278
rect 282954 157674 283574 165000
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 165000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 165000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 165000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 165000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 165000
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 165000
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 155834 315854 165000
rect 318382 164253 318442 166774
rect 318379 164252 318445 164253
rect 318379 164188 318380 164252
rect 318444 164188 318445 164252
rect 318379 164187 318445 164188
rect 315234 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 315854 155834
rect 315234 155514 315854 155598
rect 315234 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 315854 155514
rect 315234 145308 315854 155278
rect 318954 157674 319574 165000
rect 320958 164389 321018 166774
rect 323350 166774 323428 166834
rect 323350 165613 323410 166774
rect 325952 166290 326012 167106
rect 343224 166290 343284 167106
rect 325926 166230 326012 166290
rect 343222 166230 343284 166290
rect 343360 166290 343420 167106
rect 343360 166230 343466 166290
rect 323347 165612 323413 165613
rect 323347 165548 323348 165612
rect 323412 165548 323413 165612
rect 323347 165547 323413 165548
rect 325926 165477 325986 166230
rect 343222 165477 343282 166230
rect 343406 165613 343466 166230
rect 343403 165612 343469 165613
rect 343403 165548 343404 165612
rect 343468 165548 343469 165612
rect 343403 165547 343469 165548
rect 325923 165476 325989 165477
rect 325923 165412 325924 165476
rect 325988 165412 325989 165476
rect 325923 165411 325989 165412
rect 343219 165476 343285 165477
rect 343219 165412 343220 165476
rect 343284 165412 343285 165476
rect 343219 165411 343285 165412
rect 320955 164388 321021 164389
rect 320955 164324 320956 164388
rect 321020 164324 321021 164388
rect 320955 164323 321021 164324
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 165000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 165000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 165000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 165000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 165000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 165000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 155834 351854 165000
rect 351234 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 351854 155834
rect 351234 155514 351854 155598
rect 351234 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 351854 155514
rect 351234 145308 351854 155278
rect 354954 157674 355574 165000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59530 236116 60106
rect 237144 59805 237204 60106
rect 237141 59804 237207 59805
rect 237141 59740 237142 59804
rect 237206 59740 237207 59804
rect 237141 59739 237207 59740
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 235950 59470 236116 59530
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 235950 58173 236010 59470
rect 235947 58172 236013 58173
rect 235947 58108 235948 58172
rect 236012 58108 236013 58172
rect 235947 58107 236013 58108
rect 219939 56540 220005 56541
rect 219939 56476 219940 56540
rect 220004 56476 220005 56540
rect 219939 56475 220005 56476
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57901 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57901 241714 59470
rect 242942 57901 243002 59470
rect 240547 57900 240613 57901
rect 240547 57836 240548 57900
rect 240612 57836 240613 57900
rect 240547 57835 240613 57836
rect 241651 57900 241717 57901
rect 241651 57836 241652 57900
rect 241716 57836 241717 57900
rect 241651 57835 241717 57836
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57901 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 244227 57900 244293 57901
rect 244227 57836 244228 57900
rect 244292 57836 244293 57900
rect 244227 57835 244293 57836
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57901 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59666 250804 60106
rect 251288 59666 251348 60106
rect 250670 59606 250804 59666
rect 251222 59606 251348 59666
rect 250064 59470 250178 59530
rect 248278 57901 248338 59470
rect 248646 57901 248706 59470
rect 250118 57901 250178 59470
rect 250670 58581 250730 59606
rect 250667 58580 250733 58581
rect 250667 58516 250668 58580
rect 250732 58516 250733 58580
rect 250667 58515 250733 58516
rect 251222 57901 251282 59606
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59805 257060 60106
rect 256997 59804 257063 59805
rect 256997 59740 256998 59804
rect 257062 59740 257063 59804
rect 256997 59739 257063 59740
rect 258088 59669 258148 60106
rect 258085 59668 258151 59669
rect 258085 59604 258086 59668
rect 258150 59604 258151 59668
rect 258085 59603 258151 59604
rect 258496 59530 258556 60106
rect 253600 59470 253674 59530
rect 252326 57901 252386 59470
rect 253430 57901 253490 59470
rect 253614 58717 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 258398 59470 258556 59530
rect 259448 59530 259508 60106
rect 260672 59669 260732 60106
rect 260669 59668 260735 59669
rect 260669 59604 260670 59668
rect 260734 59604 260735 59668
rect 260669 59603 260735 59604
rect 261080 59530 261140 60106
rect 261760 59669 261820 60106
rect 262848 59805 262908 60106
rect 262845 59804 262911 59805
rect 262845 59740 262846 59804
rect 262910 59740 262911 59804
rect 262845 59739 262911 59740
rect 261757 59668 261823 59669
rect 261757 59604 261758 59668
rect 261822 59604 261823 59668
rect 261757 59603 261823 59604
rect 259448 59470 259562 59530
rect 253611 58716 253677 58717
rect 253611 58652 253612 58716
rect 253676 58652 253677 58716
rect 253611 58651 253677 58652
rect 247723 57900 247789 57901
rect 247723 57836 247724 57900
rect 247788 57836 247789 57900
rect 247723 57835 247789 57836
rect 248275 57900 248341 57901
rect 248275 57836 248276 57900
rect 248340 57836 248341 57900
rect 248275 57835 248341 57836
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250115 57900 250181 57901
rect 250115 57836 250116 57900
rect 250180 57836 250181 57900
rect 250115 57835 250181 57836
rect 251219 57900 251285 57901
rect 251219 57836 251220 57900
rect 251284 57836 251285 57900
rect 251219 57835 251285 57836
rect 252323 57900 252389 57901
rect 252323 57836 252324 57900
rect 252388 57836 252389 57900
rect 252323 57835 252389 57836
rect 253427 57900 253493 57901
rect 253427 57836 253428 57900
rect 253492 57836 253493 57900
rect 253427 57835 253493 57836
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57901 254594 59470
rect 254531 57900 254597 57901
rect 254531 57836 254532 57900
rect 254596 57836 254597 57900
rect 254531 57835 254597 57836
rect 256006 57357 256066 59470
rect 256003 57356 256069 57357
rect 256003 57292 256004 57356
rect 256068 57292 256069 57356
rect 256003 57291 256069 57292
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 258398 57901 258458 59470
rect 259502 58445 259562 59470
rect 260974 59470 261140 59530
rect 263528 59530 263588 60106
rect 263936 59805 263996 60106
rect 263933 59804 263999 59805
rect 263933 59740 263934 59804
rect 263998 59740 263999 59804
rect 263933 59739 263999 59740
rect 265296 59530 265356 60106
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263528 59470 263610 59530
rect 259499 58444 259565 58445
rect 259499 58380 259500 58444
rect 259564 58380 259565 58444
rect 259499 58379 259565 58380
rect 258395 57900 258461 57901
rect 258395 57836 258396 57900
rect 258460 57836 258461 57900
rect 258395 57835 258461 57836
rect 260974 57085 261034 59470
rect 263550 59397 263610 59470
rect 265206 59470 265356 59530
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59666 271068 60106
rect 270910 59606 271068 59666
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 263547 59396 263613 59397
rect 263547 59332 263548 59396
rect 263612 59332 263613 59396
rect 263547 59331 263613 59332
rect 265206 58173 265266 59470
rect 265203 58172 265269 58173
rect 265203 58108 265204 58172
rect 265268 58108 265269 58172
rect 265203 58107 265269 58108
rect 260971 57084 261037 57085
rect 260971 57020 260972 57084
rect 261036 57020 261037 57084
rect 260971 57019 261037 57020
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57221 266002 59470
rect 266310 57357 266370 59470
rect 267598 57901 267658 59470
rect 267595 57900 267661 57901
rect 267595 57836 267596 57900
rect 267660 57836 267661 57900
rect 267595 57835 267661 57836
rect 266307 57356 266373 57357
rect 266307 57292 266308 57356
rect 266372 57292 266373 57356
rect 266307 57291 266373 57292
rect 265939 57220 266005 57221
rect 265939 57156 265940 57220
rect 266004 57156 266005 57220
rect 265939 57155 266005 57156
rect 268334 56405 268394 59470
rect 268702 57901 268762 59470
rect 268699 57900 268765 57901
rect 268699 57836 268700 57900
rect 268764 57836 268765 57900
rect 268699 57835 268765 57836
rect 269806 57629 269866 59470
rect 270910 57901 270970 59606
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59666 273652 60106
rect 271094 59470 271204 59530
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59606 273652 59666
rect 271094 57901 271154 59470
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 270907 57900 270973 57901
rect 270907 57836 270908 57900
rect 270972 57836 270973 57900
rect 270907 57835 270973 57836
rect 271091 57900 271157 57901
rect 271091 57836 271092 57900
rect 271156 57836 271157 57900
rect 271091 57835 271157 57836
rect 269803 57628 269869 57629
rect 269803 57564 269804 57628
rect 269868 57564 269869 57628
rect 269803 57563 269869 57564
rect 271794 57454 272414 58000
rect 273302 57901 273362 59470
rect 273486 58989 273546 59606
rect 274408 59530 274468 60106
rect 275768 59666 275828 60106
rect 274406 59470 274468 59530
rect 275694 59606 275828 59666
rect 273483 58988 273549 58989
rect 273483 58924 273484 58988
rect 273548 58924 273549 58988
rect 273483 58923 273549 58924
rect 273299 57900 273365 57901
rect 273299 57836 273300 57900
rect 273364 57836 273365 57900
rect 273299 57835 273365 57836
rect 274406 57629 274466 59470
rect 275694 58173 275754 59606
rect 276040 59530 276100 60106
rect 276992 59530 277052 60106
rect 276040 59470 276122 59530
rect 276062 58853 276122 59470
rect 276982 59470 277052 59530
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 278080 59470 278146 59530
rect 276059 58852 276125 58853
rect 276059 58788 276060 58852
rect 276124 58788 276125 58852
rect 276059 58787 276125 58788
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57628 274469 57629
rect 274403 57564 274404 57628
rect 274468 57564 274469 57628
rect 274403 57563 274469 57564
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 268331 56404 268397 56405
rect 268331 56340 268332 56404
rect 268396 56340 268397 56404
rect 268331 56339 268397 56340
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 57901 277042 59470
rect 276979 57900 277045 57901
rect 276979 57836 276980 57900
rect 277044 57836 277045 57900
rect 276979 57835 277045 57836
rect 278086 57629 278146 59470
rect 278454 59470 278548 59530
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 279168 59470 279250 59530
rect 278454 57901 278514 59470
rect 279190 59397 279250 59470
rect 280846 59470 280996 59530
rect 283520 59530 283580 60106
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 283520 59470 283850 59530
rect 285968 59470 286058 59530
rect 279187 59396 279253 59397
rect 279187 59332 279188 59396
rect 279252 59332 279253 59396
rect 279187 59331 279253 59332
rect 280846 59261 280906 59470
rect 280843 59260 280909 59261
rect 280843 59196 280844 59260
rect 280908 59196 280909 59260
rect 280843 59195 280909 59196
rect 278451 57900 278517 57901
rect 278451 57836 278452 57900
rect 278516 57836 278517 57900
rect 278451 57835 278517 57836
rect 278083 57628 278149 57629
rect 278083 57564 278084 57628
rect 278148 57564 278149 57628
rect 278083 57563 278149 57564
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 283790 57493 283850 59470
rect 285998 59125 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59530 306020 60106
rect 308544 59669 308604 60106
rect 308541 59668 308607 59669
rect 308541 59604 308542 59668
rect 308606 59604 308607 59668
rect 308541 59603 308607 59604
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 285995 59124 286061 59125
rect 285995 59060 285996 59124
rect 286060 59060 286061 59124
rect 285995 59059 286061 59060
rect 288206 57765 288266 59470
rect 290966 59261 291026 59470
rect 290963 59260 291029 59261
rect 290963 59196 290964 59260
rect 291028 59196 291029 59260
rect 290963 59195 291029 59196
rect 288203 57764 288269 57765
rect 288203 57700 288204 57764
rect 288268 57700 288269 57764
rect 288203 57699 288269 57700
rect 283787 57492 283853 57493
rect 283787 57428 283788 57492
rect 283852 57428 283853 57492
rect 283787 57427 283853 57428
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 56677 293418 59470
rect 293355 56676 293421 56677
rect 293355 56612 293356 56676
rect 293420 56612 293421 56676
rect 293355 56611 293421 56612
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 295934 57901 295994 59470
rect 295931 57900 295997 57901
rect 295931 57836 295932 57900
rect 295996 57836 295997 57900
rect 295931 57835 295997 57836
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 298510 57901 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 305870 59470 306020 59530
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59669 315948 60106
rect 315885 59668 315951 59669
rect 315885 59604 315886 59668
rect 315950 59604 315951 59668
rect 318472 59666 318532 60106
rect 315885 59603 315951 59604
rect 318382 59606 318532 59666
rect 310992 59470 311082 59530
rect 300902 59261 300962 59470
rect 300899 59260 300965 59261
rect 300899 59196 300900 59260
rect 300964 59196 300965 59260
rect 300899 59195 300965 59196
rect 298507 57900 298573 57901
rect 298507 57836 298508 57900
rect 298572 57836 298573 57900
rect 298507 57835 298573 57836
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 303478 57901 303538 59470
rect 305870 57901 305930 59470
rect 303475 57900 303541 57901
rect 303475 57836 303476 57900
rect 303540 57836 303541 57900
rect 303475 57835 303541 57836
rect 305867 57900 305933 57901
rect 305867 57836 305868 57900
rect 305932 57836 305933 57900
rect 305867 57835 305933 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 313414 57901 313474 59470
rect 313411 57900 313477 57901
rect 313411 57836 313412 57900
rect 313476 57836 313477 57900
rect 313411 57835 313477 57836
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 318382 57901 318442 59606
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 320958 59261 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 320955 59260 321021 59261
rect 320955 59196 320956 59260
rect 321020 59196 321021 59260
rect 320955 59195 321021 59196
rect 318379 57900 318445 57901
rect 318379 57836 318380 57900
rect 318444 57836 318445 57900
rect 318379 57835 318445 57836
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 323350 57901 323410 59470
rect 325926 59261 325986 59470
rect 325923 59260 325989 59261
rect 325923 59196 325924 59260
rect 325988 59196 325989 59260
rect 325923 59195 325989 59196
rect 323347 57900 323413 57901
rect 323347 57836 323348 57900
rect 323412 57836 323413 57900
rect 323347 57835 323413 57836
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 357942 59261 358002 485555
rect 359411 482492 359477 482493
rect 359411 482428 359412 482492
rect 359476 482428 359477 482492
rect 359411 482427 359477 482428
rect 358123 478276 358189 478277
rect 358123 478212 358124 478276
rect 358188 478212 358189 478276
rect 358123 478211 358189 478212
rect 357939 59260 358005 59261
rect 357939 59196 357940 59260
rect 358004 59196 358005 59260
rect 357939 59195 358005 59196
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 358126 56677 358186 478211
rect 359414 273189 359474 482427
rect 359595 479772 359661 479773
rect 359595 479708 359596 479772
rect 359660 479708 359661 479772
rect 359595 479707 359661 479708
rect 359598 380221 359658 479707
rect 359779 475692 359845 475693
rect 359779 475628 359780 475692
rect 359844 475628 359845 475692
rect 359779 475627 359845 475628
rect 359782 380901 359842 475627
rect 360147 475556 360213 475557
rect 360147 475492 360148 475556
rect 360212 475492 360213 475556
rect 360147 475491 360213 475492
rect 359963 465900 360029 465901
rect 359963 465836 359964 465900
rect 360028 465836 360029 465900
rect 359963 465835 360029 465836
rect 359779 380900 359845 380901
rect 359779 380836 359780 380900
rect 359844 380836 359845 380900
rect 359779 380835 359845 380836
rect 359595 380220 359661 380221
rect 359595 380156 359596 380220
rect 359660 380156 359661 380220
rect 359595 380155 359661 380156
rect 359966 376685 360026 465835
rect 360150 378045 360210 475491
rect 360147 378044 360213 378045
rect 360147 377980 360148 378044
rect 360212 377980 360213 378044
rect 360147 377979 360213 377980
rect 359963 376684 360029 376685
rect 359963 376620 359964 376684
rect 360028 376620 360029 376684
rect 359963 376619 360029 376620
rect 359411 273188 359477 273189
rect 359411 273124 359412 273188
rect 359476 273124 359477 273188
rect 359411 273123 359477 273124
rect 358123 56676 358189 56677
rect 358123 56612 358124 56676
rect 358188 56612 358189 56676
rect 358123 56611 358189 56612
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 360702 3773 360762 518059
rect 361794 507454 362414 527000
rect 363459 523700 363525 523701
rect 363459 523636 363460 523700
rect 363524 523636 363525 523700
rect 363459 523635 363525 523636
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 363462 149157 363522 523635
rect 365514 511174 366134 527000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 364931 487796 364997 487797
rect 364931 487732 364932 487796
rect 364996 487732 364997 487796
rect 364931 487731 364997 487732
rect 363459 149156 363525 149157
rect 363459 149092 363460 149156
rect 363524 149092 363525 149156
rect 363459 149091 363525 149092
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 360699 3772 360765 3773
rect 360699 3708 360700 3772
rect 360764 3708 360765 3772
rect 360699 3707 360765 3708
rect 361794 3454 362414 38898
rect 364934 3637 364994 487731
rect 365115 486572 365181 486573
rect 365115 486508 365116 486572
rect 365180 486508 365181 486572
rect 365115 486507 365181 486508
rect 364931 3636 364997 3637
rect 364931 3572 364932 3636
rect 364996 3572 364997 3636
rect 364931 3571 364997 3572
rect 365118 3501 365178 486507
rect 365514 475174 366134 510618
rect 369234 514894 369854 527000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 367691 489156 367757 489157
rect 367691 489092 367692 489156
rect 367756 489092 367757 489156
rect 367691 489091 367757 489092
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 366955 472836 367021 472837
rect 366955 472772 366956 472836
rect 367020 472772 367021 472836
rect 366955 472771 367021 472772
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 365115 3500 365181 3501
rect 365115 3436 365116 3500
rect 365180 3436 365181 3500
rect 365115 3435 365181 3436
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 6618
rect 366958 3229 367018 472771
rect 367694 3365 367754 489091
rect 367875 485484 367941 485485
rect 367875 485420 367876 485484
rect 367940 485420 367941 485484
rect 367875 485419 367941 485420
rect 367878 58989 367938 485419
rect 369234 478894 369854 514338
rect 372954 518614 373574 527000
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 371739 485348 371805 485349
rect 371739 485284 371740 485348
rect 371804 485284 371805 485348
rect 371739 485283 371805 485284
rect 370451 483852 370517 483853
rect 370451 483788 370452 483852
rect 370516 483788 370517 483852
rect 370451 483787 370517 483788
rect 370083 480860 370149 480861
rect 370083 480796 370084 480860
rect 370148 480796 370149 480860
rect 370083 480795 370149 480796
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 370086 377909 370146 480795
rect 370083 377908 370149 377909
rect 370083 377844 370084 377908
rect 370148 377844 370149 377908
rect 370083 377843 370149 377844
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 367875 58988 367941 58989
rect 367875 58924 367876 58988
rect 367940 58924 367941 58988
rect 367875 58923 367941 58924
rect 369234 46894 369854 82338
rect 370454 57629 370514 483787
rect 370635 465764 370701 465765
rect 370635 465700 370636 465764
rect 370700 465700 370701 465764
rect 370635 465699 370701 465700
rect 370638 166973 370698 465699
rect 370635 166972 370701 166973
rect 370635 166908 370636 166972
rect 370700 166908 370701 166972
rect 370635 166907 370701 166908
rect 371742 59125 371802 485283
rect 372954 482614 373574 518058
rect 379794 525454 380414 527000
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 375971 485212 376037 485213
rect 375971 485148 375972 485212
rect 376036 485148 376037 485212
rect 375971 485147 376037 485148
rect 374683 485076 374749 485077
rect 374683 485012 374684 485076
rect 374748 485012 374749 485076
rect 374683 485011 374749 485012
rect 374499 483716 374565 483717
rect 374499 483652 374500 483716
rect 374564 483652 374565 483716
rect 374499 483651 374565 483652
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 371923 472700 371989 472701
rect 371923 472636 371924 472700
rect 371988 472636 371989 472700
rect 371923 472635 371989 472636
rect 371739 59124 371805 59125
rect 371739 59060 371740 59124
rect 371804 59060 371805 59124
rect 371739 59059 371805 59060
rect 370451 57628 370517 57629
rect 370451 57564 370452 57628
rect 370516 57564 370517 57628
rect 370451 57563 370517 57564
rect 371926 57357 371986 472635
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 371923 57356 371989 57357
rect 371923 57292 371924 57356
rect 371988 57292 371989 57356
rect 371923 57291 371989 57292
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 367691 3364 367757 3365
rect 367691 3300 367692 3364
rect 367756 3300 367757 3364
rect 367691 3299 367757 3300
rect 366955 3228 367021 3229
rect 366955 3164 366956 3228
rect 367020 3164 367021 3228
rect 366955 3163 367021 3164
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 86058
rect 374502 57765 374562 483651
rect 374686 58717 374746 485011
rect 375419 482356 375485 482357
rect 375419 482292 375420 482356
rect 375484 482292 375485 482356
rect 375419 482291 375485 482292
rect 375422 68917 375482 482291
rect 375419 68916 375485 68917
rect 375419 68852 375420 68916
rect 375484 68852 375485 68916
rect 375419 68851 375485 68852
rect 375974 58853 376034 485147
rect 378731 479636 378797 479637
rect 378731 479572 378732 479636
rect 378796 479572 378797 479636
rect 378731 479571 378797 479572
rect 378179 476780 378245 476781
rect 378179 476716 378180 476780
rect 378244 476716 378245 476780
rect 378179 476715 378245 476716
rect 377259 472972 377325 472973
rect 377259 472908 377260 472972
rect 377324 472908 377325 472972
rect 377259 472907 377325 472908
rect 376707 374916 376773 374917
rect 376707 374852 376708 374916
rect 376772 374852 376773 374916
rect 376707 374851 376773 374852
rect 376710 364350 376770 374851
rect 376710 364290 376954 364350
rect 376894 273325 376954 364290
rect 376891 273324 376957 273325
rect 376891 273260 376892 273324
rect 376956 273260 376957 273324
rect 376891 273259 376957 273260
rect 377262 271421 377322 472907
rect 377443 471340 377509 471341
rect 377443 471276 377444 471340
rect 377508 471276 377509 471340
rect 377443 471275 377509 471276
rect 377446 382397 377506 471275
rect 377627 471204 377693 471205
rect 377627 471140 377628 471204
rect 377692 471140 377693 471204
rect 377627 471139 377693 471140
rect 377443 382396 377509 382397
rect 377443 382332 377444 382396
rect 377508 382332 377509 382396
rect 377443 382331 377509 382332
rect 377630 378861 377690 471139
rect 377811 468484 377877 468485
rect 377811 468420 377812 468484
rect 377876 468420 377877 468484
rect 377811 468419 377877 468420
rect 377627 378860 377693 378861
rect 377627 378796 377628 378860
rect 377692 378796 377693 378860
rect 377627 378795 377693 378796
rect 377814 378725 377874 468419
rect 377811 378724 377877 378725
rect 377811 378660 377812 378724
rect 377876 378660 377877 378724
rect 377811 378659 377877 378660
rect 377443 378180 377509 378181
rect 377443 378116 377444 378180
rect 377508 378116 377509 378180
rect 377443 378115 377509 378116
rect 377259 271420 377325 271421
rect 377259 271356 377260 271420
rect 377324 271356 377325 271420
rect 377259 271355 377325 271356
rect 377446 267613 377506 378115
rect 377995 357372 378061 357373
rect 377995 357308 377996 357372
rect 378060 357308 378061 357372
rect 377995 357307 378061 357308
rect 377811 273324 377877 273325
rect 377811 273260 377812 273324
rect 377876 273260 377877 273324
rect 377811 273259 377877 273260
rect 377814 273053 377874 273259
rect 377811 273052 377877 273053
rect 377811 272988 377812 273052
rect 377876 272988 377877 273052
rect 377811 272987 377877 272988
rect 377998 272645 378058 357307
rect 378182 273325 378242 476715
rect 378179 273324 378245 273325
rect 378179 273260 378180 273324
rect 378244 273260 378245 273324
rect 378179 273259 378245 273260
rect 377995 272644 378061 272645
rect 377995 272580 377996 272644
rect 378060 272580 378061 272644
rect 377995 272579 378061 272580
rect 376891 267612 376957 267613
rect 376891 267548 376892 267612
rect 376956 267548 376957 267612
rect 376891 267547 376957 267548
rect 377443 267612 377509 267613
rect 377443 267548 377444 267612
rect 377508 267548 377509 267612
rect 377443 267547 377509 267548
rect 376894 164117 376954 267547
rect 377995 252516 378061 252517
rect 377995 252452 377996 252516
rect 378060 252452 378061 252516
rect 377995 252451 378061 252452
rect 376891 164116 376957 164117
rect 376891 164052 376892 164116
rect 376956 164052 376957 164116
rect 376891 164051 376957 164052
rect 376894 162757 376954 164051
rect 376891 162756 376957 162757
rect 376891 162692 376892 162756
rect 376956 162692 376957 162756
rect 376891 162691 376957 162692
rect 377443 147796 377509 147797
rect 377443 147732 377444 147796
rect 377508 147732 377509 147796
rect 377443 147731 377509 147732
rect 375971 58852 376037 58853
rect 375971 58788 375972 58852
rect 376036 58788 376037 58852
rect 375971 58787 376037 58788
rect 374683 58716 374749 58717
rect 374683 58652 374684 58716
rect 374748 58652 374749 58716
rect 374683 58651 374749 58652
rect 374499 57764 374565 57765
rect 374499 57700 374500 57764
rect 374564 57700 374565 57764
rect 374499 57699 374565 57700
rect 377446 56405 377506 147731
rect 377998 146301 378058 252451
rect 377995 146300 378061 146301
rect 377995 146236 377996 146300
rect 378060 146236 378061 146300
rect 377995 146235 378061 146236
rect 377627 145892 377693 145893
rect 377627 145828 377628 145892
rect 377692 145828 377693 145892
rect 377627 145827 377693 145828
rect 377630 59397 377690 145827
rect 377811 145620 377877 145621
rect 377811 145556 377812 145620
rect 377876 145556 377877 145620
rect 377811 145555 377877 145556
rect 377627 59396 377693 59397
rect 377627 59332 377628 59396
rect 377692 59332 377693 59396
rect 377627 59331 377693 59332
rect 377443 56404 377509 56405
rect 377443 56340 377444 56404
rect 377508 56340 377509 56404
rect 377443 56339 377509 56340
rect 377814 56269 377874 145555
rect 378734 57085 378794 479571
rect 379467 478140 379533 478141
rect 379467 478076 379468 478140
rect 379532 478076 379533 478140
rect 379467 478075 379533 478076
rect 378915 474060 378981 474061
rect 378915 473996 378916 474060
rect 378980 473996 378981 474060
rect 378915 473995 378981 473996
rect 378918 57221 378978 473995
rect 379099 472564 379165 472565
rect 379099 472500 379100 472564
rect 379164 472500 379165 472564
rect 379099 472499 379165 472500
rect 379102 57493 379162 472499
rect 379470 470610 379530 478075
rect 379470 470550 379714 470610
rect 379654 165205 379714 470550
rect 379794 466308 380414 488898
rect 383514 493174 384134 527000
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 466308 384134 492618
rect 387234 496894 387854 527000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 466308 387854 496338
rect 390954 500614 391574 527000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 466308 391574 500058
rect 397794 507454 398414 527000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 466308 398414 470898
rect 401514 511174 402134 527000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 466308 402134 474618
rect 405234 514894 405854 527000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 466308 405854 478338
rect 408954 518614 409574 527000
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 466308 409574 482058
rect 415794 525454 416414 527000
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 466308 416414 488898
rect 419514 493174 420134 527000
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 466308 420134 492618
rect 423234 496894 423854 527000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 466308 423854 496338
rect 426954 500614 427574 527000
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 466308 427574 500058
rect 433794 507454 434414 527000
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 466308 434414 470898
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 466308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 466308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 466308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 466308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 637000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 637000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 637000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 637000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 637000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 637000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 637000 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 637000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 637000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 637000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 637000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 476067 634948 476133 634949
rect 476067 634884 476068 634948
rect 476132 634884 476133 634948
rect 476067 634883 476133 634884
rect 488579 634948 488645 634949
rect 488579 634884 488580 634948
rect 488644 634884 488645 634948
rect 488579 634883 488645 634884
rect 506611 634948 506677 634949
rect 506611 634884 506612 634948
rect 506676 634884 506677 634948
rect 506611 634883 506677 634884
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 466308 456134 492618
rect 459234 568894 459854 583000
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 466308 459854 496338
rect 462954 572614 463574 583000
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 466308 463574 500058
rect 469794 579454 470414 583000
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 466308 470414 470898
rect 473514 547174 474134 583000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 476070 489157 476130 634883
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 477234 550894 477854 583000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 476067 489156 476133 489157
rect 476067 489092 476068 489156
rect 476132 489092 476133 489156
rect 476067 489091 476133 489092
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 466308 474134 474618
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 466308 477854 478338
rect 480954 554614 481574 583000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 466308 481574 482058
rect 487794 561454 488414 583000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 466308 488414 488898
rect 488582 486437 488642 634883
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 491514 565174 492134 583000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 488579 486436 488645 486437
rect 488579 486372 488580 486436
rect 488644 486372 488645 486436
rect 488579 486371 488645 486372
rect 491514 466308 492134 492618
rect 495234 568894 495854 583000
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 466308 495854 496338
rect 498954 572614 499574 583000
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498515 466580 498581 466581
rect 498515 466516 498516 466580
rect 498580 466516 498581 466580
rect 498515 466515 498581 466516
rect 498518 464810 498578 466515
rect 498954 466308 499574 500058
rect 505794 579454 506414 583000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 506614 472837 506674 634883
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 509514 547174 510134 583000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 506611 472836 506677 472837
rect 506611 472772 506612 472836
rect 506676 472772 506677 472836
rect 506611 472771 506677 472772
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 466580 499869 466581
rect 499803 466516 499804 466580
rect 499868 466516 499869 466580
rect 499803 466515 499869 466516
rect 499806 464810 499866 466515
rect 505794 466308 506414 470898
rect 509514 466308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 466580 510909 466581
rect 510843 466516 510844 466580
rect 510908 466516 510909 466580
rect 510843 466515 510909 466516
rect 510846 464810 510906 466515
rect 513234 466308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 466308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 464750 498578 464810
rect 499688 464750 499866 464810
rect 510840 464750 510906 464810
rect 498464 464202 498524 464750
rect 499688 464202 499748 464750
rect 510840 464202 510900 464750
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 396056 380490 396116 381106
rect 397144 380490 397204 381106
rect 396030 380430 396116 380490
rect 397134 380430 397204 380490
rect 398232 380490 398292 381106
rect 399592 380490 399652 381106
rect 400544 380490 400604 381106
rect 401768 380490 401828 381106
rect 403128 380490 403188 381106
rect 404216 380490 404276 381106
rect 405440 380629 405500 381106
rect 405437 380628 405503 380629
rect 405437 380564 405438 380628
rect 405502 380564 405503 380628
rect 405437 380563 405503 380564
rect 406528 380490 406588 381106
rect 398232 380430 398298 380490
rect 396030 379405 396090 380430
rect 397134 379405 397194 380430
rect 396027 379404 396093 379405
rect 396027 379340 396028 379404
rect 396092 379340 396093 379404
rect 396027 379339 396093 379340
rect 397131 379404 397197 379405
rect 397131 379340 397132 379404
rect 397196 379340 397197 379404
rect 397131 379339 397197 379340
rect 398238 379269 398298 380430
rect 399526 380430 399652 380490
rect 400446 380430 400604 380490
rect 401734 380430 401828 380490
rect 403022 380430 403188 380490
rect 404126 380430 404276 380490
rect 406518 380430 406588 380490
rect 407616 380490 407676 381106
rect 408296 380490 408356 381106
rect 408704 380490 408764 381106
rect 410064 380490 410124 381106
rect 410744 380765 410804 381106
rect 410741 380764 410807 380765
rect 410741 380700 410742 380764
rect 410806 380700 410807 380764
rect 410741 380699 410807 380700
rect 407616 380430 407682 380490
rect 408296 380430 408418 380490
rect 408704 380430 408786 380490
rect 399526 379269 399586 380430
rect 400446 379269 400506 380430
rect 401734 379405 401794 380430
rect 401731 379404 401797 379405
rect 401731 379340 401732 379404
rect 401796 379340 401797 379404
rect 401731 379339 401797 379340
rect 403022 379269 403082 380430
rect 404126 380221 404186 380430
rect 404123 380220 404189 380221
rect 404123 380156 404124 380220
rect 404188 380156 404189 380220
rect 404123 380155 404189 380156
rect 406518 379405 406578 380430
rect 407622 379405 407682 380430
rect 408358 379405 408418 380430
rect 406515 379404 406581 379405
rect 406515 379340 406516 379404
rect 406580 379340 406581 379404
rect 406515 379339 406581 379340
rect 407619 379404 407685 379405
rect 407619 379340 407620 379404
rect 407684 379340 407685 379404
rect 407619 379339 407685 379340
rect 408355 379404 408421 379405
rect 408355 379340 408356 379404
rect 408420 379340 408421 379404
rect 408355 379339 408421 379340
rect 398235 379268 398301 379269
rect 398235 379204 398236 379268
rect 398300 379204 398301 379268
rect 398235 379203 398301 379204
rect 399523 379268 399589 379269
rect 399523 379204 399524 379268
rect 399588 379204 399589 379268
rect 399523 379203 399589 379204
rect 400443 379268 400509 379269
rect 400443 379204 400444 379268
rect 400508 379204 400509 379268
rect 400443 379203 400509 379204
rect 403019 379268 403085 379269
rect 403019 379204 403020 379268
rect 403084 379204 403085 379268
rect 403019 379203 403085 379204
rect 379794 364394 380414 379000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 359308 380414 363838
rect 383514 368114 384134 379000
rect 383514 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 384134 368114
rect 383514 367794 384134 367878
rect 383514 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 384134 367794
rect 383514 359308 384134 367558
rect 387234 369954 387854 379000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 359308 387854 369398
rect 390954 373674 391574 379000
rect 390954 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 391574 373674
rect 390954 373354 391574 373438
rect 390954 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 391574 373354
rect 390954 359308 391574 373118
rect 397794 363454 398414 379000
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 359308 398414 362898
rect 401514 367174 402134 379000
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 359308 402134 366618
rect 405234 370894 405854 379000
rect 408726 378181 408786 380430
rect 410014 380430 410124 380490
rect 411288 380490 411348 381106
rect 412376 380490 412436 381106
rect 413464 380629 413524 381106
rect 413461 380628 413527 380629
rect 413461 380564 413462 380628
rect 413526 380564 413527 380628
rect 413461 380563 413527 380564
rect 413600 380490 413660 381106
rect 411288 380430 411362 380490
rect 412376 380430 412466 380490
rect 410014 379269 410074 380430
rect 411302 379405 411362 380430
rect 412406 379405 412466 380430
rect 413510 380430 413660 380490
rect 414552 380490 414612 381106
rect 415912 380490 415972 381106
rect 414552 380430 414674 380490
rect 411299 379404 411365 379405
rect 411299 379340 411300 379404
rect 411364 379340 411365 379404
rect 411299 379339 411365 379340
rect 412403 379404 412469 379405
rect 412403 379340 412404 379404
rect 412468 379340 412469 379404
rect 412403 379339 412469 379340
rect 410011 379268 410077 379269
rect 410011 379204 410012 379268
rect 410076 379204 410077 379268
rect 410011 379203 410077 379204
rect 408723 378180 408789 378181
rect 408723 378116 408724 378180
rect 408788 378116 408789 378180
rect 408723 378115 408789 378116
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 359308 405854 370338
rect 408954 374614 409574 379000
rect 413510 378589 413570 380430
rect 414614 378589 414674 380430
rect 415902 380430 415972 380490
rect 416048 380490 416108 381106
rect 417000 380490 417060 381106
rect 418088 380490 418148 381106
rect 418496 380490 418556 381106
rect 419448 380629 419508 381106
rect 419445 380628 419511 380629
rect 419445 380564 419446 380628
rect 419510 380564 419511 380628
rect 419445 380563 419511 380564
rect 416048 380430 416146 380490
rect 417000 380430 417066 380490
rect 418088 380430 418170 380490
rect 415902 379269 415962 380430
rect 416086 379405 416146 380430
rect 416083 379404 416149 379405
rect 416083 379340 416084 379404
rect 416148 379340 416149 379404
rect 416083 379339 416149 379340
rect 417006 379269 417066 380430
rect 415899 379268 415965 379269
rect 415899 379204 415900 379268
rect 415964 379204 415965 379268
rect 415899 379203 415965 379204
rect 417003 379268 417069 379269
rect 417003 379204 417004 379268
rect 417068 379204 417069 379268
rect 417003 379203 417069 379204
rect 413507 378588 413573 378589
rect 413507 378524 413508 378588
rect 413572 378524 413573 378588
rect 413507 378523 413573 378524
rect 414611 378588 414677 378589
rect 414611 378524 414612 378588
rect 414676 378524 414677 378588
rect 414611 378523 414677 378524
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 359308 409574 374058
rect 415794 364394 416414 379000
rect 418110 378181 418170 380430
rect 418478 380430 418556 380490
rect 420672 380490 420732 381106
rect 421080 380765 421140 381106
rect 421077 380764 421143 380765
rect 421077 380700 421078 380764
rect 421142 380700 421143 380764
rect 421077 380699 421143 380700
rect 421760 380490 421820 381106
rect 422848 380490 422908 381106
rect 423528 380490 423588 381106
rect 420672 380430 420746 380490
rect 421760 380430 421850 380490
rect 422848 380430 422954 380490
rect 418478 378589 418538 380430
rect 418475 378588 418541 378589
rect 418475 378524 418476 378588
rect 418540 378524 418541 378588
rect 418475 378523 418541 378524
rect 418107 378180 418173 378181
rect 418107 378116 418108 378180
rect 418172 378116 418173 378180
rect 418107 378115 418173 378116
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 359308 416414 363838
rect 419514 368114 420134 379000
rect 420686 378181 420746 380430
rect 421790 378181 421850 380430
rect 422894 378181 422954 380430
rect 423446 380430 423588 380490
rect 423936 380490 423996 381106
rect 425296 380490 425356 381106
rect 423936 380430 424058 380490
rect 423446 379269 423506 380430
rect 423443 379268 423509 379269
rect 423443 379204 423444 379268
rect 423508 379204 423509 379268
rect 423443 379203 423509 379204
rect 420683 378180 420749 378181
rect 420683 378116 420684 378180
rect 420748 378116 420749 378180
rect 420683 378115 420749 378116
rect 421787 378180 421853 378181
rect 421787 378116 421788 378180
rect 421852 378116 421853 378180
rect 421787 378115 421853 378116
rect 422891 378180 422957 378181
rect 422891 378116 422892 378180
rect 422956 378116 422957 378180
rect 422891 378115 422957 378116
rect 419514 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 420134 368114
rect 419514 367794 420134 367878
rect 419514 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 420134 367794
rect 419514 359308 420134 367558
rect 423234 369954 423854 379000
rect 423998 378181 424058 380430
rect 425286 380430 425356 380490
rect 425976 380490 426036 381106
rect 426384 380493 426444 381106
rect 426384 380492 426453 380493
rect 425976 380430 426082 380490
rect 426384 380430 426388 380492
rect 425286 378181 425346 380430
rect 426022 379405 426082 380430
rect 426387 380428 426388 380430
rect 426452 380428 426453 380492
rect 427608 380490 427668 381106
rect 428288 380901 428348 381106
rect 428285 380900 428351 380901
rect 428285 380836 428286 380900
rect 428350 380836 428351 380900
rect 428285 380835 428351 380836
rect 428696 380490 428756 381106
rect 429784 380490 429844 381106
rect 431008 380490 431068 381106
rect 431144 380901 431204 381106
rect 431141 380900 431207 380901
rect 431141 380836 431142 380900
rect 431206 380836 431207 380900
rect 431141 380835 431207 380836
rect 427608 380430 427738 380490
rect 426387 380427 426453 380428
rect 426019 379404 426085 379405
rect 426019 379340 426020 379404
rect 426084 379340 426085 379404
rect 426019 379339 426085 379340
rect 423995 378180 424061 378181
rect 423995 378116 423996 378180
rect 424060 378116 424061 378180
rect 423995 378115 424061 378116
rect 425283 378180 425349 378181
rect 425283 378116 425284 378180
rect 425348 378116 425349 378180
rect 425283 378115 425349 378116
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 359308 423854 369398
rect 426954 373674 427574 379000
rect 427678 378861 427738 380430
rect 428598 380430 428756 380490
rect 429702 380430 429844 380490
rect 430990 380430 431068 380490
rect 432232 380490 432292 381106
rect 433320 380490 433380 381106
rect 433592 380901 433652 381106
rect 433589 380900 433655 380901
rect 433589 380836 433590 380900
rect 433654 380836 433655 380900
rect 433589 380835 433655 380836
rect 434408 380629 434468 381106
rect 434405 380628 434471 380629
rect 434405 380564 434406 380628
rect 434470 380564 434471 380628
rect 434405 380563 434471 380564
rect 435768 380490 435828 381106
rect 436040 380765 436100 381106
rect 436037 380764 436103 380765
rect 436037 380700 436038 380764
rect 436102 380700 436103 380764
rect 436037 380699 436103 380700
rect 436992 380490 437052 381106
rect 438080 380490 438140 381106
rect 438488 380901 438548 381106
rect 438485 380900 438551 380901
rect 438485 380836 438486 380900
rect 438550 380836 438551 380900
rect 438485 380835 438551 380836
rect 439168 380490 439228 381106
rect 440936 380765 440996 381106
rect 443520 380765 443580 381106
rect 440933 380764 440999 380765
rect 440933 380700 440934 380764
rect 440998 380700 440999 380764
rect 440933 380699 440999 380700
rect 443517 380764 443583 380765
rect 443517 380700 443518 380764
rect 443582 380700 443583 380764
rect 443517 380699 443583 380700
rect 445968 380490 446028 381106
rect 432232 380430 432338 380490
rect 433320 380430 433442 380490
rect 435768 380430 435834 380490
rect 427675 378860 427741 378861
rect 427675 378796 427676 378860
rect 427740 378796 427741 378860
rect 427675 378795 427741 378796
rect 428598 378181 428658 380430
rect 429702 378181 429762 380430
rect 430990 378861 431050 380430
rect 430987 378860 431053 378861
rect 430987 378796 430988 378860
rect 431052 378796 431053 378860
rect 430987 378795 431053 378796
rect 432278 378317 432338 380430
rect 433382 378725 433442 380430
rect 435774 379405 435834 380430
rect 436878 380430 437052 380490
rect 437982 380430 438140 380490
rect 439086 380430 439228 380490
rect 445894 380430 446028 380490
rect 448280 380490 448340 381106
rect 451000 380490 451060 381106
rect 453448 380490 453508 381106
rect 455896 380490 455956 381106
rect 458480 380490 458540 381106
rect 448280 380430 448346 380490
rect 451000 380430 451106 380490
rect 435771 379404 435837 379405
rect 435771 379340 435772 379404
rect 435836 379340 435837 379404
rect 435771 379339 435837 379340
rect 433379 378724 433445 378725
rect 433379 378660 433380 378724
rect 433444 378660 433445 378724
rect 433379 378659 433445 378660
rect 432275 378316 432341 378317
rect 432275 378252 432276 378316
rect 432340 378252 432341 378316
rect 432275 378251 432341 378252
rect 428595 378180 428661 378181
rect 428595 378116 428596 378180
rect 428660 378116 428661 378180
rect 428595 378115 428661 378116
rect 429699 378180 429765 378181
rect 429699 378116 429700 378180
rect 429764 378116 429765 378180
rect 429699 378115 429765 378116
rect 426954 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 427574 373674
rect 426954 373354 427574 373438
rect 426954 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 427574 373354
rect 426954 359308 427574 373118
rect 433794 363454 434414 379000
rect 436878 378725 436938 380430
rect 437982 379405 438042 380430
rect 437979 379404 438045 379405
rect 437979 379340 437980 379404
rect 438044 379340 438045 379404
rect 437979 379339 438045 379340
rect 436875 378724 436941 378725
rect 436875 378660 436876 378724
rect 436940 378660 436941 378724
rect 436875 378659 436941 378660
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 359308 434414 362898
rect 437514 367174 438134 379000
rect 439086 378181 439146 380430
rect 445894 379405 445954 380430
rect 448286 379405 448346 380430
rect 451046 379405 451106 380430
rect 453438 380430 453508 380490
rect 455830 380430 455956 380490
rect 458406 380430 458540 380490
rect 460928 380490 460988 381106
rect 463512 380490 463572 381106
rect 465960 380490 466020 381106
rect 468544 380490 468604 381106
rect 470992 380490 471052 381106
rect 460928 380430 461042 380490
rect 463512 380430 463618 380490
rect 453438 379405 453498 380430
rect 455830 379405 455890 380430
rect 458406 379405 458466 380430
rect 460982 379405 461042 380430
rect 445891 379404 445957 379405
rect 445891 379340 445892 379404
rect 445956 379340 445957 379404
rect 445891 379339 445957 379340
rect 448283 379404 448349 379405
rect 448283 379340 448284 379404
rect 448348 379340 448349 379404
rect 448283 379339 448349 379340
rect 451043 379404 451109 379405
rect 451043 379340 451044 379404
rect 451108 379340 451109 379404
rect 451043 379339 451109 379340
rect 453435 379404 453501 379405
rect 453435 379340 453436 379404
rect 453500 379340 453501 379404
rect 453435 379339 453501 379340
rect 455827 379404 455893 379405
rect 455827 379340 455828 379404
rect 455892 379340 455893 379404
rect 455827 379339 455893 379340
rect 458403 379404 458469 379405
rect 458403 379340 458404 379404
rect 458468 379340 458469 379404
rect 458403 379339 458469 379340
rect 460979 379404 461045 379405
rect 460979 379340 460980 379404
rect 461044 379340 461045 379404
rect 460979 379339 461045 379340
rect 463558 379269 463618 380430
rect 465950 380430 466020 380490
rect 468526 380430 468604 380490
rect 470918 380430 471052 380490
rect 473440 380490 473500 381106
rect 475888 380490 475948 381106
rect 478472 380490 478532 381106
rect 480920 380490 480980 381106
rect 473440 380430 473554 380490
rect 463555 379268 463621 379269
rect 463555 379204 463556 379268
rect 463620 379204 463621 379268
rect 463555 379203 463621 379204
rect 439083 378180 439149 378181
rect 439083 378116 439084 378180
rect 439148 378116 439149 378180
rect 439083 378115 439149 378116
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 359308 438134 366618
rect 441234 370894 441854 379000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 359308 441854 370338
rect 444954 374614 445574 379000
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 359308 445574 374058
rect 451794 364394 452414 379000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 359308 452414 363838
rect 455514 368114 456134 379000
rect 455514 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 456134 368114
rect 455514 367794 456134 367878
rect 455514 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 456134 367794
rect 455514 359308 456134 367558
rect 459234 369954 459854 379000
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 359308 459854 369398
rect 462954 373674 463574 379000
rect 465950 378997 466010 380430
rect 465947 378996 466013 378997
rect 465947 378932 465948 378996
rect 466012 378932 466013 378996
rect 465947 378931 466013 378932
rect 468526 378725 468586 380430
rect 468523 378724 468589 378725
rect 468523 378660 468524 378724
rect 468588 378660 468589 378724
rect 468523 378659 468589 378660
rect 462954 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 463574 373674
rect 462954 373354 463574 373438
rect 462954 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 463574 373354
rect 462954 359308 463574 373118
rect 469794 363454 470414 379000
rect 470918 378861 470978 380430
rect 473494 379269 473554 380430
rect 475886 380430 475948 380490
rect 478462 380430 478532 380490
rect 480670 380430 480980 380490
rect 483368 380490 483428 381106
rect 485952 380629 486012 381106
rect 485949 380628 486015 380629
rect 485949 380564 485950 380628
rect 486014 380564 486015 380628
rect 485949 380563 486015 380564
rect 503224 380490 503284 381106
rect 483368 380430 483490 380490
rect 475886 379405 475946 380430
rect 475883 379404 475949 379405
rect 475883 379340 475884 379404
rect 475948 379340 475949 379404
rect 475883 379339 475949 379340
rect 473491 379268 473557 379269
rect 473491 379204 473492 379268
rect 473556 379204 473557 379268
rect 473491 379203 473557 379204
rect 470915 378860 470981 378861
rect 470915 378796 470916 378860
rect 470980 378796 470981 378860
rect 470915 378795 470981 378796
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 359308 470414 362898
rect 473514 367174 474134 379000
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 359308 474134 366618
rect 477234 370894 477854 379000
rect 478462 378997 478522 380430
rect 478459 378996 478525 378997
rect 478459 378932 478460 378996
rect 478524 378932 478525 378996
rect 478459 378931 478525 378932
rect 480670 378181 480730 380430
rect 480667 378180 480733 378181
rect 480667 378116 480668 378180
rect 480732 378116 480733 378180
rect 480667 378115 480733 378116
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 359308 477854 370338
rect 480954 374614 481574 379000
rect 483430 378861 483490 380430
rect 503118 380430 503284 380490
rect 503360 380490 503420 381106
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 503360 380430 503546 380490
rect 503118 379269 503178 380430
rect 503486 379269 503546 380430
rect 503115 379268 503181 379269
rect 503115 379204 503116 379268
rect 503180 379204 503181 379268
rect 503115 379203 503181 379204
rect 503483 379268 503549 379269
rect 503483 379204 503484 379268
rect 503548 379204 503549 379268
rect 503483 379203 503549 379204
rect 483427 378860 483493 378861
rect 483427 378796 483428 378860
rect 483492 378796 483493 378860
rect 483427 378795 483493 378796
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 359308 481574 374058
rect 487794 364394 488414 379000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 359308 488414 363838
rect 491514 368114 492134 379000
rect 491514 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 491514 367794 492134 367878
rect 491514 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 491514 359308 492134 367558
rect 495234 369954 495854 379000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 359308 495854 369398
rect 498954 373674 499574 379000
rect 498954 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 498954 373354 499574 373438
rect 498954 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 498954 359308 499574 373118
rect 505794 363454 506414 379000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 359308 506414 362898
rect 509514 367174 510134 379000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 359308 510134 366618
rect 513234 370894 513854 379000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 359308 513854 370338
rect 516954 374614 517574 379000
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 359308 517574 374058
rect 498515 358868 498581 358869
rect 498515 358804 498516 358868
rect 498580 358804 498581 358868
rect 498515 358803 498581 358804
rect 499803 358868 499869 358869
rect 499803 358804 499804 358868
rect 499868 358804 499869 358868
rect 499803 358803 499869 358804
rect 510843 358868 510909 358869
rect 510843 358804 510844 358868
rect 510908 358804 510909 358868
rect 510843 358803 510909 358804
rect 498518 358050 498578 358803
rect 499806 358050 499866 358803
rect 510846 358050 510906 358803
rect 498464 357990 498578 358050
rect 499688 357990 499866 358050
rect 510840 357990 510906 358050
rect 498464 357202 498524 357990
rect 499688 357202 499748 357990
rect 510840 357202 510900 357990
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 396056 273730 396116 274040
rect 397144 273730 397204 274040
rect 398232 273730 398292 274040
rect 399592 273730 399652 274040
rect 400544 273730 400604 274040
rect 401768 273730 401828 274040
rect 403128 273730 403188 274040
rect 404216 273730 404276 274040
rect 405440 273730 405500 274040
rect 406528 273730 406588 274040
rect 396030 273670 396116 273730
rect 397134 273670 397204 273730
rect 397502 273670 398292 273730
rect 399526 273670 399652 273730
rect 400446 273670 400604 273730
rect 401734 273670 401828 273730
rect 403022 273670 403188 273730
rect 404126 273670 404276 273730
rect 405046 273670 405500 273730
rect 406518 273670 406588 273730
rect 407616 273730 407676 274040
rect 408296 273730 408356 274040
rect 407616 273670 407682 273730
rect 379794 256394 380414 272000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 252308 380414 255838
rect 383514 260114 384134 272000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 252308 384134 259558
rect 387234 261954 387854 272000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 252308 387854 261398
rect 390954 265674 391574 272000
rect 396030 271285 396090 273670
rect 396027 271284 396093 271285
rect 396027 271220 396028 271284
rect 396092 271220 396093 271284
rect 396027 271219 396093 271220
rect 397134 271149 397194 273670
rect 397131 271148 397197 271149
rect 397131 271084 397132 271148
rect 397196 271084 397197 271148
rect 397131 271083 397197 271084
rect 397502 270605 397562 273670
rect 397499 270604 397565 270605
rect 397499 270540 397500 270604
rect 397564 270540 397565 270604
rect 397499 270539 397565 270540
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 252308 391574 265118
rect 397794 255454 398414 272000
rect 399526 270605 399586 273670
rect 400446 270605 400506 273670
rect 401734 272237 401794 273670
rect 401731 272236 401797 272237
rect 401731 272172 401732 272236
rect 401796 272172 401797 272236
rect 401731 272171 401797 272172
rect 399523 270604 399589 270605
rect 399523 270540 399524 270604
rect 399588 270540 399589 270604
rect 399523 270539 399589 270540
rect 400443 270604 400509 270605
rect 400443 270540 400444 270604
rect 400508 270540 400509 270604
rect 400443 270539 400509 270540
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252308 398414 254898
rect 401514 259174 402134 272000
rect 403022 270605 403082 273670
rect 404126 270605 404186 273670
rect 405046 270605 405106 273670
rect 403019 270604 403085 270605
rect 403019 270540 403020 270604
rect 403084 270540 403085 270604
rect 403019 270539 403085 270540
rect 404123 270604 404189 270605
rect 404123 270540 404124 270604
rect 404188 270540 404189 270604
rect 404123 270539 404189 270540
rect 405043 270604 405109 270605
rect 405043 270540 405044 270604
rect 405108 270540 405109 270604
rect 405043 270539 405109 270540
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252308 402134 258618
rect 405234 262894 405854 272000
rect 406518 270877 406578 273670
rect 406515 270876 406581 270877
rect 406515 270812 406516 270876
rect 406580 270812 406581 270876
rect 406515 270811 406581 270812
rect 407622 270605 407682 273670
rect 408174 273670 408356 273730
rect 408704 273730 408764 274040
rect 410064 273730 410124 274040
rect 408704 273670 408786 273730
rect 408174 271421 408234 273670
rect 408171 271420 408237 271421
rect 408171 271356 408172 271420
rect 408236 271356 408237 271420
rect 408171 271355 408237 271356
rect 408726 270605 408786 273670
rect 410014 273670 410124 273730
rect 410744 273730 410804 274040
rect 411288 273730 411348 274040
rect 412376 273730 412436 274040
rect 413464 273730 413524 274040
rect 410744 273670 410810 273730
rect 411288 273670 411362 273730
rect 412376 273670 412466 273730
rect 407619 270604 407685 270605
rect 407619 270540 407620 270604
rect 407684 270540 407685 270604
rect 407619 270539 407685 270540
rect 408723 270604 408789 270605
rect 408723 270540 408724 270604
rect 408788 270540 408789 270604
rect 408723 270539 408789 270540
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252308 405854 262338
rect 408954 266614 409574 272000
rect 410014 270605 410074 273670
rect 410750 271149 410810 273670
rect 410747 271148 410813 271149
rect 410747 271084 410748 271148
rect 410812 271084 410813 271148
rect 410747 271083 410813 271084
rect 411302 270741 411362 273670
rect 411299 270740 411365 270741
rect 411299 270676 411300 270740
rect 411364 270676 411365 270740
rect 411299 270675 411365 270676
rect 412406 270605 412466 273670
rect 413326 273670 413524 273730
rect 413600 273730 413660 274040
rect 414552 273730 414612 274040
rect 415912 273730 415972 274040
rect 413600 273670 413754 273730
rect 413326 270605 413386 273670
rect 413694 271149 413754 273670
rect 414430 273670 414612 273730
rect 415902 273670 415972 273730
rect 416048 273730 416108 274040
rect 417000 273730 417060 274040
rect 418088 273730 418148 274040
rect 418496 273730 418556 274040
rect 419448 273730 419508 274040
rect 416048 273670 416146 273730
rect 417000 273670 417066 273730
rect 418088 273670 418170 273730
rect 413691 271148 413757 271149
rect 413691 271084 413692 271148
rect 413756 271084 413757 271148
rect 413691 271083 413757 271084
rect 414430 270605 414490 273670
rect 415902 272237 415962 273670
rect 416086 272237 416146 273670
rect 415899 272236 415965 272237
rect 415899 272172 415900 272236
rect 415964 272172 415965 272236
rect 415899 272171 415965 272172
rect 416083 272236 416149 272237
rect 416083 272172 416084 272236
rect 416148 272172 416149 272236
rect 416083 272171 416149 272172
rect 410011 270604 410077 270605
rect 410011 270540 410012 270604
rect 410076 270540 410077 270604
rect 410011 270539 410077 270540
rect 412403 270604 412469 270605
rect 412403 270540 412404 270604
rect 412468 270540 412469 270604
rect 412403 270539 412469 270540
rect 413323 270604 413389 270605
rect 413323 270540 413324 270604
rect 413388 270540 413389 270604
rect 413323 270539 413389 270540
rect 414427 270604 414493 270605
rect 414427 270540 414428 270604
rect 414492 270540 414493 270604
rect 414427 270539 414493 270540
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252308 409574 266058
rect 415794 256394 416414 272000
rect 417006 270605 417066 273670
rect 418110 270605 418170 273670
rect 418478 273670 418556 273730
rect 419214 273670 419508 273730
rect 420672 273730 420732 274040
rect 420672 273670 420746 273730
rect 418478 271149 418538 273670
rect 418475 271148 418541 271149
rect 418475 271084 418476 271148
rect 418540 271084 418541 271148
rect 418475 271083 418541 271084
rect 417003 270604 417069 270605
rect 417003 270540 417004 270604
rect 417068 270540 417069 270604
rect 417003 270539 417069 270540
rect 418107 270604 418173 270605
rect 418107 270540 418108 270604
rect 418172 270540 418173 270604
rect 418107 270539 418173 270540
rect 419214 269925 419274 273670
rect 419211 269924 419277 269925
rect 419211 269860 419212 269924
rect 419276 269860 419277 269924
rect 419211 269859 419277 269860
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 252308 416414 255838
rect 419514 260114 420134 272000
rect 420686 270605 420746 273670
rect 421080 273597 421140 274040
rect 421760 273730 421820 274040
rect 422848 273730 422908 274040
rect 423528 273730 423588 274040
rect 423936 273730 423996 274040
rect 425296 273730 425356 274040
rect 421760 273670 421850 273730
rect 422848 273670 422954 273730
rect 421077 273596 421143 273597
rect 421077 273532 421078 273596
rect 421142 273532 421143 273596
rect 421077 273531 421143 273532
rect 421790 270605 421850 273670
rect 422894 273189 422954 273670
rect 423446 273670 423588 273730
rect 423814 273670 423996 273730
rect 425286 273670 425356 273730
rect 425976 273730 426036 274040
rect 426384 273869 426444 274040
rect 426381 273868 426447 273869
rect 426381 273804 426382 273868
rect 426446 273804 426447 273868
rect 426381 273803 426447 273804
rect 427608 273730 427668 274040
rect 428288 273730 428348 274040
rect 428696 273730 428756 274040
rect 429784 273730 429844 274040
rect 431008 273730 431068 274040
rect 425976 273670 426082 273730
rect 427608 273670 427738 273730
rect 423446 273189 423506 273670
rect 422891 273188 422957 273189
rect 422891 273124 422892 273188
rect 422956 273124 422957 273188
rect 422891 273123 422957 273124
rect 423443 273188 423509 273189
rect 423443 273124 423444 273188
rect 423508 273124 423509 273188
rect 423443 273123 423509 273124
rect 423814 272509 423874 273670
rect 425286 273053 425346 273670
rect 426022 273189 426082 273670
rect 426019 273188 426085 273189
rect 426019 273124 426020 273188
rect 426084 273124 426085 273188
rect 426019 273123 426085 273124
rect 425283 273052 425349 273053
rect 425283 272988 425284 273052
rect 425348 272988 425349 273052
rect 425283 272987 425349 272988
rect 423811 272508 423877 272509
rect 423811 272444 423812 272508
rect 423876 272444 423877 272508
rect 423811 272443 423877 272444
rect 420683 270604 420749 270605
rect 420683 270540 420684 270604
rect 420748 270540 420749 270604
rect 420683 270539 420749 270540
rect 421787 270604 421853 270605
rect 421787 270540 421788 270604
rect 421852 270540 421853 270604
rect 421787 270539 421853 270540
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 252308 420134 259558
rect 423234 261954 423854 272000
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 252308 423854 261398
rect 426954 265674 427574 272000
rect 427678 269789 427738 273670
rect 428230 273670 428348 273730
rect 428598 273670 428756 273730
rect 429702 273670 429844 273730
rect 430990 273670 431068 273730
rect 428230 272917 428290 273670
rect 428227 272916 428293 272917
rect 428227 272852 428228 272916
rect 428292 272852 428293 272916
rect 428227 272851 428293 272852
rect 428598 271829 428658 273670
rect 428595 271828 428661 271829
rect 428595 271764 428596 271828
rect 428660 271764 428661 271828
rect 428595 271763 428661 271764
rect 429702 270741 429762 273670
rect 430990 273461 431050 273670
rect 431144 273597 431204 274040
rect 432232 273730 432292 274040
rect 432232 273670 432338 273730
rect 431141 273596 431207 273597
rect 431141 273532 431142 273596
rect 431206 273532 431207 273596
rect 431141 273531 431207 273532
rect 430987 273460 431053 273461
rect 430987 273396 430988 273460
rect 431052 273396 431053 273460
rect 430987 273395 431053 273396
rect 432278 270877 432338 273670
rect 433320 273597 433380 274040
rect 433592 273730 433652 274040
rect 433566 273670 433652 273730
rect 434408 273730 434468 274040
rect 435768 273730 435828 274040
rect 436040 273730 436100 274040
rect 436992 273730 437052 274040
rect 434408 273670 434730 273730
rect 435768 273670 435834 273730
rect 433317 273596 433383 273597
rect 433317 273532 433318 273596
rect 433382 273532 433383 273596
rect 433317 273531 433383 273532
rect 433566 271829 433626 273670
rect 433563 271828 433629 271829
rect 433563 271764 433564 271828
rect 433628 271764 433629 271828
rect 433563 271763 433629 271764
rect 432275 270876 432341 270877
rect 432275 270812 432276 270876
rect 432340 270812 432341 270876
rect 432275 270811 432341 270812
rect 429699 270740 429765 270741
rect 429699 270676 429700 270740
rect 429764 270676 429765 270740
rect 429699 270675 429765 270676
rect 427675 269788 427741 269789
rect 427675 269724 427676 269788
rect 427740 269724 427741 269788
rect 427675 269723 427741 269724
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 252308 427574 265118
rect 433794 255454 434414 272000
rect 434670 270877 434730 273670
rect 434667 270876 434733 270877
rect 434667 270812 434668 270876
rect 434732 270812 434733 270876
rect 434667 270811 434733 270812
rect 435774 270469 435834 273670
rect 435958 273670 436100 273730
rect 436878 273670 437052 273730
rect 438080 273730 438140 274040
rect 438488 273730 438548 274040
rect 439168 273730 439228 274040
rect 440936 273730 440996 274040
rect 443520 273730 443580 274040
rect 445968 273730 446028 274040
rect 438080 273670 438410 273730
rect 438488 273670 438594 273730
rect 435958 271285 436018 273670
rect 436878 271829 436938 273670
rect 436875 271828 436941 271829
rect 436875 271764 436876 271828
rect 436940 271764 436941 271828
rect 436875 271763 436941 271764
rect 435955 271284 436021 271285
rect 435955 271220 435956 271284
rect 436020 271220 436021 271284
rect 435955 271219 436021 271220
rect 435771 270468 435837 270469
rect 435771 270404 435772 270468
rect 435836 270404 435837 270468
rect 435771 270403 435837 270404
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 252308 434414 254898
rect 437514 259174 438134 272000
rect 438350 270877 438410 273670
rect 438534 271829 438594 273670
rect 439086 273670 439228 273730
rect 440926 273670 440996 273730
rect 443502 273670 443580 273730
rect 445894 273670 446028 273730
rect 448280 273730 448340 274040
rect 451000 273730 451060 274040
rect 448280 273670 448346 273730
rect 451000 273670 451106 273730
rect 438531 271828 438597 271829
rect 438531 271764 438532 271828
rect 438596 271764 438597 271828
rect 438531 271763 438597 271764
rect 439086 270877 439146 273670
rect 440926 271421 440986 273670
rect 440923 271420 440989 271421
rect 440923 271356 440924 271420
rect 440988 271356 440989 271420
rect 440923 271355 440989 271356
rect 438347 270876 438413 270877
rect 438347 270812 438348 270876
rect 438412 270812 438413 270876
rect 438347 270811 438413 270812
rect 439083 270876 439149 270877
rect 439083 270812 439084 270876
rect 439148 270812 439149 270876
rect 439083 270811 439149 270812
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 252308 438134 258618
rect 441234 262894 441854 272000
rect 443502 271829 443562 273670
rect 443499 271828 443565 271829
rect 443499 271764 443500 271828
rect 443564 271764 443565 271828
rect 443499 271763 443565 271764
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 252308 441854 262338
rect 444954 266614 445574 272000
rect 445894 271829 445954 273670
rect 448286 271829 448346 273670
rect 451046 271829 451106 273670
rect 453448 273597 453508 274040
rect 455896 273730 455956 274040
rect 458480 273730 458540 274040
rect 455830 273670 455956 273730
rect 458406 273670 458540 273730
rect 460928 273730 460988 274040
rect 463512 273730 463572 274040
rect 465960 273730 466020 274040
rect 468544 273730 468604 274040
rect 470992 273730 471052 274040
rect 460928 273670 461042 273730
rect 453445 273596 453511 273597
rect 453445 273532 453446 273596
rect 453510 273532 453511 273596
rect 453445 273531 453511 273532
rect 455830 272237 455890 273670
rect 455827 272236 455893 272237
rect 455827 272172 455828 272236
rect 455892 272172 455893 272236
rect 455827 272171 455893 272172
rect 445891 271828 445957 271829
rect 445891 271764 445892 271828
rect 445956 271764 445957 271828
rect 445891 271763 445957 271764
rect 448283 271828 448349 271829
rect 448283 271764 448284 271828
rect 448348 271764 448349 271828
rect 448283 271763 448349 271764
rect 451043 271828 451109 271829
rect 451043 271764 451044 271828
rect 451108 271764 451109 271828
rect 451043 271763 451109 271764
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 252308 445574 266058
rect 451794 256394 452414 272000
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 252308 452414 255838
rect 455514 260114 456134 272000
rect 458406 271829 458466 273670
rect 458403 271828 458469 271829
rect 458403 271764 458404 271828
rect 458468 271764 458469 271828
rect 458403 271763 458469 271764
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 252308 456134 259558
rect 459234 261954 459854 272000
rect 460982 271557 461042 273670
rect 462638 273670 463572 273730
rect 465950 273670 466020 273730
rect 468526 273670 468604 273730
rect 470918 273670 471052 273730
rect 473440 273730 473500 274040
rect 475888 273730 475948 274040
rect 478472 273730 478532 274040
rect 480920 273730 480980 274040
rect 483368 273730 483428 274040
rect 473440 273670 473554 273730
rect 460979 271556 461045 271557
rect 460979 271492 460980 271556
rect 461044 271492 461045 271556
rect 460979 271491 461045 271492
rect 462638 271013 462698 273670
rect 462635 271012 462701 271013
rect 462635 270948 462636 271012
rect 462700 270948 462701 271012
rect 462635 270947 462701 270948
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 252308 459854 261398
rect 462954 265674 463574 272000
rect 465950 271693 466010 273670
rect 468526 273053 468586 273670
rect 470918 273053 470978 273670
rect 468523 273052 468589 273053
rect 468523 272988 468524 273052
rect 468588 272988 468589 273052
rect 468523 272987 468589 272988
rect 470915 273052 470981 273053
rect 470915 272988 470916 273052
rect 470980 272988 470981 273052
rect 470915 272987 470981 272988
rect 473494 272917 473554 273670
rect 475886 273670 475948 273730
rect 478462 273670 478532 273730
rect 480854 273670 480980 273730
rect 483246 273670 483428 273730
rect 485952 273730 486012 274040
rect 503224 273730 503284 274040
rect 485952 273670 486066 273730
rect 475886 272917 475946 273670
rect 473491 272916 473557 272917
rect 473491 272852 473492 272916
rect 473556 272852 473557 272916
rect 473491 272851 473557 272852
rect 475883 272916 475949 272917
rect 475883 272852 475884 272916
rect 475948 272852 475949 272916
rect 475883 272851 475949 272852
rect 478462 272781 478522 273670
rect 480854 272781 480914 273670
rect 478459 272780 478525 272781
rect 478459 272716 478460 272780
rect 478524 272716 478525 272780
rect 478459 272715 478525 272716
rect 480851 272780 480917 272781
rect 480851 272716 480852 272780
rect 480916 272716 480917 272780
rect 480851 272715 480917 272716
rect 483246 272645 483306 273670
rect 486006 272645 486066 273670
rect 503118 273670 503284 273730
rect 503360 273730 503420 274040
rect 503360 273670 503546 273730
rect 483243 272644 483309 272645
rect 483243 272580 483244 272644
rect 483308 272580 483309 272644
rect 483243 272579 483309 272580
rect 486003 272644 486069 272645
rect 486003 272580 486004 272644
rect 486068 272580 486069 272644
rect 486003 272579 486069 272580
rect 465947 271692 466013 271693
rect 465947 271628 465948 271692
rect 466012 271628 466013 271692
rect 465947 271627 466013 271628
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 252308 463574 265118
rect 469794 255454 470414 272000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 252308 470414 254898
rect 473514 259174 474134 272000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 252308 474134 258618
rect 477234 262894 477854 272000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 252308 477854 262338
rect 480954 266614 481574 272000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 252308 481574 266058
rect 487794 256394 488414 272000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 252308 488414 255838
rect 491514 260114 492134 272000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 252308 492134 259558
rect 495234 261954 495854 272000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 252308 495854 261398
rect 498954 265674 499574 272000
rect 503118 271693 503178 273670
rect 503115 271692 503181 271693
rect 503115 271628 503116 271692
rect 503180 271628 503181 271692
rect 503115 271627 503181 271628
rect 503486 271285 503546 273670
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 503483 271284 503549 271285
rect 503483 271220 503484 271284
rect 503548 271220 503549 271284
rect 503483 271219 503549 271220
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498515 252788 498581 252789
rect 498515 252724 498516 252788
rect 498580 252724 498581 252788
rect 498515 252723 498581 252724
rect 498518 250610 498578 252723
rect 498954 252308 499574 265118
rect 505794 255454 506414 272000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 499803 253332 499869 253333
rect 499803 253268 499804 253332
rect 499868 253268 499869 253332
rect 499803 253267 499869 253268
rect 499806 250610 499866 253267
rect 505794 252308 506414 254898
rect 509514 259174 510134 272000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 252308 510134 258618
rect 513234 262894 513854 272000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 510843 252652 510909 252653
rect 510843 252588 510844 252652
rect 510908 252588 510909 252652
rect 510843 252587 510909 252588
rect 510846 250610 510906 252587
rect 513234 252308 513854 262338
rect 516954 266614 517574 272000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 252308 517574 266058
rect 498464 250550 498578 250610
rect 499688 250550 499866 250610
rect 510840 250550 510906 250610
rect 498464 250240 498524 250550
rect 499688 250240 499748 250550
rect 510840 250240 510900 250550
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 396056 167010 396116 167106
rect 397144 167010 397204 167106
rect 396030 166950 396116 167010
rect 397134 166950 397204 167010
rect 398232 167010 398292 167106
rect 399592 167010 399652 167106
rect 400544 167010 400604 167106
rect 401768 167010 401828 167106
rect 403128 167010 403188 167106
rect 404216 167010 404276 167106
rect 405440 167010 405500 167106
rect 406528 167010 406588 167106
rect 398232 166950 398298 167010
rect 379651 165204 379717 165205
rect 379651 165140 379652 165204
rect 379716 165140 379717 165204
rect 379651 165139 379717 165140
rect 379794 148394 380414 165000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379794 145308 380414 147838
rect 383514 152114 384134 165000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 155834 387854 165000
rect 387234 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 387854 155834
rect 387234 155514 387854 155598
rect 387234 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 387854 155514
rect 387234 145308 387854 155278
rect 390954 157674 391574 165000
rect 396030 164253 396090 166950
rect 397134 164389 397194 166950
rect 398238 165613 398298 166950
rect 399526 166950 399652 167010
rect 400446 166950 400604 167010
rect 401734 166950 401828 167010
rect 403022 166950 403188 167010
rect 404126 166950 404276 167010
rect 405414 166950 405500 167010
rect 406518 166950 406588 167010
rect 407616 167010 407676 167106
rect 408296 167010 408356 167106
rect 407616 166950 407682 167010
rect 398235 165612 398301 165613
rect 398235 165548 398236 165612
rect 398300 165548 398301 165612
rect 398235 165547 398301 165548
rect 397131 164388 397197 164389
rect 397131 164324 397132 164388
rect 397196 164324 397197 164388
rect 397131 164323 397197 164324
rect 396027 164252 396093 164253
rect 396027 164188 396028 164252
rect 396092 164188 396093 164252
rect 396027 164187 396093 164188
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 165000
rect 399526 164253 399586 166950
rect 400446 164253 400506 166950
rect 401734 165613 401794 166950
rect 401731 165612 401797 165613
rect 401731 165548 401732 165612
rect 401796 165548 401797 165612
rect 401731 165547 401797 165548
rect 399523 164252 399589 164253
rect 399523 164188 399524 164252
rect 399588 164188 399589 164252
rect 399523 164187 399589 164188
rect 400443 164252 400509 164253
rect 400443 164188 400444 164252
rect 400508 164188 400509 164252
rect 400443 164187 400509 164188
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 165000
rect 403022 164253 403082 166950
rect 404126 164389 404186 166950
rect 405414 165613 405474 166950
rect 405411 165612 405477 165613
rect 405411 165548 405412 165612
rect 405476 165548 405477 165612
rect 405411 165547 405477 165548
rect 404123 164388 404189 164389
rect 404123 164324 404124 164388
rect 404188 164324 404189 164388
rect 404123 164323 404189 164324
rect 403019 164252 403085 164253
rect 403019 164188 403020 164252
rect 403084 164188 403085 164252
rect 403019 164187 403085 164188
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 165000
rect 406518 164253 406578 166950
rect 407622 164253 407682 166950
rect 408174 166950 408356 167010
rect 408704 167010 408764 167106
rect 410064 167010 410124 167106
rect 408704 166950 408786 167010
rect 408174 164933 408234 166950
rect 408171 164932 408237 164933
rect 408171 164868 408172 164932
rect 408236 164868 408237 164932
rect 408171 164867 408237 164868
rect 408726 164253 408786 166950
rect 410014 166950 410124 167010
rect 410744 167010 410804 167106
rect 411288 167010 411348 167106
rect 412376 167010 412436 167106
rect 413464 167010 413524 167106
rect 410744 166950 410810 167010
rect 411288 166950 411362 167010
rect 412376 166950 412466 167010
rect 406515 164252 406581 164253
rect 406515 164188 406516 164252
rect 406580 164188 406581 164252
rect 406515 164187 406581 164188
rect 407619 164252 407685 164253
rect 407619 164188 407620 164252
rect 407684 164188 407685 164252
rect 407619 164187 407685 164188
rect 408723 164252 408789 164253
rect 408723 164188 408724 164252
rect 408788 164188 408789 164252
rect 408723 164187 408789 164188
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 165000
rect 410014 164253 410074 166950
rect 410750 165613 410810 166950
rect 410747 165612 410813 165613
rect 410747 165548 410748 165612
rect 410812 165548 410813 165612
rect 410747 165547 410813 165548
rect 411302 164253 411362 166950
rect 412406 164389 412466 166950
rect 413326 166950 413524 167010
rect 413600 167010 413660 167106
rect 414552 167010 414612 167106
rect 415912 167010 415972 167106
rect 413600 166950 413754 167010
rect 412403 164388 412469 164389
rect 412403 164324 412404 164388
rect 412468 164324 412469 164388
rect 412403 164323 412469 164324
rect 413326 164253 413386 166950
rect 413694 164797 413754 166950
rect 414430 166950 414612 167010
rect 415902 166950 415972 167010
rect 416048 167010 416108 167106
rect 417000 167010 417060 167106
rect 418088 167010 418148 167106
rect 418496 167010 418556 167106
rect 419448 167010 419508 167106
rect 416048 166950 416146 167010
rect 417000 166950 417066 167010
rect 418088 166950 418354 167010
rect 413691 164796 413757 164797
rect 413691 164732 413692 164796
rect 413756 164732 413757 164796
rect 413691 164731 413757 164732
rect 414430 164253 414490 166950
rect 415902 165613 415962 166950
rect 416086 165613 416146 166950
rect 415899 165612 415965 165613
rect 415899 165548 415900 165612
rect 415964 165548 415965 165612
rect 415899 165547 415965 165548
rect 416083 165612 416149 165613
rect 416083 165548 416084 165612
rect 416148 165548 416149 165612
rect 416083 165547 416149 165548
rect 410011 164252 410077 164253
rect 410011 164188 410012 164252
rect 410076 164188 410077 164252
rect 410011 164187 410077 164188
rect 411299 164252 411365 164253
rect 411299 164188 411300 164252
rect 411364 164188 411365 164252
rect 411299 164187 411365 164188
rect 413323 164252 413389 164253
rect 413323 164188 413324 164252
rect 413388 164188 413389 164252
rect 413323 164187 413389 164188
rect 414427 164252 414493 164253
rect 414427 164188 414428 164252
rect 414492 164188 414493 164252
rect 414427 164187 414493 164188
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 165000
rect 417006 164253 417066 166950
rect 418294 164253 418354 166950
rect 418478 166950 418556 167010
rect 419398 166950 419508 167010
rect 420672 167010 420732 167106
rect 421080 167010 421140 167106
rect 420672 166950 420746 167010
rect 418478 166837 418538 166950
rect 418475 166836 418541 166837
rect 418475 166772 418476 166836
rect 418540 166772 418541 166836
rect 418475 166771 418541 166772
rect 419398 165613 419458 166950
rect 419395 165612 419461 165613
rect 419395 165548 419396 165612
rect 419460 165548 419461 165612
rect 419395 165547 419461 165548
rect 417003 164252 417069 164253
rect 417003 164188 417004 164252
rect 417068 164188 417069 164252
rect 417003 164187 417069 164188
rect 418291 164252 418357 164253
rect 418291 164188 418292 164252
rect 418356 164188 418357 164252
rect 418291 164187 418357 164188
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 165000
rect 420686 164253 420746 166950
rect 421054 166950 421140 167010
rect 421760 167010 421820 167106
rect 422848 167010 422908 167106
rect 423528 167010 423588 167106
rect 423936 167010 423996 167106
rect 425296 167010 425356 167106
rect 421760 166950 421850 167010
rect 422848 166950 422954 167010
rect 421054 166837 421114 166950
rect 421051 166836 421117 166837
rect 421051 166772 421052 166836
rect 421116 166772 421117 166836
rect 421051 166771 421117 166772
rect 421790 164797 421850 166950
rect 421787 164796 421853 164797
rect 421787 164732 421788 164796
rect 421852 164732 421853 164796
rect 421787 164731 421853 164732
rect 422894 164253 422954 166950
rect 423446 166950 423588 167010
rect 423814 166950 423996 167010
rect 425286 166950 425356 167010
rect 425976 167010 426036 167106
rect 426384 167010 426444 167106
rect 427608 167010 427668 167106
rect 428288 167010 428348 167106
rect 425976 166950 426082 167010
rect 426384 166950 426450 167010
rect 427608 166950 427738 167010
rect 423446 166837 423506 166950
rect 423443 166836 423509 166837
rect 423443 166772 423444 166836
rect 423508 166772 423509 166836
rect 423443 166771 423509 166772
rect 423814 165613 423874 166950
rect 423811 165612 423877 165613
rect 423811 165548 423812 165612
rect 423876 165548 423877 165612
rect 423811 165547 423877 165548
rect 420683 164252 420749 164253
rect 420683 164188 420684 164252
rect 420748 164188 420749 164252
rect 420683 164187 420749 164188
rect 422891 164252 422957 164253
rect 422891 164188 422892 164252
rect 422956 164188 422957 164252
rect 422891 164187 422957 164188
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 155834 423854 165000
rect 425286 164253 425346 166950
rect 426022 165069 426082 166950
rect 426019 165068 426085 165069
rect 426019 165004 426020 165068
rect 426084 165004 426085 165068
rect 426019 165003 426085 165004
rect 426390 164389 426450 166950
rect 426387 164388 426453 164389
rect 426387 164324 426388 164388
rect 426452 164324 426453 164388
rect 426387 164323 426453 164324
rect 425283 164252 425349 164253
rect 425283 164188 425284 164252
rect 425348 164188 425349 164252
rect 425283 164187 425349 164188
rect 423234 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 423854 155834
rect 423234 155514 423854 155598
rect 423234 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 423854 155514
rect 423234 145308 423854 155278
rect 426954 157674 427574 165000
rect 427678 164253 427738 166950
rect 428230 166950 428348 167010
rect 428696 167010 428756 167106
rect 429784 167010 429844 167106
rect 431008 167010 431068 167106
rect 428696 166950 428842 167010
rect 428230 166837 428290 166950
rect 428227 166836 428293 166837
rect 428227 166772 428228 166836
rect 428292 166772 428293 166836
rect 428227 166771 428293 166772
rect 428782 164253 428842 166950
rect 429702 166950 429844 167010
rect 430990 166950 431068 167010
rect 431144 167010 431204 167106
rect 432232 167010 432292 167106
rect 433320 167010 433380 167106
rect 433592 167010 433652 167106
rect 434408 167010 434468 167106
rect 431144 166950 431234 167010
rect 432232 166950 432338 167010
rect 433320 166950 433442 167010
rect 429702 164389 429762 166950
rect 429699 164388 429765 164389
rect 429699 164324 429700 164388
rect 429764 164324 429765 164388
rect 429699 164323 429765 164324
rect 430990 164253 431050 166950
rect 431174 164797 431234 166950
rect 431171 164796 431237 164797
rect 431171 164732 431172 164796
rect 431236 164732 431237 164796
rect 431171 164731 431237 164732
rect 432278 164253 432338 166950
rect 433382 164253 433442 166950
rect 433566 166950 433652 167010
rect 434302 166950 434468 167010
rect 435768 167010 435828 167106
rect 436040 167010 436100 167106
rect 436992 167010 437052 167106
rect 438080 167010 438140 167106
rect 435768 166950 435834 167010
rect 433566 164933 433626 166950
rect 434302 165613 434362 166950
rect 434299 165612 434365 165613
rect 434299 165548 434300 165612
rect 434364 165548 434365 165612
rect 434299 165547 434365 165548
rect 433563 164932 433629 164933
rect 433563 164868 433564 164932
rect 433628 164868 433629 164932
rect 433563 164867 433629 164868
rect 427675 164252 427741 164253
rect 427675 164188 427676 164252
rect 427740 164188 427741 164252
rect 427675 164187 427741 164188
rect 428779 164252 428845 164253
rect 428779 164188 428780 164252
rect 428844 164188 428845 164252
rect 428779 164187 428845 164188
rect 430987 164252 431053 164253
rect 430987 164188 430988 164252
rect 431052 164188 431053 164252
rect 430987 164187 431053 164188
rect 432275 164252 432341 164253
rect 432275 164188 432276 164252
rect 432340 164188 432341 164252
rect 432275 164187 432341 164188
rect 433379 164252 433445 164253
rect 433379 164188 433380 164252
rect 433444 164188 433445 164252
rect 433379 164187 433445 164188
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 165000
rect 435774 164253 435834 166950
rect 435958 166950 436100 167010
rect 436878 166950 437052 167010
rect 437798 166950 438140 167010
rect 438488 167010 438548 167106
rect 439168 167010 439228 167106
rect 440936 167010 440996 167106
rect 443520 167010 443580 167106
rect 445968 167010 446028 167106
rect 438488 166950 438594 167010
rect 439168 166950 439330 167010
rect 435958 165613 436018 166950
rect 436878 165613 436938 166950
rect 437798 165613 437858 166950
rect 438534 165613 438594 166950
rect 439270 165613 439330 166950
rect 440926 166950 440996 167010
rect 443502 166950 443580 167010
rect 445894 166950 446028 167010
rect 448280 167010 448340 167106
rect 451000 167010 451060 167106
rect 453448 167010 453508 167106
rect 455896 167010 455956 167106
rect 448280 166950 448346 167010
rect 451000 166950 451106 167010
rect 435955 165612 436021 165613
rect 435955 165548 435956 165612
rect 436020 165548 436021 165612
rect 435955 165547 436021 165548
rect 436875 165612 436941 165613
rect 436875 165548 436876 165612
rect 436940 165548 436941 165612
rect 436875 165547 436941 165548
rect 437795 165612 437861 165613
rect 437795 165548 437796 165612
rect 437860 165548 437861 165612
rect 437795 165547 437861 165548
rect 438531 165612 438597 165613
rect 438531 165548 438532 165612
rect 438596 165548 438597 165612
rect 438531 165547 438597 165548
rect 439267 165612 439333 165613
rect 439267 165548 439268 165612
rect 439332 165548 439333 165612
rect 439267 165547 439333 165548
rect 440926 165069 440986 166950
rect 443502 165613 443562 166950
rect 445894 166837 445954 166950
rect 445891 166836 445957 166837
rect 445891 166772 445892 166836
rect 445956 166772 445957 166836
rect 445891 166771 445957 166772
rect 448286 165613 448346 166950
rect 451046 165613 451106 166950
rect 453438 166950 453508 167010
rect 455830 166950 455956 167010
rect 453438 165613 453498 166950
rect 455830 165613 455890 166950
rect 458480 166290 458540 167106
rect 458406 166230 458540 166290
rect 460928 166290 460988 167106
rect 463512 166290 463572 167106
rect 465960 166290 466020 167106
rect 468544 166290 468604 167106
rect 470992 166837 471052 167106
rect 473440 166837 473500 167106
rect 475888 166837 475948 167106
rect 478472 166837 478532 167106
rect 480920 166837 480980 167106
rect 470989 166836 471055 166837
rect 470989 166772 470990 166836
rect 471054 166772 471055 166836
rect 470989 166771 471055 166772
rect 473437 166836 473503 166837
rect 473437 166772 473438 166836
rect 473502 166772 473503 166836
rect 473437 166771 473503 166772
rect 475885 166836 475951 166837
rect 475885 166772 475886 166836
rect 475950 166772 475951 166836
rect 475885 166771 475951 166772
rect 478469 166836 478535 166837
rect 478469 166772 478470 166836
rect 478534 166772 478535 166836
rect 478469 166771 478535 166772
rect 480917 166836 480983 166837
rect 480917 166772 480918 166836
rect 480982 166772 480983 166836
rect 480917 166771 480983 166772
rect 483368 166701 483428 167106
rect 485952 166701 486012 167106
rect 483365 166700 483431 166701
rect 483365 166636 483366 166700
rect 483430 166636 483431 166700
rect 483365 166635 483431 166636
rect 485949 166700 486015 166701
rect 485949 166636 485950 166700
rect 486014 166636 486015 166700
rect 485949 166635 486015 166636
rect 503224 166565 503284 167106
rect 503221 166564 503287 166565
rect 503221 166500 503222 166564
rect 503286 166500 503287 166564
rect 503221 166499 503287 166500
rect 503360 166290 503420 167106
rect 460928 166230 461042 166290
rect 463512 166230 463618 166290
rect 458406 165613 458466 166230
rect 443499 165612 443565 165613
rect 443499 165548 443500 165612
rect 443564 165548 443565 165612
rect 443499 165547 443565 165548
rect 448283 165612 448349 165613
rect 448283 165548 448284 165612
rect 448348 165548 448349 165612
rect 448283 165547 448349 165548
rect 451043 165612 451109 165613
rect 451043 165548 451044 165612
rect 451108 165548 451109 165612
rect 451043 165547 451109 165548
rect 453435 165612 453501 165613
rect 453435 165548 453436 165612
rect 453500 165548 453501 165612
rect 453435 165547 453501 165548
rect 455827 165612 455893 165613
rect 455827 165548 455828 165612
rect 455892 165548 455893 165612
rect 455827 165547 455893 165548
rect 458403 165612 458469 165613
rect 458403 165548 458404 165612
rect 458468 165548 458469 165612
rect 458403 165547 458469 165548
rect 460982 165205 461042 166230
rect 463558 165341 463618 166230
rect 465950 166230 466020 166290
rect 468526 166230 468604 166290
rect 503302 166230 503420 166290
rect 463555 165340 463621 165341
rect 463555 165276 463556 165340
rect 463620 165276 463621 165340
rect 463555 165275 463621 165276
rect 460979 165204 461045 165205
rect 460979 165140 460980 165204
rect 461044 165140 461045 165204
rect 460979 165139 461045 165140
rect 440923 165068 440989 165069
rect 440923 165004 440924 165068
rect 440988 165004 440989 165068
rect 440923 165003 440989 165004
rect 435771 164252 435837 164253
rect 435771 164188 435772 164252
rect 435836 164188 435837 164252
rect 435771 164187 435837 164188
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 165000
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 165000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 165000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 165000
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 165000
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 155834 459854 165000
rect 459234 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 459854 155834
rect 459234 155514 459854 155598
rect 459234 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 459854 155514
rect 459234 145308 459854 155278
rect 462954 157674 463574 165000
rect 465950 164661 466010 166230
rect 468526 165477 468586 166230
rect 503302 165613 503362 166230
rect 503299 165612 503365 165613
rect 503299 165548 503300 165612
rect 503364 165548 503365 165612
rect 503299 165547 503365 165548
rect 468523 165476 468589 165477
rect 468523 165412 468524 165476
rect 468588 165412 468589 165476
rect 468523 165411 468589 165412
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 465947 164660 466013 164661
rect 465947 164596 465948 164660
rect 466012 164596 466013 164660
rect 465947 164595 466013 164596
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 165000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 165000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 165000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 165000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 165000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 165000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 155834 495854 165000
rect 495234 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 495234 155514 495854 155598
rect 495234 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 495234 145308 495854 155278
rect 498954 157674 499574 165000
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 165000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 165000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 165000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 145484 510909 145485
rect 510843 145420 510844 145484
rect 510908 145420 510909 145484
rect 510843 145419 510909 145420
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 145419
rect 513234 145308 513854 154338
rect 516954 158614 517574 165000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 397141 59739 397207 59740
rect 398232 59530 398292 60106
rect 399592 59666 399652 60106
rect 400544 59666 400604 60106
rect 399526 59606 399652 59666
rect 400446 59606 400604 59666
rect 398232 59470 398298 59530
rect 398238 58173 398298 59470
rect 398235 58172 398301 58173
rect 398235 58108 398236 58172
rect 398300 58108 398301 58172
rect 398235 58107 398301 58108
rect 379099 57492 379165 57493
rect 379099 57428 379100 57492
rect 379164 57428 379165 57492
rect 379099 57427 379165 57428
rect 379794 57454 380414 58000
rect 378915 57220 378981 57221
rect 378915 57156 378916 57220
rect 378980 57156 378981 57220
rect 378915 57155 378981 57156
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 378731 57084 378797 57085
rect 378731 57020 378732 57084
rect 378796 57020 378797 57084
rect 378731 57019 378797 57020
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 377811 56268 377877 56269
rect 377811 56204 377812 56268
rect 377876 56204 377877 56268
rect 377811 56203 377877 56204
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59606
rect 400446 57901 400506 59606
rect 401768 59530 401828 60106
rect 403128 59669 403188 60106
rect 404216 59669 404276 60106
rect 403125 59668 403191 59669
rect 403125 59604 403126 59668
rect 403190 59604 403191 59668
rect 403125 59603 403191 59604
rect 404213 59668 404279 59669
rect 404213 59604 404214 59668
rect 404278 59604 404279 59668
rect 404213 59603 404279 59604
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 405414 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 405414 58173 405474 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 405411 58172 405477 58173
rect 405411 58108 405412 58172
rect 405476 58108 405477 58172
rect 405411 58107 405477 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59533 410804 60106
rect 410744 59532 410813 59533
rect 410744 59470 410748 59532
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410747 59468 410748 59470
rect 410812 59468 410813 59532
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59669 413524 60106
rect 413461 59668 413527 59669
rect 413461 59604 413462 59668
rect 413526 59604 413527 59668
rect 413461 59603 413527 59604
rect 413600 59530 413660 60106
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 410747 59467 410813 59468
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 59470 413660 59530
rect 414552 59530 414612 60106
rect 415912 59530 415972 60106
rect 416048 59669 416108 60106
rect 417000 59805 417060 60106
rect 416997 59804 417063 59805
rect 416997 59740 416998 59804
rect 417062 59740 417063 59804
rect 416997 59739 417063 59740
rect 416045 59668 416111 59669
rect 416045 59604 416046 59668
rect 416110 59604 416111 59668
rect 416045 59603 416111 59604
rect 414552 59470 414674 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413510 57085 413570 59470
rect 414614 57901 414674 59470
rect 415534 59470 415972 59530
rect 418088 59533 418148 60106
rect 418088 59532 418173 59533
rect 418088 59470 418108 59532
rect 415534 57901 415594 59470
rect 418107 59468 418108 59470
rect 418172 59468 418173 59532
rect 418496 59530 418556 60106
rect 419448 59669 419508 60106
rect 419445 59668 419511 59669
rect 419445 59604 419446 59668
rect 419510 59604 419511 59668
rect 419445 59603 419511 59604
rect 418107 59467 418173 59468
rect 418478 59470 418556 59530
rect 420672 59533 420732 60106
rect 420672 59532 420749 59533
rect 420672 59470 420684 59532
rect 414611 57900 414677 57901
rect 414611 57836 414612 57900
rect 414676 57836 414677 57900
rect 414611 57835 414677 57836
rect 415531 57900 415597 57901
rect 415531 57836 415532 57900
rect 415596 57836 415597 57900
rect 415531 57835 415597 57836
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 418478 57221 418538 59470
rect 420683 59468 420684 59470
rect 420748 59468 420749 59532
rect 421080 59530 421140 60106
rect 421760 59669 421820 60106
rect 421757 59668 421823 59669
rect 421757 59604 421758 59668
rect 421822 59604 421823 59668
rect 421757 59603 421823 59604
rect 420683 59467 420749 59468
rect 421054 59470 421140 59530
rect 422848 59530 422908 60106
rect 423528 59805 423588 60106
rect 423936 59805 423996 60106
rect 423525 59804 423591 59805
rect 423525 59740 423526 59804
rect 423590 59740 423591 59804
rect 423525 59739 423591 59740
rect 423933 59804 423999 59805
rect 423933 59740 423934 59804
rect 423998 59740 423999 59804
rect 423933 59739 423999 59740
rect 425296 59530 425356 60106
rect 422848 59470 422954 59530
rect 415794 57134 416414 57218
rect 418475 57220 418541 57221
rect 418475 57156 418476 57220
rect 418540 57156 418541 57220
rect 418475 57155 418541 57156
rect 413507 57084 413573 57085
rect 413507 57020 413508 57084
rect 413572 57020 413573 57084
rect 413507 57019 413573 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 421054 56541 421114 59470
rect 422894 59397 422954 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 422891 59396 422957 59397
rect 422891 59332 422892 59396
rect 422956 59332 422957 59396
rect 422891 59331 422957 59332
rect 421051 56540 421117 56541
rect 421051 56476 421052 56540
rect 421116 56476 421117 56540
rect 421051 56475 421117 56476
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 425286 56269 425346 59470
rect 426022 59397 426082 59470
rect 426019 59396 426085 59397
rect 426019 59332 426020 59396
rect 426084 59332 426085 59396
rect 426019 59331 426085 59332
rect 426390 57901 426450 59470
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 425283 56268 425349 56269
rect 425283 56204 425284 56268
rect 425348 56204 425349 56268
rect 425283 56203 425349 56204
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57901 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 427675 57900 427741 57901
rect 427675 57836 427676 57900
rect 427740 57836 427741 57900
rect 427675 57835 427741 57836
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430990 57221 431050 59470
rect 431174 57901 431234 59470
rect 432278 57901 432338 59470
rect 431171 57900 431237 57901
rect 431171 57836 431172 57900
rect 431236 57836 431237 57900
rect 431171 57835 431237 57836
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433382 57629 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433379 57628 433445 57629
rect 433379 57564 433380 57628
rect 433444 57564 433445 57628
rect 433379 57563 433445 57564
rect 433566 57357 433626 59470
rect 433563 57356 433629 57357
rect 433563 57292 433564 57356
rect 433628 57292 433629 57356
rect 433563 57291 433629 57292
rect 430987 57220 431053 57221
rect 430987 57156 430988 57220
rect 431052 57156 431053 57220
rect 430987 57155 431053 57156
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57901 434730 59470
rect 434667 57900 434733 57901
rect 434667 57836 434668 57900
rect 434732 57836 434733 57900
rect 434667 57835 434733 57836
rect 435774 57629 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 436878 57901 436938 59470
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436875 57900 436941 57901
rect 436875 57836 436876 57900
rect 436940 57836 436941 57900
rect 436875 57835 436941 57836
rect 435771 57628 435837 57629
rect 435771 57564 435772 57628
rect 435836 57564 435837 57628
rect 435771 57563 435837 57564
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 57629 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 455896 59530 455956 60106
rect 458480 59669 458540 60106
rect 458477 59668 458543 59669
rect 458477 59604 458478 59668
rect 458542 59604 458543 59668
rect 458477 59603 458543 59604
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 438347 57628 438413 57629
rect 438347 57564 438348 57628
rect 438412 57564 438413 57628
rect 438347 57563 438413 57564
rect 439086 56677 439146 59470
rect 440926 57221 440986 59470
rect 440923 57220 440989 57221
rect 440923 57156 440924 57220
rect 440988 57156 440989 57220
rect 440923 57155 440989 57156
rect 439083 56676 439149 56677
rect 439083 56612 439084 56676
rect 439148 56612 439149 56676
rect 439083 56611 439149 56612
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 56813 443562 59470
rect 443499 56812 443565 56813
rect 443499 56748 443500 56812
rect 443564 56748 443565 56812
rect 443499 56747 443565 56748
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57901 445954 59470
rect 445891 57900 445957 57901
rect 445891 57836 445892 57900
rect 445956 57836 445957 57900
rect 445891 57835 445957 57836
rect 448286 57493 448346 59470
rect 451046 57901 451106 59470
rect 453438 59470 453508 59530
rect 455830 59470 455956 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 453438 59397 453498 59470
rect 453435 59396 453501 59397
rect 453435 59332 453436 59396
rect 453500 59332 453501 59396
rect 453435 59331 453501 59332
rect 455830 58173 455890 59470
rect 455827 58172 455893 58173
rect 455827 58108 455828 58172
rect 455892 58108 455893 58172
rect 455827 58107 455893 58108
rect 451043 57900 451109 57901
rect 451043 57836 451044 57900
rect 451108 57836 451109 57900
rect 451043 57835 451109 57836
rect 448283 57492 448349 57493
rect 448283 57428 448284 57492
rect 448348 57428 448349 57492
rect 448283 57427 448349 57428
rect 451794 57454 452414 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 57901 461042 59470
rect 463558 58717 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59530 480980 60106
rect 473440 59470 473554 59530
rect 463555 58716 463621 58717
rect 463555 58652 463556 58716
rect 463620 58652 463621 58716
rect 463555 58651 463621 58652
rect 460979 57900 461045 57901
rect 460979 57836 460980 57900
rect 461044 57836 461045 57900
rect 460979 57835 461045 57836
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 465950 57901 466010 59470
rect 468526 58989 468586 59470
rect 468523 58988 468589 58989
rect 468523 58924 468524 58988
rect 468588 58924 468589 58988
rect 468523 58923 468589 58924
rect 465947 57900 466013 57901
rect 465947 57836 465948 57900
rect 466012 57836 466013 57900
rect 465947 57835 466013 57836
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 470918 57901 470978 59470
rect 473494 58853 473554 59470
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 480854 59470 480980 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59669 503284 60106
rect 503221 59668 503287 59669
rect 503221 59604 503222 59668
rect 503286 59604 503287 59668
rect 503221 59603 503287 59604
rect 503360 59530 503420 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 475886 58989 475946 59470
rect 475883 58988 475949 58989
rect 475883 58924 475884 58988
rect 475948 58924 475949 58988
rect 475883 58923 475949 58924
rect 473491 58852 473557 58853
rect 473491 58788 473492 58852
rect 473556 58788 473557 58852
rect 473491 58787 473557 58788
rect 470915 57900 470981 57901
rect 470915 57836 470916 57900
rect 470980 57836 470981 57900
rect 470915 57835 470981 57836
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 478462 57901 478522 59470
rect 480854 59261 480914 59470
rect 480851 59260 480917 59261
rect 480851 59196 480852 59260
rect 480916 59196 480917 59260
rect 480851 59195 480917 59196
rect 483430 59125 483490 59470
rect 483427 59124 483493 59125
rect 483427 59060 483428 59124
rect 483492 59060 483493 59124
rect 483427 59059 483493 59060
rect 478459 57900 478525 57901
rect 478459 57836 478460 57900
rect 478524 57836 478525 57900
rect 478459 57835 478525 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 486006 57901 486066 59470
rect 503302 59470 503420 59530
rect 486003 57900 486069 57901
rect 486003 57836 486004 57900
rect 486068 57836 486069 57900
rect 486003 57835 486069 57836
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503302 57901 503362 59470
rect 503299 57900 503365 57901
rect 503299 57836 503300 57900
rect 503364 57836 503365 57900
rect 503299 57835 503365 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 79610 633218 79846 633454
rect 79610 632898 79846 633134
rect 110330 633218 110566 633454
rect 110330 632898 110566 633134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 562158 74062 562394
rect 74146 562158 74382 562394
rect 73826 561838 74062 562074
rect 74146 561838 74382 562074
rect 77546 563998 77782 564234
rect 77866 563998 78102 564234
rect 77546 563678 77782 563914
rect 77866 563678 78102 563914
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 562158 110062 562394
rect 110146 562158 110382 562394
rect 109826 561838 110062 562074
rect 110146 561838 110382 562074
rect 113546 563998 113782 564234
rect 113866 563998 114102 564234
rect 113546 563678 113782 563914
rect 113866 563678 114102 563914
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 169610 633218 169846 633454
rect 169610 632898 169846 633134
rect 200330 633218 200566 633454
rect 200330 632898 200566 633134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 154250 615218 154486 615454
rect 154250 614898 154486 615134
rect 184970 615218 185206 615454
rect 184970 614898 185206 615134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 169610 597218 169846 597454
rect 169610 596898 169846 597134
rect 200330 597218 200566 597454
rect 200330 596898 200566 597134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 154250 579218 154486 579454
rect 154250 578898 154486 579134
rect 184970 579218 185206 579454
rect 184970 578898 185206 579134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 145826 562158 146062 562394
rect 146146 562158 146382 562394
rect 145826 561838 146062 562074
rect 146146 561838 146382 562074
rect 149546 563998 149782 564234
rect 149866 563998 150102 564234
rect 149546 563678 149782 563914
rect 149866 563678 150102 563914
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 562158 182062 562394
rect 182146 562158 182382 562394
rect 181826 561838 182062 562074
rect 182146 561838 182382 562074
rect 185546 563998 185782 564234
rect 185866 563998 186102 564234
rect 185546 563678 185782 563914
rect 185866 563678 186102 563914
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 562158 218062 562394
rect 218146 562158 218382 562394
rect 217826 561838 218062 562074
rect 218146 561838 218382 562074
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 563998 221782 564234
rect 221866 563998 222102 564234
rect 221546 563678 221782 563914
rect 221866 563678 222102 563914
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 259610 633218 259846 633454
rect 259610 632898 259846 633134
rect 290330 633218 290566 633454
rect 290330 632898 290566 633134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 244250 615218 244486 615454
rect 244250 614898 244486 615134
rect 274970 615218 275206 615454
rect 274970 614898 275206 615134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 259610 597218 259846 597454
rect 259610 596898 259846 597134
rect 290330 597218 290566 597454
rect 290330 596898 290566 597134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 244250 579218 244486 579454
rect 244250 578898 244486 579134
rect 274970 579218 275206 579454
rect 274970 578898 275206 579134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 562158 254062 562394
rect 254146 562158 254382 562394
rect 253826 561838 254062 562074
rect 254146 561838 254382 562074
rect 257546 563998 257782 564234
rect 257866 563998 258102 564234
rect 257546 563678 257782 563914
rect 257866 563678 258102 563914
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 562158 290062 562394
rect 290146 562158 290382 562394
rect 289826 561838 290062 562074
rect 290146 561838 290382 562074
rect 293546 563998 293782 564234
rect 293866 563998 294102 564234
rect 293546 563678 293782 563914
rect 293866 563678 294102 563914
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 64250 543218 64486 543454
rect 64250 542898 64486 543134
rect 94970 543218 95206 543454
rect 94970 542898 95206 543134
rect 125690 543218 125926 543454
rect 125690 542898 125926 543134
rect 156410 543218 156646 543454
rect 156410 542898 156646 543134
rect 187130 543218 187366 543454
rect 187130 542898 187366 543134
rect 217850 543218 218086 543454
rect 217850 542898 218086 543134
rect 248570 543218 248806 543454
rect 248570 542898 248806 543134
rect 279290 543218 279526 543454
rect 279290 542898 279526 543134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 475878 59782 476114
rect 59866 475878 60102 476114
rect 59546 475558 59782 475794
rect 59866 475558 60102 475794
rect 63266 477718 63502 477954
rect 63586 477718 63822 477954
rect 63266 477398 63502 477634
rect 63586 477398 63822 477634
rect 66986 481438 67222 481674
rect 67306 481438 67542 481674
rect 66986 481118 67222 481354
rect 67306 481118 67542 481354
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 472158 92062 472394
rect 92146 472158 92382 472394
rect 91826 471838 92062 472074
rect 92146 471838 92382 472074
rect 95546 475878 95782 476114
rect 95866 475878 96102 476114
rect 95546 475558 95782 475794
rect 95866 475558 96102 475794
rect 99266 477718 99502 477954
rect 99586 477718 99822 477954
rect 99266 477398 99502 477634
rect 99586 477398 99822 477634
rect 102986 481438 103222 481674
rect 103306 481438 103542 481674
rect 102986 481118 103222 481354
rect 103306 481118 103542 481354
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 472158 128062 472394
rect 128146 472158 128382 472394
rect 127826 471838 128062 472074
rect 128146 471838 128382 472074
rect 131546 475878 131782 476114
rect 131866 475878 132102 476114
rect 131546 475558 131782 475794
rect 131866 475558 132102 475794
rect 135266 477718 135502 477954
rect 135586 477718 135822 477954
rect 135266 477398 135502 477634
rect 135586 477398 135822 477634
rect 138986 481438 139222 481674
rect 139306 481438 139542 481674
rect 138986 481118 139222 481354
rect 139306 481118 139542 481354
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 472158 164062 472394
rect 164146 472158 164382 472394
rect 163826 471838 164062 472074
rect 164146 471838 164382 472074
rect 167546 475878 167782 476114
rect 167866 475878 168102 476114
rect 167546 475558 167782 475794
rect 167866 475558 168102 475794
rect 171266 477718 171502 477954
rect 171586 477718 171822 477954
rect 171266 477398 171502 477634
rect 171586 477398 171822 477634
rect 174986 481438 175222 481674
rect 175306 481438 175542 481674
rect 174986 481118 175222 481354
rect 175306 481118 175542 481354
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 59546 367878 59782 368114
rect 59866 367878 60102 368114
rect 59546 367558 59782 367794
rect 59866 367558 60102 367794
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 373438 67222 373674
rect 67306 373438 67542 373674
rect 66986 373118 67222 373354
rect 67306 373118 67542 373354
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 367878 95782 368114
rect 95866 367878 96102 368114
rect 95546 367558 95782 367794
rect 95866 367558 96102 367794
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 373438 103222 373674
rect 103306 373438 103542 373674
rect 102986 373118 103222 373354
rect 103306 373118 103542 373354
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 367878 131782 368114
rect 131866 367878 132102 368114
rect 131546 367558 131782 367794
rect 131866 367558 132102 367794
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 373438 139222 373674
rect 139306 373438 139542 373674
rect 138986 373118 139222 373354
rect 139306 373118 139542 373354
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 367878 167782 368114
rect 167866 367878 168102 368114
rect 167546 367558 167782 367794
rect 167866 367558 168102 367794
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 373438 175222 373674
rect 175306 373438 175542 373674
rect 174986 373118 175222 373354
rect 175306 373118 175542 373354
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 155598 63502 155834
rect 63586 155598 63822 155834
rect 63266 155278 63502 155514
rect 63586 155278 63822 155514
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 155598 99502 155834
rect 99586 155598 99822 155834
rect 99266 155278 99502 155514
rect 99586 155278 99822 155514
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 155598 135502 155834
rect 135586 155598 135822 155834
rect 135266 155278 135502 155514
rect 135586 155278 135822 155514
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 155598 171502 155834
rect 171586 155598 171822 155834
rect 171266 155278 171502 155514
rect 171586 155278 171822 155514
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 199826 472158 200062 472394
rect 200146 472158 200382 472394
rect 199826 471838 200062 472074
rect 200146 471838 200382 472074
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 203546 475878 203782 476114
rect 203866 475878 204102 476114
rect 203546 475558 203782 475794
rect 203866 475558 204102 475794
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 367878 203782 368114
rect 203866 367878 204102 368114
rect 203546 367558 203782 367794
rect 203866 367558 204102 367794
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 207266 477718 207502 477954
rect 207586 477718 207822 477954
rect 207266 477398 207502 477634
rect 207586 477398 207822 477634
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 155598 207502 155834
rect 207586 155598 207822 155834
rect 207266 155278 207502 155514
rect 207586 155278 207822 155514
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 210986 481438 211222 481674
rect 211306 481438 211542 481674
rect 210986 481118 211222 481354
rect 211306 481118 211542 481354
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 373438 211222 373674
rect 211306 373438 211542 373674
rect 210986 373118 211222 373354
rect 211306 373118 211542 373354
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 472158 236062 472394
rect 236146 472158 236382 472394
rect 235826 471838 236062 472074
rect 236146 471838 236382 472074
rect 239546 475878 239782 476114
rect 239866 475878 240102 476114
rect 239546 475558 239782 475794
rect 239866 475558 240102 475794
rect 243266 477718 243502 477954
rect 243586 477718 243822 477954
rect 243266 477398 243502 477634
rect 243586 477398 243822 477634
rect 246986 481438 247222 481674
rect 247306 481438 247542 481674
rect 246986 481118 247222 481354
rect 247306 481118 247542 481354
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 472158 272062 472394
rect 272146 472158 272382 472394
rect 271826 471838 272062 472074
rect 272146 471838 272382 472074
rect 275546 475878 275782 476114
rect 275866 475878 276102 476114
rect 275546 475558 275782 475794
rect 275866 475558 276102 475794
rect 279266 477718 279502 477954
rect 279586 477718 279822 477954
rect 279266 477398 279502 477634
rect 279586 477398 279822 477634
rect 282986 481438 283222 481674
rect 283306 481438 283542 481674
rect 282986 481118 283222 481354
rect 283306 481118 283542 481354
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 344610 633218 344846 633454
rect 344610 632898 344846 633134
rect 375330 633218 375566 633454
rect 375330 632898 375566 633134
rect 406050 633218 406286 633454
rect 406050 632898 406286 633134
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 329250 615218 329486 615454
rect 329250 614898 329486 615134
rect 359970 615218 360206 615454
rect 359970 614898 360206 615134
rect 390690 615218 390926 615454
rect 390690 614898 390926 615134
rect 421410 615218 421646 615454
rect 421410 614898 421646 615134
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 344610 597218 344846 597454
rect 344610 596898 344846 597134
rect 375330 597218 375566 597454
rect 375330 596898 375566 597134
rect 406050 597218 406286 597454
rect 406050 596898 406286 597134
rect 329250 579218 329486 579454
rect 329250 578898 329486 579134
rect 359970 579218 360206 579454
rect 359970 578898 360206 579134
rect 390690 579218 390926 579454
rect 390690 578898 390926 579134
rect 421410 579218 421646 579454
rect 421410 578898 421646 579134
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 344610 561218 344846 561454
rect 344610 560898 344846 561134
rect 375330 561218 375566 561454
rect 375330 560898 375566 561134
rect 406050 561218 406286 561454
rect 406050 560898 406286 561134
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 329250 543218 329486 543454
rect 329250 542898 329486 543134
rect 359970 543218 360206 543454
rect 359970 542898 360206 543134
rect 390690 543218 390926 543454
rect 390690 542898 390926 543134
rect 421410 543218 421646 543454
rect 421410 542898 421646 543134
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 367878 239782 368114
rect 239866 367878 240102 368114
rect 239546 367558 239782 367794
rect 239866 367558 240102 367794
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 373438 247222 373674
rect 247306 373438 247542 373674
rect 246986 373118 247222 373354
rect 247306 373118 247542 373354
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 367878 275782 368114
rect 275866 367878 276102 368114
rect 275546 367558 275782 367794
rect 275866 367558 276102 367794
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 373438 283222 373674
rect 283306 373438 283542 373674
rect 282986 373118 283222 373354
rect 283306 373118 283542 373354
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 367878 311782 368114
rect 311866 367878 312102 368114
rect 311546 367558 311782 367794
rect 311866 367558 312102 367794
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 373438 319222 373674
rect 319306 373438 319542 373674
rect 318986 373118 319222 373354
rect 319306 373118 319542 373354
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 367878 347782 368114
rect 347866 367878 348102 368114
rect 347546 367558 347782 367794
rect 347866 367558 348102 367794
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 373438 355222 373674
rect 355306 373438 355542 373674
rect 354986 373118 355222 373354
rect 355306 373118 355542 373354
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 155598 243502 155834
rect 243586 155598 243822 155834
rect 243266 155278 243502 155514
rect 243586 155278 243822 155514
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 155598 279502 155834
rect 279586 155598 279822 155834
rect 279266 155278 279502 155514
rect 279586 155278 279822 155514
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 155598 315502 155834
rect 315586 155598 315822 155834
rect 315266 155278 315502 155514
rect 315586 155278 315822 155514
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 155598 351502 155834
rect 351586 155598 351822 155834
rect 351266 155278 351502 155514
rect 351586 155278 351822 155514
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 367878 383782 368114
rect 383866 367878 384102 368114
rect 383546 367558 383782 367794
rect 383866 367558 384102 367794
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 373438 391222 373674
rect 391306 373438 391542 373674
rect 390986 373118 391222 373354
rect 391306 373118 391542 373354
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 367878 419782 368114
rect 419866 367878 420102 368114
rect 419546 367558 419782 367794
rect 419866 367558 420102 367794
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 373438 427222 373674
rect 427306 373438 427542 373674
rect 426986 373118 427222 373354
rect 427306 373118 427542 373354
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 367878 455782 368114
rect 455866 367878 456102 368114
rect 455546 367558 455782 367794
rect 455866 367558 456102 367794
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 373438 463222 373674
rect 463306 373438 463542 373674
rect 462986 373118 463222 373354
rect 463306 373118 463542 373354
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 367878 491782 368114
rect 491866 367878 492102 368114
rect 491546 367558 491782 367794
rect 491866 367558 492102 367794
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 373438 499222 373674
rect 499306 373438 499542 373674
rect 498986 373118 499222 373354
rect 499306 373118 499542 373354
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 155598 387502 155834
rect 387586 155598 387822 155834
rect 387266 155278 387502 155514
rect 387586 155278 387822 155514
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 155598 423502 155834
rect 423586 155598 423822 155834
rect 423266 155278 423502 155514
rect 423586 155278 423822 155514
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 459266 155598 459502 155834
rect 459586 155598 459822 155834
rect 459266 155278 459502 155514
rect 459586 155278 459822 155514
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 155598 495502 155834
rect 495586 155598 495822 155834
rect 495266 155278 495502 155514
rect 495586 155278 495822 155514
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 79610 633454
rect 79846 633218 110330 633454
rect 110566 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 169610 633454
rect 169846 633218 200330 633454
rect 200566 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 259610 633454
rect 259846 633218 290330 633454
rect 290566 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 344610 633454
rect 344846 633218 375330 633454
rect 375566 633218 406050 633454
rect 406286 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 79610 633134
rect 79846 632898 110330 633134
rect 110566 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 169610 633134
rect 169846 632898 200330 633134
rect 200566 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 259610 633134
rect 259846 632898 290330 633134
rect 290566 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 344610 633134
rect 344846 632898 375330 633134
rect 375566 632898 406050 633134
rect 406286 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 154250 615454
rect 154486 615218 184970 615454
rect 185206 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 244250 615454
rect 244486 615218 274970 615454
rect 275206 615218 329250 615454
rect 329486 615218 359970 615454
rect 360206 615218 390690 615454
rect 390926 615218 421410 615454
rect 421646 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 154250 615134
rect 154486 614898 184970 615134
rect 185206 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 244250 615134
rect 244486 614898 274970 615134
rect 275206 614898 329250 615134
rect 329486 614898 359970 615134
rect 360206 614898 390690 615134
rect 390926 614898 421410 615134
rect 421646 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 169610 597454
rect 169846 597218 200330 597454
rect 200566 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 259610 597454
rect 259846 597218 290330 597454
rect 290566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 344610 597454
rect 344846 597218 375330 597454
rect 375566 597218 406050 597454
rect 406286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 169610 597134
rect 169846 596898 200330 597134
rect 200566 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 259610 597134
rect 259846 596898 290330 597134
rect 290566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 344610 597134
rect 344846 596898 375330 597134
rect 375566 596898 406050 597134
rect 406286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 154250 579454
rect 154486 579218 184970 579454
rect 185206 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 244250 579454
rect 244486 579218 274970 579454
rect 275206 579218 329250 579454
rect 329486 579218 359970 579454
rect 360206 579218 390690 579454
rect 390926 579218 421410 579454
rect 421646 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 154250 579134
rect 154486 578898 184970 579134
rect 185206 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 244250 579134
rect 244486 578898 274970 579134
rect 275206 578898 329250 579134
rect 329486 578898 359970 579134
rect 360206 578898 390690 579134
rect 390926 578898 421410 579134
rect 421646 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect 77514 564234 294134 564266
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 293546 564234
rect 293782 563998 293866 564234
rect 294102 563998 294134 564234
rect 77514 563914 294134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 293546 563914
rect 293782 563678 293866 563914
rect 294102 563678 294134 563914
rect 77514 563646 294134 563678
rect 73794 562394 290414 562426
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 289826 562394
rect 290062 562158 290146 562394
rect 290382 562158 290414 562394
rect 73794 562074 290414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 289826 562074
rect 290062 561838 290146 562074
rect 290382 561838 290414 562074
rect 73794 561806 290414 561838
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 344610 561454
rect 344846 561218 375330 561454
rect 375566 561218 406050 561454
rect 406286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 344610 561134
rect 344846 560898 375330 561134
rect 375566 560898 406050 561134
rect 406286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64250 543454
rect 64486 543218 94970 543454
rect 95206 543218 125690 543454
rect 125926 543218 156410 543454
rect 156646 543218 187130 543454
rect 187366 543218 217850 543454
rect 218086 543218 248570 543454
rect 248806 543218 279290 543454
rect 279526 543218 329250 543454
rect 329486 543218 359970 543454
rect 360206 543218 390690 543454
rect 390926 543218 421410 543454
rect 421646 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64250 543134
rect 64486 542898 94970 543134
rect 95206 542898 125690 543134
rect 125926 542898 156410 543134
rect 156646 542898 187130 543134
rect 187366 542898 217850 543134
rect 218086 542898 248570 543134
rect 248806 542898 279290 543134
rect 279526 542898 329250 543134
rect 329486 542898 359970 543134
rect 360206 542898 390690 543134
rect 390926 542898 421410 543134
rect 421646 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect 66954 481674 283574 481706
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 66954 481354 283574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 66954 481086 283574 481118
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect 63234 477954 279854 477986
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 63234 477634 279854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 63234 477366 279854 477398
rect 59514 476114 276134 476146
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 59514 475794 276134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 59514 475526 276134 475558
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect 91794 472394 272414 472426
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 91794 472074 272414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 91794 471806 272414 471838
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect 66954 373674 499574 373706
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 66954 373354 499574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 66954 373086 499574 373118
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect 59514 368114 492134 368146
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 59514 367794 492134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 59514 367526 492134 367558
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect 63234 155834 495854 155866
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 63234 155514 495854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 63234 155246 495854 155278
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 381000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 575000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 240000 0 1 575000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 150000 0 1 575000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 488000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 325000 0 1 529000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 585000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s 73794 561806 290414 562426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 252308 74414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 252308 110414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 252308 146414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 252308 182414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252308 218414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252308 254414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252308 290414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252308 326414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252308 398414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 252308 434414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 252308 470414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 252308 506414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 359308 74414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 359308 110414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 359308 146414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 359308 182414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 359308 218414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 359308 254414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 359308 290414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 359308 326414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 359308 398414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 359308 434414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 359308 470414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 359308 506414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 466308 74414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 466308 110414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 466308 146414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 466308 182414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 466308 218414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 466308 254414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 466308 290414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 466308 326414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 466308 398414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 466308 434414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 550000 74414 573000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 550000 110414 573000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 550000 182414 573000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 550000 254414 573000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 550000 290414 573000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 466308 470414 583000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 466308 506414 583000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 640099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 640099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 550000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 640099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 550000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 640099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 640099 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 642033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 642033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 642033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 642033 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 637000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 637000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s 77514 563646 294134 564266 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 252308 78134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 252308 114134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 252308 150134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 252308 186134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252308 222134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252308 258134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252308 294134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252308 330134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252308 402134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 252308 438134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 252308 474134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 252308 510134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 359308 78134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 359308 114134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 359308 150134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 359308 186134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 359308 222134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 359308 258134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 359308 294134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 359308 330134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 359308 402134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 359308 438134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 359308 474134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 359308 510134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 466308 78134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 466308 114134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 466308 150134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 466308 186134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 466308 222134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 466308 258134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 466308 294134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 466308 330134 527000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 527000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 466308 402134 527000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 550000 78134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 550000 114134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 550000 150134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 550000 186134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 550000 258134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 550000 294134 573000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 466308 474134 583000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 466308 510134 583000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 640099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 640099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 640099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 640099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 550000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 640099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 640099 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 642033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 642033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 642033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 466308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 637000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 637000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 252308 81854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 252308 117854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 252308 153854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252308 189854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252308 225854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252308 261854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252308 297854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252308 333854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252308 405854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 252308 441854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 252308 477854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 252308 513854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 359308 81854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 359308 117854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 359308 153854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 359308 189854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 359308 225854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 359308 261854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 359308 297854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 359308 333854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 359308 405854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 359308 441854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 359308 477854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 359308 513854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 466308 81854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 466308 117854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 466308 153854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 466308 189854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 466308 225854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 466308 261854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 466308 297854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 466308 333854 527000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 527000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 466308 405854 527000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 550000 81854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 550000 117854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 550000 153854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 550000 189854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 550000 261854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 550000 297854 573000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 466308 477854 583000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 640099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 640099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 640099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 640099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 550000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 640099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 640099 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 642033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 642033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 642033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 466308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 637000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 466308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 252308 85574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 252308 121574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 252308 157574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252308 193574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252308 229574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252308 265574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252308 301574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252308 337574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252308 409574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 252308 445574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 252308 481574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 252308 517574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 359308 85574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 359308 121574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 359308 157574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 359308 193574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 359308 229574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 359308 265574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 359308 301574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 359308 337574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 359308 409574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 359308 445574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 359308 481574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 359308 517574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 466308 85574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 466308 121574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 466308 157574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 466308 193574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 466308 229574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 466308 265574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 466308 301574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 466308 337574 527000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 527000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 466308 409574 527000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 550000 85574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 550000 121574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 550000 157574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 550000 193574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 550000 265574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 550000 301574 573000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 466308 481574 583000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 640099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 640099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 640099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 640099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 550000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 640099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 640099 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 642033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 642033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 642033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 466308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 637000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 466308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 155246 495854 155866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 477366 279854 477986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 252308 63854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 252308 99854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 252308 135854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 252308 171854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252308 243854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252308 279854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252308 315854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252308 351854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252308 387854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 252308 423854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 252308 459854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 252308 495854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 359308 63854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 359308 99854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 359308 135854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 359308 171854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 359308 243854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 359308 279854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 359308 315854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 359308 351854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 359308 387854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 359308 423854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 359308 459854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 359308 495854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 466308 63854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 466308 99854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 466308 135854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 466308 171854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 466308 243854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 466308 279854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 466308 351854 527000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 466308 387854 527000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 466308 423854 527000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 550000 63854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 550000 99854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 550000 171854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 550000 207854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 550000 243854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 550000 279854 573000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 466308 459854 583000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 466308 495854 583000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 640099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 640099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 550000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 640099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 640099 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 640099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 640099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 466308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 642033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 642033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 642033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 637000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 637000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 373086 499574 373706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 481086 283574 481706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 252308 67574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 252308 103574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 252308 139574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 252308 175574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252308 247574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252308 283574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252308 319574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252308 355574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252308 391574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 252308 427574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 252308 463574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 252308 499574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 359308 67574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 359308 103574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 359308 139574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 359308 175574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 359308 247574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 359308 283574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 359308 319574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 359308 355574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 359308 391574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 359308 427574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 359308 463574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 359308 499574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 466308 67574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 466308 103574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 466308 139574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 466308 175574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 466308 247574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 466308 283574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 466308 355574 527000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 466308 391574 527000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 466308 427574 527000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 550000 67574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 550000 103574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 550000 175574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 550000 211574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 550000 247574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 550000 283574 573000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 466308 463574 583000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 466308 499574 583000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 640099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 640099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 550000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 640099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 640099 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 640099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 640099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 466308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 642033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 642033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 642033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 637000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 637000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 471806 272414 472426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 252308 92414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 252308 128414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 252308 164414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252308 236414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252308 272414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252308 308414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252308 344414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252308 380414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 252308 416414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 252308 452414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 252308 488414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 359308 92414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 359308 128414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 359308 164414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 359308 236414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 359308 272414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 359308 308414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 359308 344414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 359308 380414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 359308 416414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 359308 452414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 359308 488414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 466308 92414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 466308 128414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 466308 164414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 466308 236414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 466308 272414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 466308 344414 527000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 466308 380414 527000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 466308 416414 527000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 550000 92414 573000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 550000 164414 573000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 550000 200414 573000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 550000 272414 573000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 466308 488414 583000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 640099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 550000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 640099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 640099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 550000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 640099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 466308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 642033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 642033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 642033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 466308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 637000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 367526 492134 368146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 252308 60134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 252308 96134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 252308 132134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 252308 168134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252308 240134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252308 276134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252308 312134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252308 348134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252308 384134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 252308 420134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 252308 456134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 252308 492134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 359308 60134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 359308 96134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 359308 132134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 359308 168134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 359308 240134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 359308 276134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 359308 312134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 359308 348134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 359308 384134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 359308 420134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 359308 456134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 359308 492134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 466308 60134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 466308 96134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 466308 132134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 466308 168134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 466308 240134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 466308 276134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 466308 348134 527000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 466308 384134 527000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 466308 420134 527000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 550000 60134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 550000 96134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 550000 168134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 550000 204134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 550000 240134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 550000 276134 573000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 466308 492134 583000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 640099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 640099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 550000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 640099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 640099 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 640099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 640099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 466308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 642033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 642033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 642033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 466308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 637000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
